magic
tech EFS8A
magscale 1 2
timestamp 1602873233
<< locali >>
rect 9631 28577 9758 28611
rect 2599 25449 2605 25483
rect 2599 25381 2633 25449
rect 4163 24599 4197 24667
rect 4163 24565 4169 24599
rect 11287 23137 11322 23171
rect 2329 22967 2363 23069
rect 5543 22185 5549 22219
rect 5543 22117 5577 22185
rect 8211 20009 8217 20043
rect 6411 19941 6456 19975
rect 8211 19941 8245 20009
rect 8211 18921 8217 18955
rect 8211 18853 8245 18921
rect 4439 17833 4445 17867
rect 4439 17765 4473 17833
rect 2605 16983 2639 17289
rect 4445 14943 4479 15113
rect 8395 14807 8429 14875
rect 8395 14773 8401 14807
rect 5457 13719 5491 14025
rect 7113 13855 7147 13957
rect 3617 13175 3651 13481
rect 4439 13481 4445 13515
rect 4439 13413 4473 13481
rect 5181 13175 5215 13481
rect 3427 12631 3461 12699
rect 8769 12631 8803 12869
rect 3427 12597 3433 12631
rect 4439 12393 4445 12427
rect 4439 12325 4473 12393
rect 3157 12087 3191 12189
rect 3519 11543 3553 11611
rect 9689 11543 9723 11645
rect 3519 11509 3525 11543
rect 1547 11305 1685 11339
rect 11287 10081 11322 10115
rect 6009 9571 6043 9605
rect 5917 9537 6043 9571
rect 2139 8279 2173 8347
rect 6469 8279 6503 8585
rect 2139 8245 2145 8279
rect 4899 8041 4905 8075
rect 4899 7973 4933 8041
rect 3893 6103 3927 6273
rect 11287 4641 11322 4675
rect 2507 3689 2513 3723
rect 2507 3621 2541 3689
rect 8585 3519 8619 3621
rect 13311 3553 13346 3587
rect 7757 2567 7791 2601
rect 7665 2533 7791 2567
<< viali >>
rect 7849 35241 7883 35275
rect 7665 35105 7699 35139
rect 8493 34697 8527 34731
rect 9873 34697 9907 34731
rect 13369 34697 13403 34731
rect 4721 34629 4755 34663
rect 7021 34629 7055 34663
rect 6561 34561 6595 34595
rect 4537 34493 4571 34527
rect 6837 34493 6871 34527
rect 8309 34493 8343 34527
rect 8861 34493 8895 34527
rect 9689 34493 9723 34527
rect 10241 34493 10275 34527
rect 13185 34493 13219 34527
rect 13737 34493 13771 34527
rect 5181 34357 5215 34391
rect 7757 34357 7791 34391
rect 8309 34153 8343 34187
rect 8125 34017 8159 34051
rect 8125 33269 8159 33303
rect 1547 30345 1581 30379
rect 1476 30141 1510 30175
rect 1961 30005 1995 30039
rect 7297 30005 7331 30039
rect 7619 29801 7653 29835
rect 6101 29733 6135 29767
rect 7548 29665 7582 29699
rect 6009 29597 6043 29631
rect 6653 29597 6687 29631
rect 8493 29461 8527 29495
rect 6285 29257 6319 29291
rect 7849 29257 7883 29291
rect 4859 29121 4893 29155
rect 8769 29121 8803 29155
rect 4772 29053 4806 29087
rect 5784 29053 5818 29087
rect 5871 28985 5905 29019
rect 6929 28985 6963 29019
rect 7021 28985 7055 29019
rect 7573 28985 7607 29019
rect 8493 28985 8527 29019
rect 8585 28985 8619 29019
rect 5181 28917 5215 28951
rect 5641 28917 5675 28951
rect 6653 28917 6687 28951
rect 8309 28917 8343 28951
rect 5043 28713 5077 28747
rect 5825 28713 5859 28747
rect 6929 28713 6963 28747
rect 7297 28713 7331 28747
rect 6101 28645 6135 28679
rect 7573 28645 7607 28679
rect 7665 28645 7699 28679
rect 4940 28577 4974 28611
rect 9597 28577 9631 28611
rect 6009 28509 6043 28543
rect 6653 28509 6687 28543
rect 7849 28509 7883 28543
rect 5365 28373 5399 28407
rect 9827 28373 9861 28407
rect 10333 28373 10367 28407
rect 3295 28169 3329 28203
rect 4629 28169 4663 28203
rect 4997 28169 5031 28203
rect 8125 28169 8159 28203
rect 10057 28169 10091 28203
rect 3709 28101 3743 28135
rect 7849 28101 7883 28135
rect 10333 28033 10367 28067
rect 10609 28033 10643 28067
rect 3224 27965 3258 27999
rect 4215 27965 4249 27999
rect 6929 27965 6963 27999
rect 5273 27897 5307 27931
rect 5365 27897 5399 27931
rect 5917 27897 5951 27931
rect 7250 27897 7284 27931
rect 8769 27897 8803 27931
rect 8861 27897 8895 27931
rect 9413 27897 9447 27931
rect 10425 27897 10459 27931
rect 4307 27829 4341 27863
rect 6193 27829 6227 27863
rect 6653 27829 6687 27863
rect 8585 27829 8619 27863
rect 9781 27829 9815 27863
rect 4997 27625 5031 27659
rect 6285 27625 6319 27659
rect 8309 27625 8343 27659
rect 5410 27557 5444 27591
rect 7751 27557 7785 27591
rect 9781 27557 9815 27591
rect 9873 27557 9907 27591
rect 3024 27489 3058 27523
rect 4144 27489 4178 27523
rect 6009 27489 6043 27523
rect 11288 27489 11322 27523
rect 3111 27421 3145 27455
rect 5089 27421 5123 27455
rect 7389 27421 7423 27455
rect 8769 27421 8803 27455
rect 11391 27421 11425 27455
rect 10333 27353 10367 27387
rect 3525 27285 3559 27319
rect 4215 27285 4249 27319
rect 7021 27285 7055 27319
rect 3249 27081 3283 27115
rect 4445 27081 4479 27115
rect 5917 27081 5951 27115
rect 10333 27081 10367 27115
rect 11253 27081 11287 27115
rect 3525 26945 3559 26979
rect 6193 26945 6227 26979
rect 7113 26945 7147 26979
rect 7389 26945 7423 26979
rect 10057 26945 10091 26979
rect 2488 26877 2522 26911
rect 4997 26877 5031 26911
rect 7573 26877 7607 26911
rect 8493 26877 8527 26911
rect 9137 26877 9171 26911
rect 3617 26809 3651 26843
rect 4169 26809 4203 26843
rect 5318 26809 5352 26843
rect 7894 26809 7928 26843
rect 9413 26809 9447 26843
rect 9505 26809 9539 26843
rect 2559 26741 2593 26775
rect 2973 26741 3007 26775
rect 4813 26741 4847 26775
rect 6653 26741 6687 26775
rect 8769 26741 8803 26775
rect 2329 26537 2363 26571
rect 4215 26537 4249 26571
rect 6285 26537 6319 26571
rect 8493 26537 8527 26571
rect 9873 26537 9907 26571
rect 2513 26469 2547 26503
rect 2605 26469 2639 26503
rect 5686 26469 5720 26503
rect 7935 26469 7969 26503
rect 4144 26401 4178 26435
rect 6653 26401 6687 26435
rect 3157 26333 3191 26367
rect 5365 26333 5399 26367
rect 7113 26333 7147 26367
rect 7573 26333 7607 26367
rect 3525 26197 3559 26231
rect 4629 26197 4663 26231
rect 5089 26197 5123 26231
rect 7481 26197 7515 26231
rect 9413 26197 9447 26231
rect 4169 25993 4203 26027
rect 6653 25993 6687 26027
rect 1685 25925 1719 25959
rect 1915 25857 1949 25891
rect 4905 25857 4939 25891
rect 6929 25857 6963 25891
rect 7297 25857 7331 25891
rect 8585 25857 8619 25891
rect 1812 25789 1846 25823
rect 2237 25789 2271 25823
rect 2789 25789 2823 25823
rect 3709 25789 3743 25823
rect 3111 25721 3145 25755
rect 4629 25721 4663 25755
rect 4721 25721 4755 25755
rect 7021 25721 7055 25755
rect 8401 25721 8435 25755
rect 8677 25721 8711 25755
rect 9229 25721 9263 25755
rect 2605 25653 2639 25687
rect 5549 25653 5583 25687
rect 6009 25653 6043 25687
rect 7941 25653 7975 25687
rect 2605 25449 2639 25483
rect 5089 25449 5123 25483
rect 7297 25449 7331 25483
rect 10333 25449 10367 25483
rect 4261 25381 4295 25415
rect 5825 25381 5859 25415
rect 7481 25313 7515 25347
rect 7665 25313 7699 25347
rect 10149 25313 10183 25347
rect 2237 25245 2271 25279
rect 3893 25245 3927 25279
rect 4169 25245 4203 25279
rect 4445 25245 4479 25279
rect 5733 25245 5767 25279
rect 6009 25245 6043 25279
rect 3157 25177 3191 25211
rect 3433 25109 3467 25143
rect 6837 25109 6871 25143
rect 8401 25109 8435 25143
rect 8861 25109 8895 25143
rect 10057 25109 10091 25143
rect 3341 24905 3375 24939
rect 4997 24905 5031 24939
rect 5457 24905 5491 24939
rect 10977 24905 11011 24939
rect 4721 24837 4755 24871
rect 2973 24769 3007 24803
rect 6009 24769 6043 24803
rect 10057 24769 10091 24803
rect 1777 24701 1811 24735
rect 2237 24701 2271 24735
rect 2789 24701 2823 24735
rect 3801 24701 3835 24735
rect 5616 24701 5650 24735
rect 6837 24701 6871 24735
rect 7297 24701 7331 24735
rect 8401 24701 8435 24735
rect 8861 24701 8895 24735
rect 6561 24633 6595 24667
rect 10149 24633 10183 24667
rect 10701 24633 10735 24667
rect 2145 24565 2179 24599
rect 3709 24565 3743 24599
rect 4169 24565 4203 24599
rect 5687 24565 5721 24599
rect 6929 24565 6963 24599
rect 7849 24565 7883 24599
rect 8217 24565 8251 24599
rect 8493 24565 8527 24599
rect 9781 24565 9815 24599
rect 2145 24361 2179 24395
rect 2329 24361 2363 24395
rect 7297 24361 7331 24395
rect 7573 24361 7607 24395
rect 11437 24361 11471 24395
rect 4261 24293 4295 24327
rect 4813 24293 4847 24327
rect 6101 24293 6135 24327
rect 9873 24293 9907 24327
rect 2513 24225 2547 24259
rect 2697 24225 2731 24259
rect 7481 24225 7515 24259
rect 7941 24225 7975 24259
rect 11253 24225 11287 24259
rect 4169 24157 4203 24191
rect 6009 24157 6043 24191
rect 6653 24157 6687 24191
rect 9781 24157 9815 24191
rect 10057 24157 10091 24191
rect 3893 24021 3927 24055
rect 5641 24021 5675 24055
rect 8493 24021 8527 24055
rect 1961 23817 1995 23851
rect 4629 23817 4663 23851
rect 6561 23817 6595 23851
rect 7297 23817 7331 23851
rect 8677 23817 8711 23851
rect 10885 23817 10919 23851
rect 9321 23749 9355 23783
rect 2789 23681 2823 23715
rect 4169 23681 4203 23715
rect 5089 23681 5123 23715
rect 7757 23681 7791 23715
rect 2053 23613 2087 23647
rect 2605 23613 2639 23647
rect 3617 23613 3651 23647
rect 4077 23613 4111 23647
rect 9505 23613 9539 23647
rect 9965 23613 9999 23647
rect 11136 23613 11170 23647
rect 3433 23545 3467 23579
rect 5273 23545 5307 23579
rect 5374 23545 5408 23579
rect 5917 23545 5951 23579
rect 7665 23545 7699 23579
rect 8078 23545 8112 23579
rect 3157 23477 3191 23511
rect 6193 23477 6227 23511
rect 8953 23477 8987 23511
rect 9597 23477 9631 23511
rect 10517 23477 10551 23511
rect 11207 23477 11241 23511
rect 11621 23477 11655 23511
rect 11989 23477 12023 23511
rect 1547 23273 1581 23307
rect 4399 23273 4433 23307
rect 4813 23273 4847 23307
rect 5273 23273 5307 23307
rect 6377 23273 6411 23307
rect 6929 23273 6963 23307
rect 7481 23273 7515 23307
rect 8677 23273 8711 23307
rect 10793 23273 10827 23307
rect 5778 23205 5812 23239
rect 8078 23205 8112 23239
rect 1476 23137 1510 23171
rect 2973 23137 3007 23171
rect 4328 23137 4362 23171
rect 9781 23137 9815 23171
rect 10149 23137 10183 23171
rect 11253 23137 11287 23171
rect 2329 23069 2363 23103
rect 3617 23069 3651 23103
rect 5457 23069 5491 23103
rect 7757 23069 7791 23103
rect 10241 23069 10275 23103
rect 11391 23001 11425 23035
rect 2053 22933 2087 22967
rect 2329 22933 2363 22967
rect 2421 22933 2455 22967
rect 3157 22933 3191 22967
rect 2053 22729 2087 22763
rect 3065 22729 3099 22763
rect 3525 22729 3559 22763
rect 7849 22661 7883 22695
rect 4077 22593 4111 22627
rect 4353 22593 4387 22627
rect 5733 22593 5767 22627
rect 6929 22593 6963 22627
rect 7389 22593 7423 22627
rect 8953 22593 8987 22627
rect 10057 22593 10091 22627
rect 10701 22593 10735 22627
rect 5089 22525 5123 22559
rect 8585 22525 8619 22559
rect 8861 22525 8895 22559
rect 4169 22457 4203 22491
rect 6561 22457 6595 22491
rect 7021 22457 7055 22491
rect 10149 22457 10183 22491
rect 1685 22389 1719 22423
rect 2237 22389 2271 22423
rect 3893 22389 3927 22423
rect 5549 22389 5583 22423
rect 6285 22389 6319 22423
rect 8309 22389 8343 22423
rect 9689 22389 9723 22423
rect 11345 22389 11379 22423
rect 2329 22185 2363 22219
rect 5549 22185 5583 22219
rect 6101 22185 6135 22219
rect 7021 22185 7055 22219
rect 9827 22185 9861 22219
rect 10517 22185 10551 22219
rect 1547 22117 1581 22151
rect 2513 22117 2547 22151
rect 2605 22117 2639 22151
rect 1460 22049 1494 22083
rect 4169 22049 4203 22083
rect 7205 22049 7239 22083
rect 7389 22049 7423 22083
rect 8528 22049 8562 22083
rect 9724 22049 9758 22083
rect 10701 22049 10735 22083
rect 3157 21981 3191 22015
rect 5181 21981 5215 22015
rect 8631 21981 8665 22015
rect 10885 21913 10919 21947
rect 1869 21845 1903 21879
rect 4353 21845 4387 21879
rect 5089 21845 5123 21879
rect 8033 21845 8067 21879
rect 9045 21845 9079 21879
rect 10149 21845 10183 21879
rect 2421 21641 2455 21675
rect 4261 21641 4295 21675
rect 5917 21641 5951 21675
rect 7849 21641 7883 21675
rect 9689 21641 9723 21675
rect 6561 21505 6595 21539
rect 10701 21505 10735 21539
rect 1685 21437 1719 21471
rect 1869 21437 1903 21471
rect 2145 21437 2179 21471
rect 2973 21437 3007 21471
rect 4997 21437 5031 21471
rect 6837 21437 6871 21471
rect 7297 21437 7331 21471
rect 8401 21437 8435 21471
rect 8861 21437 8895 21471
rect 2881 21369 2915 21403
rect 3335 21369 3369 21403
rect 5318 21369 5352 21403
rect 9965 21369 9999 21403
rect 3893 21301 3927 21335
rect 4813 21301 4847 21335
rect 6193 21301 6227 21335
rect 6929 21301 6963 21335
rect 8217 21301 8251 21335
rect 8493 21301 8527 21335
rect 1685 21097 1719 21131
rect 2973 21097 3007 21131
rect 3249 21097 3283 21131
rect 4997 21097 5031 21131
rect 5917 21097 5951 21131
rect 7297 21097 7331 21131
rect 8493 21097 8527 21131
rect 2415 21029 2449 21063
rect 3801 21029 3835 21063
rect 4439 21029 4473 21063
rect 5733 21029 5767 21063
rect 8769 21029 8803 21063
rect 9873 21029 9907 21063
rect 5825 20961 5859 20995
rect 6377 20961 6411 20995
rect 7665 20961 7699 20995
rect 7849 20961 7883 20995
rect 11253 20961 11287 20995
rect 2053 20893 2087 20927
rect 4077 20893 4111 20927
rect 7941 20893 7975 20927
rect 9781 20893 9815 20927
rect 10425 20893 10459 20927
rect 5365 20757 5399 20791
rect 6929 20757 6963 20791
rect 10701 20757 10735 20791
rect 11437 20757 11471 20791
rect 2881 20553 2915 20587
rect 4813 20553 4847 20587
rect 5917 20553 5951 20587
rect 9045 20553 9079 20587
rect 9781 20553 9815 20587
rect 6561 20485 6595 20519
rect 1777 20417 1811 20451
rect 3801 20417 3835 20451
rect 4261 20417 4295 20451
rect 9965 20417 9999 20451
rect 1869 20349 1903 20383
rect 2421 20349 2455 20383
rect 5641 20349 5675 20383
rect 5733 20349 5767 20383
rect 7148 20349 7182 20383
rect 7573 20349 7607 20383
rect 8125 20349 8159 20383
rect 9321 20349 9355 20383
rect 2605 20281 2639 20315
rect 3617 20281 3651 20315
rect 3893 20281 3927 20315
rect 6193 20281 6227 20315
rect 7251 20281 7285 20315
rect 8446 20281 8480 20315
rect 10057 20281 10091 20315
rect 10609 20281 10643 20315
rect 8033 20213 8067 20247
rect 10885 20213 10919 20247
rect 11253 20213 11287 20247
rect 1593 20009 1627 20043
rect 3433 20009 3467 20043
rect 8217 20009 8251 20043
rect 8769 20009 8803 20043
rect 9781 20009 9815 20043
rect 13001 20009 13035 20043
rect 3157 19941 3191 19975
rect 4261 19941 4295 19975
rect 4629 19941 4663 19975
rect 4721 19941 4755 19975
rect 6377 19941 6411 19975
rect 10701 19941 10735 19975
rect 11437 19941 11471 19975
rect 1409 19873 1443 19907
rect 2697 19873 2731 19907
rect 2881 19873 2915 19907
rect 7849 19873 7883 19907
rect 9689 19873 9723 19907
rect 10149 19873 10183 19907
rect 12817 19873 12851 19907
rect 4905 19805 4939 19839
rect 6101 19805 6135 19839
rect 7481 19805 7515 19839
rect 11345 19805 11379 19839
rect 11897 19737 11931 19771
rect 1869 19669 1903 19703
rect 2329 19669 2363 19703
rect 7021 19669 7055 19703
rect 9045 19669 9079 19703
rect 9505 19669 9539 19703
rect 1777 19465 1811 19499
rect 4905 19465 4939 19499
rect 5273 19465 5307 19499
rect 6653 19465 6687 19499
rect 7113 19465 7147 19499
rect 10977 19465 11011 19499
rect 11713 19465 11747 19499
rect 12587 19465 12621 19499
rect 3341 19329 3375 19363
rect 6285 19329 6319 19363
rect 7757 19329 7791 19363
rect 8125 19329 8159 19363
rect 9413 19329 9447 19363
rect 10057 19329 10091 19363
rect 2145 19261 2179 19295
rect 2513 19261 2547 19295
rect 2789 19261 2823 19295
rect 4537 19261 4571 19295
rect 5733 19261 5767 19295
rect 7272 19261 7306 19295
rect 8217 19261 8251 19295
rect 10701 19261 10735 19295
rect 12484 19261 12518 19295
rect 12909 19261 12943 19295
rect 2973 19193 3007 19227
rect 3893 19193 3927 19227
rect 3994 19193 4028 19227
rect 8538 19193 8572 19227
rect 10149 19193 10183 19227
rect 11345 19193 11379 19227
rect 13277 19193 13311 19227
rect 3709 19125 3743 19159
rect 5641 19125 5675 19159
rect 5917 19125 5951 19159
rect 7343 19125 7377 19159
rect 9137 19125 9171 19159
rect 9781 19125 9815 19159
rect 1593 18921 1627 18955
rect 6285 18921 6319 18955
rect 8217 18921 8251 18955
rect 9781 18921 9815 18955
rect 10701 18921 10735 18955
rect 4629 18853 4663 18887
rect 11437 18853 11471 18887
rect 1409 18785 1443 18819
rect 2421 18785 2455 18819
rect 2881 18785 2915 18819
rect 6193 18785 6227 18819
rect 6745 18785 6779 18819
rect 7849 18785 7883 18819
rect 8769 18785 8803 18819
rect 9689 18785 9723 18819
rect 10149 18785 10183 18819
rect 12884 18785 12918 18819
rect 1961 18717 1995 18751
rect 2973 18717 3007 18751
rect 3893 18717 3927 18751
rect 4537 18717 4571 18751
rect 4813 18717 4847 18751
rect 11345 18717 11379 18751
rect 11621 18717 11655 18751
rect 2237 18581 2271 18615
rect 9045 18581 9079 18615
rect 12955 18581 12989 18615
rect 2053 18377 2087 18411
rect 3801 18377 3835 18411
rect 4169 18377 4203 18411
rect 6561 18377 6595 18411
rect 7343 18377 7377 18411
rect 12081 18377 12115 18411
rect 13277 18377 13311 18411
rect 6285 18309 6319 18343
rect 7113 18309 7147 18343
rect 8033 18309 8067 18343
rect 9137 18309 9171 18343
rect 11345 18309 11379 18343
rect 2881 18241 2915 18275
rect 5733 18241 5767 18275
rect 8217 18241 8251 18275
rect 10057 18241 10091 18275
rect 11713 18241 11747 18275
rect 1869 18173 1903 18207
rect 5365 18173 5399 18207
rect 7272 18173 7306 18207
rect 10977 18173 11011 18207
rect 12484 18173 12518 18207
rect 12909 18173 12943 18207
rect 13528 18173 13562 18207
rect 3202 18105 3236 18139
rect 4721 18105 4755 18139
rect 4813 18105 4847 18139
rect 7757 18105 7791 18139
rect 8538 18105 8572 18139
rect 10149 18105 10183 18139
rect 10701 18105 10735 18139
rect 1777 18037 1811 18071
rect 2329 18037 2363 18071
rect 2789 18037 2823 18071
rect 4537 18037 4571 18071
rect 9689 18037 9723 18071
rect 12587 18037 12621 18071
rect 13599 18037 13633 18071
rect 13921 18037 13955 18071
rect 3341 17833 3375 17867
rect 4445 17833 4479 17867
rect 4997 17833 5031 17867
rect 8493 17833 8527 17867
rect 2145 17765 2179 17799
rect 3709 17765 3743 17799
rect 6009 17765 6043 17799
rect 8125 17765 8159 17799
rect 9873 17765 9907 17799
rect 10701 17765 10735 17799
rect 11345 17765 11379 17799
rect 11437 17765 11471 17799
rect 4077 17697 4111 17731
rect 7389 17697 7423 17731
rect 7941 17697 7975 17731
rect 10425 17697 10459 17731
rect 12884 17697 12918 17731
rect 2053 17629 2087 17663
rect 2973 17629 3007 17663
rect 5733 17629 5767 17663
rect 5917 17629 5951 17663
rect 6193 17629 6227 17663
rect 9781 17629 9815 17663
rect 2605 17561 2639 17595
rect 11897 17561 11931 17595
rect 1685 17493 1719 17527
rect 5365 17493 5399 17527
rect 8953 17493 8987 17527
rect 12955 17493 12989 17527
rect 2605 17289 2639 17323
rect 6009 17289 6043 17323
rect 9873 17289 9907 17323
rect 10241 17289 10275 17323
rect 11621 17289 11655 17323
rect 13277 17289 13311 17323
rect 1685 17085 1719 17119
rect 1961 17085 1995 17119
rect 13599 17221 13633 17255
rect 6561 17153 6595 17187
rect 7205 17153 7239 17187
rect 8033 17153 8067 17187
rect 8769 17153 8803 17187
rect 8953 17153 8987 17187
rect 10563 17153 10597 17187
rect 11345 17153 11379 17187
rect 2973 17085 3007 17119
rect 4813 17085 4847 17119
rect 7573 17085 7607 17119
rect 7849 17085 7883 17119
rect 8861 17085 8895 17119
rect 9137 17085 9171 17119
rect 10476 17085 10510 17119
rect 10885 17085 10919 17119
rect 12484 17085 12518 17119
rect 12909 17085 12943 17119
rect 13528 17085 13562 17119
rect 13921 17085 13955 17119
rect 2789 17017 2823 17051
rect 3294 17017 3328 17051
rect 4169 17017 4203 17051
rect 4629 17017 4663 17051
rect 5134 17017 5168 17051
rect 12587 17017 12621 17051
rect 1685 16949 1719 16983
rect 2421 16949 2455 16983
rect 2605 16949 2639 16983
rect 3893 16949 3927 16983
rect 5733 16949 5767 16983
rect 8401 16949 8435 16983
rect 9321 16949 9355 16983
rect 2605 16745 2639 16779
rect 3801 16745 3835 16779
rect 5181 16745 5215 16779
rect 7297 16745 7331 16779
rect 12403 16745 12437 16779
rect 2047 16677 2081 16711
rect 4261 16677 4295 16711
rect 5549 16677 5583 16711
rect 5825 16677 5859 16711
rect 8309 16677 8343 16711
rect 1685 16609 1719 16643
rect 7205 16609 7239 16643
rect 7757 16609 7791 16643
rect 9689 16609 9723 16643
rect 9965 16609 9999 16643
rect 11253 16609 11287 16643
rect 12332 16609 12366 16643
rect 4169 16541 4203 16575
rect 4813 16541 4847 16575
rect 5733 16541 5767 16575
rect 6193 16541 6227 16575
rect 10149 16541 10183 16575
rect 8861 16473 8895 16507
rect 9781 16473 9815 16507
rect 11437 16473 11471 16507
rect 3065 16405 3099 16439
rect 3341 16405 3375 16439
rect 6837 16405 6871 16439
rect 9413 16405 9447 16439
rect 2237 16201 2271 16235
rect 4261 16201 4295 16235
rect 4721 16201 4755 16235
rect 5825 16201 5859 16235
rect 6285 16201 6319 16235
rect 7849 16201 7883 16235
rect 8861 16201 8895 16235
rect 11069 16201 11103 16235
rect 12633 16201 12667 16235
rect 1547 16065 1581 16099
rect 5181 16065 5215 16099
rect 7297 16065 7331 16099
rect 9229 16065 9263 16099
rect 9413 16065 9447 16099
rect 10333 16065 10367 16099
rect 1460 15997 1494 16031
rect 2973 15997 3007 16031
rect 6837 15997 6871 16031
rect 6929 15997 6963 16031
rect 7113 15997 7147 16031
rect 10885 15997 10919 16031
rect 11713 15997 11747 16031
rect 1961 15929 1995 15963
rect 2881 15929 2915 15963
rect 3335 15929 3369 15963
rect 4905 15929 4939 15963
rect 4997 15929 5031 15963
rect 6653 15929 6687 15963
rect 9505 15929 9539 15963
rect 10057 15929 10091 15963
rect 11345 15929 11379 15963
rect 3893 15861 3927 15895
rect 8217 15861 8251 15895
rect 1869 15657 1903 15691
rect 3525 15657 3559 15691
rect 5273 15657 5307 15691
rect 12955 15657 12989 15691
rect 1409 15589 1443 15623
rect 3157 15589 3191 15623
rect 4261 15589 4295 15623
rect 4813 15589 4847 15623
rect 9413 15589 9447 15623
rect 9873 15589 9907 15623
rect 11253 15589 11287 15623
rect 2421 15521 2455 15555
rect 2973 15521 3007 15555
rect 6377 15521 6411 15555
rect 7297 15521 7331 15555
rect 7573 15521 7607 15555
rect 11437 15521 11471 15555
rect 12884 15521 12918 15555
rect 3893 15453 3927 15487
rect 4169 15453 4203 15487
rect 6469 15453 6503 15487
rect 7757 15453 7791 15487
rect 9781 15453 9815 15487
rect 10425 15453 10459 15487
rect 2329 15385 2363 15419
rect 6929 15385 6963 15419
rect 7389 15385 7423 15419
rect 8309 15317 8343 15351
rect 8769 15317 8803 15351
rect 1685 15113 1719 15147
rect 4445 15113 4479 15147
rect 4721 15113 4755 15147
rect 7389 15113 7423 15147
rect 7757 15113 7791 15147
rect 9321 15113 9355 15147
rect 10701 15113 10735 15147
rect 11345 15113 11379 15147
rect 2053 15045 2087 15079
rect 2421 15045 2455 15079
rect 3617 15045 3651 15079
rect 3985 15045 4019 15079
rect 3065 14977 3099 15011
rect 6285 14977 6319 15011
rect 8033 14977 8067 15011
rect 1501 14909 1535 14943
rect 2513 14909 2547 14943
rect 2973 14909 3007 14943
rect 4169 14909 4203 14943
rect 4445 14909 4479 14943
rect 5089 14909 5123 14943
rect 5181 14909 5215 14943
rect 5733 14909 5767 14943
rect 5917 14909 5951 14943
rect 6653 14909 6687 14943
rect 6837 14909 6871 14943
rect 9781 14909 9815 14943
rect 12265 14909 12299 14943
rect 12449 14909 12483 14943
rect 12909 14909 12943 14943
rect 9597 14841 9631 14875
rect 10102 14841 10136 14875
rect 4353 14773 4387 14807
rect 7021 14773 7055 14807
rect 8401 14773 8435 14807
rect 8953 14773 8987 14807
rect 12541 14773 12575 14807
rect 13461 14773 13495 14807
rect 4629 14569 4663 14603
rect 7389 14569 7423 14603
rect 9505 14569 9539 14603
rect 11345 14569 11379 14603
rect 1547 14501 1581 14535
rect 3801 14501 3835 14535
rect 4997 14501 5031 14535
rect 9873 14501 9907 14535
rect 10425 14501 10459 14535
rect 12449 14501 12483 14535
rect 1460 14433 1494 14467
rect 2421 14433 2455 14467
rect 2697 14433 2731 14467
rect 3157 14433 3191 14467
rect 6377 14433 6411 14467
rect 6469 14433 6503 14467
rect 6653 14433 6687 14467
rect 7941 14433 7975 14467
rect 8493 14433 8527 14467
rect 11529 14433 11563 14467
rect 11713 14433 11747 14467
rect 12868 14433 12902 14467
rect 1961 14365 1995 14399
rect 4905 14365 4939 14399
rect 6837 14365 6871 14399
rect 8677 14365 8711 14399
rect 9781 14365 9815 14399
rect 12955 14365 12989 14399
rect 2513 14297 2547 14331
rect 5457 14297 5491 14331
rect 2329 14229 2363 14263
rect 3433 14229 3467 14263
rect 4353 14229 4387 14263
rect 9137 14229 9171 14263
rect 2513 14025 2547 14059
rect 5273 14025 5307 14059
rect 5457 14025 5491 14059
rect 5733 14025 5767 14059
rect 6469 14025 6503 14059
rect 7849 14025 7883 14059
rect 9597 14025 9631 14059
rect 9873 14025 9907 14059
rect 11345 14025 11379 14059
rect 12587 14025 12621 14059
rect 13277 14025 13311 14059
rect 4169 13957 4203 13991
rect 4353 13889 4387 13923
rect 1685 13821 1719 13855
rect 2697 13821 2731 13855
rect 3249 13821 3283 13855
rect 4445 13753 4479 13787
rect 4997 13753 5031 13787
rect 7021 13957 7055 13991
rect 7113 13957 7147 13991
rect 7389 13957 7423 13991
rect 9229 13957 9263 13991
rect 8309 13889 8343 13923
rect 10425 13889 10459 13923
rect 11713 13889 11747 13923
rect 6009 13821 6043 13855
rect 6837 13821 6871 13855
rect 7113 13821 7147 13855
rect 12500 13821 12534 13855
rect 13528 13821 13562 13855
rect 8125 13753 8159 13787
rect 8630 13753 8664 13787
rect 10149 13753 10183 13787
rect 10241 13753 10275 13787
rect 13921 13753 13955 13787
rect 1869 13685 1903 13719
rect 2973 13685 3007 13719
rect 3709 13685 3743 13719
rect 5457 13685 5491 13719
rect 12909 13685 12943 13719
rect 13599 13685 13633 13719
rect 3617 13481 3651 13515
rect 3433 13413 3467 13447
rect 2697 13345 2731 13379
rect 2881 13345 2915 13379
rect 1409 13277 1443 13311
rect 3157 13277 3191 13311
rect 4445 13481 4479 13515
rect 5181 13481 5215 13515
rect 7481 13481 7515 13515
rect 8769 13481 8803 13515
rect 9505 13481 9539 13515
rect 10793 13481 10827 13515
rect 4077 13277 4111 13311
rect 3801 13209 3835 13243
rect 4997 13209 5031 13243
rect 1869 13141 1903 13175
rect 2329 13141 2363 13175
rect 3617 13141 3651 13175
rect 6009 13413 6043 13447
rect 6561 13413 6595 13447
rect 8401 13413 8435 13447
rect 9873 13413 9907 13447
rect 11437 13413 11471 13447
rect 7389 13345 7423 13379
rect 7849 13345 7883 13379
rect 5917 13277 5951 13311
rect 9781 13277 9815 13311
rect 10425 13277 10459 13311
rect 11345 13277 11379 13311
rect 11621 13277 11655 13311
rect 5181 13141 5215 13175
rect 5365 13141 5399 13175
rect 8953 12937 8987 12971
rect 13599 12937 13633 12971
rect 13921 12937 13955 12971
rect 8769 12869 8803 12903
rect 11897 12869 11931 12903
rect 4997 12801 5031 12835
rect 7757 12801 7791 12835
rect 1777 12733 1811 12767
rect 2053 12733 2087 12767
rect 3065 12733 3099 12767
rect 7665 12733 7699 12767
rect 8677 12733 8711 12767
rect 2237 12665 2271 12699
rect 4353 12665 4387 12699
rect 4905 12665 4939 12699
rect 5359 12665 5393 12699
rect 6653 12665 6687 12699
rect 8078 12665 8112 12699
rect 9597 12801 9631 12835
rect 10885 12801 10919 12835
rect 11207 12801 11241 12835
rect 12587 12801 12621 12835
rect 11104 12733 11138 12767
rect 11529 12733 11563 12767
rect 12484 12733 12518 12767
rect 12909 12733 12943 12767
rect 13528 12733 13562 12767
rect 9413 12665 9447 12699
rect 9689 12665 9723 12699
rect 10241 12665 10275 12699
rect 2605 12597 2639 12631
rect 2973 12597 3007 12631
rect 3433 12597 3467 12631
rect 3985 12597 4019 12631
rect 5917 12597 5951 12631
rect 6193 12597 6227 12631
rect 7205 12597 7239 12631
rect 8769 12597 8803 12631
rect 10517 12597 10551 12631
rect 2881 12393 2915 12427
rect 3893 12393 3927 12427
rect 4445 12393 4479 12427
rect 4997 12393 5031 12427
rect 5365 12393 5399 12427
rect 8769 12393 8803 12427
rect 11713 12393 11747 12427
rect 12403 12393 12437 12427
rect 2047 12325 2081 12359
rect 6009 12325 6043 12359
rect 8170 12325 8204 12359
rect 9505 12325 9539 12359
rect 9873 12325 9907 12359
rect 10425 12325 10459 12359
rect 4077 12257 4111 12291
rect 11288 12257 11322 12291
rect 12300 12257 12334 12291
rect 1685 12189 1719 12223
rect 3157 12189 3191 12223
rect 3249 12189 3283 12223
rect 5917 12189 5951 12223
rect 6193 12189 6227 12223
rect 6837 12189 6871 12223
rect 7849 12189 7883 12223
rect 9781 12189 9815 12223
rect 5641 12121 5675 12155
rect 11391 12121 11425 12155
rect 2605 12053 2639 12087
rect 3157 12053 3191 12087
rect 7481 12053 7515 12087
rect 3065 11849 3099 11883
rect 4445 11849 4479 11883
rect 4813 11849 4847 11883
rect 6009 11849 6043 11883
rect 8677 11849 8711 11883
rect 9505 11849 9539 11883
rect 12909 11849 12943 11883
rect 4077 11781 4111 11815
rect 6561 11781 6595 11815
rect 1685 11713 1719 11747
rect 2605 11713 2639 11747
rect 3157 11713 3191 11747
rect 4997 11713 5031 11747
rect 6929 11713 6963 11747
rect 7205 11713 7239 11747
rect 2329 11645 2363 11679
rect 5641 11645 5675 11679
rect 8493 11645 8527 11679
rect 9689 11645 9723 11679
rect 9965 11645 9999 11679
rect 10425 11645 10459 11679
rect 12484 11645 12518 11679
rect 13277 11645 13311 11679
rect 1777 11577 1811 11611
rect 5089 11577 5123 11611
rect 7021 11577 7055 11611
rect 12587 11577 12621 11611
rect 3525 11509 3559 11543
rect 7941 11509 7975 11543
rect 8217 11509 8251 11543
rect 9689 11509 9723 11543
rect 9781 11509 9815 11543
rect 10057 11509 10091 11543
rect 11253 11509 11287 11543
rect 1685 11305 1719 11339
rect 2329 11305 2363 11339
rect 3433 11305 3467 11339
rect 4261 11305 4295 11339
rect 4997 11305 5031 11339
rect 9413 11305 9447 11339
rect 9781 11305 9815 11339
rect 11437 11305 11471 11339
rect 3157 11237 3191 11271
rect 5733 11237 5767 11271
rect 6285 11237 6319 11271
rect 8211 11237 8245 11271
rect 9137 11237 9171 11271
rect 1476 11169 1510 11203
rect 2513 11169 2547 11203
rect 2881 11169 2915 11203
rect 4445 11169 4479 11203
rect 9965 11169 9999 11203
rect 10149 11169 10183 11203
rect 11253 11169 11287 11203
rect 3801 11101 3835 11135
rect 5641 11101 5675 11135
rect 7849 11101 7883 11135
rect 4629 11033 4663 11067
rect 6929 11033 6963 11067
rect 7757 11033 7791 11067
rect 1961 10965 1995 10999
rect 7205 10965 7239 10999
rect 8769 10965 8803 10999
rect 2789 10761 2823 10795
rect 3985 10761 4019 10795
rect 5549 10761 5583 10795
rect 10241 10761 10275 10795
rect 10931 10761 10965 10795
rect 5825 10693 5859 10727
rect 3617 10625 3651 10659
rect 4445 10625 4479 10659
rect 7941 10625 7975 10659
rect 8585 10625 8619 10659
rect 1777 10557 1811 10591
rect 2237 10557 2271 10591
rect 3157 10557 3191 10591
rect 5641 10557 5675 10591
rect 6837 10557 6871 10591
rect 7297 10557 7331 10591
rect 7665 10557 7699 10591
rect 9873 10557 9907 10591
rect 10860 10557 10894 10591
rect 11621 10557 11655 10591
rect 1685 10489 1719 10523
rect 4158 10489 4192 10523
rect 4261 10489 4295 10523
rect 9965 10489 9999 10523
rect 1869 10421 1903 10455
rect 5181 10421 5215 10455
rect 6193 10421 6227 10455
rect 6653 10421 6687 10455
rect 8309 10421 8343 10455
rect 9137 10421 9171 10455
rect 11253 10421 11287 10455
rect 1869 10217 1903 10251
rect 2605 10217 2639 10251
rect 4169 10217 4203 10251
rect 6009 10217 6043 10251
rect 8309 10217 8343 10251
rect 12403 10217 12437 10251
rect 2145 10149 2179 10183
rect 9873 10149 9907 10183
rect 2605 10081 2639 10115
rect 2881 10081 2915 10115
rect 4077 10081 4111 10115
rect 4629 10081 4663 10115
rect 6561 10081 6595 10115
rect 7389 10081 7423 10115
rect 11253 10081 11287 10115
rect 12300 10081 12334 10115
rect 3893 10013 3927 10047
rect 7297 10013 7331 10047
rect 8585 10013 8619 10047
rect 9781 10013 9815 10047
rect 7481 9945 7515 9979
rect 10333 9945 10367 9979
rect 5181 9877 5215 9911
rect 5641 9877 5675 9911
rect 6377 9877 6411 9911
rect 9321 9877 9355 9911
rect 10701 9877 10735 9911
rect 11391 9877 11425 9911
rect 3065 9673 3099 9707
rect 4629 9673 4663 9707
rect 7113 9673 7147 9707
rect 9781 9673 9815 9707
rect 12633 9673 12667 9707
rect 6009 9605 6043 9639
rect 3433 9537 3467 9571
rect 8217 9537 8251 9571
rect 10333 9537 10367 9571
rect 1961 9469 1995 9503
rect 2329 9469 2363 9503
rect 2605 9469 2639 9503
rect 3617 9469 3651 9503
rect 4077 9469 4111 9503
rect 5169 9469 5203 9503
rect 5273 9469 5307 9503
rect 5457 9469 5491 9503
rect 7021 9469 7055 9503
rect 7665 9469 7699 9503
rect 4353 9401 4387 9435
rect 5089 9401 5123 9435
rect 6285 9401 6319 9435
rect 6837 9401 6871 9435
rect 8538 9401 8572 9435
rect 10057 9401 10091 9435
rect 10149 9401 10183 9435
rect 2145 9333 2179 9367
rect 6653 9333 6687 9367
rect 8125 9333 8159 9367
rect 9137 9333 9171 9367
rect 11253 9333 11287 9367
rect 2053 9129 2087 9163
rect 3157 9129 3191 9163
rect 3709 9129 3743 9163
rect 7297 9129 7331 9163
rect 9505 9129 9539 9163
rect 11253 9129 11287 9163
rect 2329 9061 2363 9095
rect 4261 9061 4295 9095
rect 7843 9061 7877 9095
rect 9781 9061 9815 9095
rect 9873 9061 9907 9095
rect 5641 8993 5675 9027
rect 5917 8993 5951 9027
rect 6377 8993 6411 9027
rect 7481 8993 7515 9027
rect 10425 8993 10459 9027
rect 10701 8993 10735 9027
rect 12300 8993 12334 9027
rect 2237 8925 2271 8959
rect 4169 8925 4203 8959
rect 4445 8925 4479 8959
rect 8769 8925 8803 8959
rect 2789 8857 2823 8891
rect 5733 8857 5767 8891
rect 5365 8789 5399 8823
rect 6929 8789 6963 8823
rect 8401 8789 8435 8823
rect 12403 8789 12437 8823
rect 4445 8585 4479 8619
rect 4905 8585 4939 8619
rect 6469 8585 6503 8619
rect 7941 8585 7975 8619
rect 9505 8585 9539 8619
rect 10977 8585 11011 8619
rect 6193 8517 6227 8551
rect 5273 8449 5307 8483
rect 5917 8449 5951 8483
rect 1777 8381 1811 8415
rect 3341 8381 3375 8415
rect 3525 8381 3559 8415
rect 5549 8381 5583 8415
rect 1685 8313 1719 8347
rect 2973 8313 3007 8347
rect 3846 8313 3880 8347
rect 5365 8313 5399 8347
rect 8493 8449 8527 8483
rect 9137 8449 9171 8483
rect 10333 8449 10367 8483
rect 12173 8449 12207 8483
rect 7113 8381 7147 8415
rect 7297 8381 7331 8415
rect 12484 8381 12518 8415
rect 12909 8381 12943 8415
rect 8585 8313 8619 8347
rect 10057 8313 10091 8347
rect 10149 8313 10183 8347
rect 2145 8245 2179 8279
rect 2697 8245 2731 8279
rect 6469 8245 6503 8279
rect 6561 8245 6595 8279
rect 6929 8245 6963 8279
rect 8217 8245 8251 8279
rect 9781 8245 9815 8279
rect 12587 8245 12621 8279
rect 2145 8041 2179 8075
rect 3525 8041 3559 8075
rect 3893 8041 3927 8075
rect 4261 8041 4295 8075
rect 4905 8041 4939 8075
rect 6745 8041 6779 8075
rect 7481 8041 7515 8075
rect 10793 8041 10827 8075
rect 2558 7973 2592 8007
rect 8769 7973 8803 8007
rect 10425 7973 10459 8007
rect 2237 7905 2271 7939
rect 4537 7905 4571 7939
rect 6285 7905 6319 7939
rect 6561 7905 6595 7939
rect 8125 7905 8159 7939
rect 9689 7905 9723 7939
rect 9965 7905 9999 7939
rect 11253 7905 11287 7939
rect 5457 7769 5491 7803
rect 6377 7769 6411 7803
rect 9781 7769 9815 7803
rect 1777 7701 1811 7735
rect 3157 7701 3191 7735
rect 5825 7701 5859 7735
rect 6193 7701 6227 7735
rect 11437 7701 11471 7735
rect 6009 7497 6043 7531
rect 7941 7497 7975 7531
rect 11253 7497 11287 7531
rect 6377 7429 6411 7463
rect 8217 7429 8251 7463
rect 1593 7361 1627 7395
rect 2605 7361 2639 7395
rect 3801 7361 3835 7395
rect 4537 7361 4571 7395
rect 6929 7361 6963 7395
rect 8401 7361 8435 7395
rect 8493 7293 8527 7327
rect 9689 7293 9723 7327
rect 10057 7293 10091 7327
rect 2926 7225 2960 7259
rect 4858 7225 4892 7259
rect 7021 7225 7055 7259
rect 7573 7225 7607 7259
rect 2145 7157 2179 7191
rect 2421 7157 2455 7191
rect 3525 7157 3559 7191
rect 4353 7157 4387 7191
rect 5457 7157 5491 7191
rect 10425 7157 10459 7191
rect 2237 6953 2271 6987
rect 4077 6953 4111 6987
rect 4905 6953 4939 6987
rect 6929 6953 6963 6987
rect 9505 6953 9539 6987
rect 9873 6953 9907 6987
rect 10149 6953 10183 6987
rect 10517 6953 10551 6987
rect 1547 6885 1581 6919
rect 1961 6885 1995 6919
rect 2605 6885 2639 6919
rect 5457 6885 5491 6919
rect 6377 6885 6411 6919
rect 1460 6817 1494 6851
rect 3893 6817 3927 6851
rect 7389 6817 7423 6851
rect 7481 6817 7515 6851
rect 7757 6817 7791 6851
rect 8217 6817 8251 6851
rect 9689 6817 9723 6851
rect 2513 6749 2547 6783
rect 2789 6749 2823 6783
rect 5365 6749 5399 6783
rect 3433 6681 3467 6715
rect 5917 6681 5951 6715
rect 7573 6681 7607 6715
rect 4629 6613 4663 6647
rect 9045 6613 9079 6647
rect 2513 6409 2547 6443
rect 5549 6409 5583 6443
rect 3617 6341 3651 6375
rect 4445 6341 4479 6375
rect 1961 6273 1995 6307
rect 3065 6273 3099 6307
rect 3893 6273 3927 6307
rect 10747 6273 10781 6307
rect 1685 6205 1719 6239
rect 1869 6205 1903 6239
rect 3157 6137 3191 6171
rect 4721 6205 4755 6239
rect 4997 6205 5031 6239
rect 8125 6205 8159 6239
rect 9045 6205 9079 6239
rect 9137 6205 9171 6239
rect 9321 6205 9355 6239
rect 10644 6205 10678 6239
rect 11069 6205 11103 6239
rect 8217 6137 8251 6171
rect 8493 6137 8527 6171
rect 8861 6137 8895 6171
rect 2881 6069 2915 6103
rect 3893 6069 3927 6103
rect 3985 6069 4019 6103
rect 4629 6069 4663 6103
rect 5917 6069 5951 6103
rect 6653 6069 6687 6103
rect 7389 6069 7423 6103
rect 9505 6069 9539 6103
rect 10149 6069 10183 6103
rect 1777 5865 1811 5899
rect 2329 5865 2363 5899
rect 3157 5865 3191 5899
rect 6285 5865 6319 5899
rect 7757 5865 7791 5899
rect 10149 5865 10183 5899
rect 3801 5797 3835 5831
rect 2329 5729 2363 5763
rect 2513 5729 2547 5763
rect 4077 5729 4111 5763
rect 4629 5729 4663 5763
rect 6101 5729 6135 5763
rect 7113 5729 7147 5763
rect 8401 5729 8435 5763
rect 9689 5729 9723 5763
rect 9965 5729 9999 5763
rect 4721 5661 4755 5695
rect 7481 5661 7515 5695
rect 7389 5593 7423 5627
rect 9137 5593 9171 5627
rect 9781 5593 9815 5627
rect 3433 5525 3467 5559
rect 5181 5525 5215 5559
rect 6929 5525 6963 5559
rect 7278 5525 7312 5559
rect 4261 5321 4295 5355
rect 6285 5321 6319 5355
rect 9413 5321 9447 5355
rect 9781 5321 9815 5355
rect 10977 5321 11011 5355
rect 2789 5253 2823 5287
rect 4629 5253 4663 5287
rect 6653 5253 6687 5287
rect 6929 5253 6963 5287
rect 8309 5253 8343 5287
rect 8493 5253 8527 5287
rect 10057 5253 10091 5287
rect 11345 5253 11379 5287
rect 3617 5185 3651 5219
rect 10425 5185 10459 5219
rect 1869 5117 1903 5151
rect 2237 5117 2271 5151
rect 4813 5117 4847 5151
rect 5365 5117 5399 5151
rect 5917 5117 5951 5151
rect 6837 5117 6871 5151
rect 7113 5117 7147 5151
rect 8401 5117 8435 5151
rect 8677 5117 8711 5151
rect 9965 5117 9999 5151
rect 10241 5117 10275 5151
rect 2421 5049 2455 5083
rect 3341 5049 3375 5083
rect 3433 5049 3467 5083
rect 9137 5049 9171 5083
rect 3065 4981 3099 5015
rect 4905 4981 4939 5015
rect 7297 4981 7331 5015
rect 7941 4981 7975 5015
rect 1961 4777 1995 4811
rect 2329 4777 2363 4811
rect 4721 4777 4755 4811
rect 6101 4777 6135 4811
rect 7757 4777 7791 4811
rect 9781 4777 9815 4811
rect 2605 4709 2639 4743
rect 5226 4709 5260 4743
rect 6837 4709 6871 4743
rect 7389 4709 7423 4743
rect 8769 4709 8803 4743
rect 9413 4709 9447 4743
rect 1476 4641 1510 4675
rect 4905 4641 4939 4675
rect 8217 4641 8251 4675
rect 9965 4641 9999 4675
rect 10241 4641 10275 4675
rect 11253 4641 11287 4675
rect 2513 4573 2547 4607
rect 3157 4573 3191 4607
rect 4353 4573 4387 4607
rect 6745 4573 6779 4607
rect 8033 4573 8067 4607
rect 1547 4437 1581 4471
rect 3525 4437 3559 4471
rect 5825 4437 5859 4471
rect 6561 4437 6595 4471
rect 8401 4437 8435 4471
rect 10701 4437 10735 4471
rect 11391 4437 11425 4471
rect 6193 4233 6227 4267
rect 6561 4233 6595 4267
rect 7849 4233 7883 4267
rect 8677 4233 8711 4267
rect 9781 4233 9815 4267
rect 10149 4233 10183 4267
rect 1915 4165 1949 4199
rect 10609 4165 10643 4199
rect 1685 4097 1719 4131
rect 3341 4097 3375 4131
rect 4445 4097 4479 4131
rect 6929 4097 6963 4131
rect 7205 4097 7239 4131
rect 1844 4029 1878 4063
rect 8309 4029 8343 4063
rect 8769 4029 8803 4063
rect 9965 4029 9999 4063
rect 11104 4029 11138 4063
rect 12484 4029 12518 4063
rect 12909 4029 12943 4063
rect 2329 3961 2363 3995
rect 2881 3961 2915 3995
rect 2973 3961 3007 3995
rect 4807 3961 4841 3995
rect 5641 3961 5675 3995
rect 7021 3961 7055 3995
rect 11897 3961 11931 3995
rect 2605 3893 2639 3927
rect 3801 3893 3835 3927
rect 4353 3893 4387 3927
rect 5365 3893 5399 3927
rect 11207 3893 11241 3927
rect 11529 3893 11563 3927
rect 12587 3893 12621 3927
rect 2513 3689 2547 3723
rect 4353 3689 4387 3723
rect 5733 3689 5767 3723
rect 7573 3689 7607 3723
rect 9873 3689 9907 3723
rect 10241 3689 10275 3723
rect 2053 3621 2087 3655
rect 4807 3621 4841 3655
rect 6377 3621 6411 3655
rect 7941 3621 7975 3655
rect 8585 3621 8619 3655
rect 8861 3621 8895 3655
rect 3801 3553 3835 3587
rect 10057 3553 10091 3587
rect 11161 3553 11195 3587
rect 12300 3553 12334 3587
rect 13277 3553 13311 3587
rect 2145 3485 2179 3519
rect 4445 3485 4479 3519
rect 6101 3485 6135 3519
rect 6285 3485 6319 3519
rect 7849 3485 7883 3519
rect 8585 3485 8619 3519
rect 13415 3485 13449 3519
rect 6837 3417 6871 3451
rect 8401 3417 8435 3451
rect 11345 3417 11379 3451
rect 3065 3349 3099 3383
rect 3433 3349 3467 3383
rect 5365 3349 5399 3383
rect 7205 3349 7239 3383
rect 12403 3349 12437 3383
rect 3249 3145 3283 3179
rect 3525 3145 3559 3179
rect 4721 3145 4755 3179
rect 6285 3145 6319 3179
rect 6561 3145 6595 3179
rect 7941 3145 7975 3179
rect 9873 3145 9907 3179
rect 10609 3145 10643 3179
rect 11069 3145 11103 3179
rect 12173 3145 12207 3179
rect 13599 3145 13633 3179
rect 7481 3077 7515 3111
rect 10149 3077 10183 3111
rect 11345 3077 11379 3111
rect 2329 3009 2363 3043
rect 3893 3009 3927 3043
rect 5273 3009 5307 3043
rect 5917 3009 5951 3043
rect 6929 3009 6963 3043
rect 8769 3009 8803 3043
rect 11713 3009 11747 3043
rect 4077 2941 4111 2975
rect 9965 2941 9999 2975
rect 11161 2941 11195 2975
rect 12484 2941 12518 2975
rect 12909 2941 12943 2975
rect 13528 2941 13562 2975
rect 13921 2941 13955 2975
rect 1869 2873 1903 2907
rect 2237 2873 2271 2907
rect 2691 2873 2725 2907
rect 5365 2873 5399 2907
rect 7021 2873 7055 2907
rect 8493 2873 8527 2907
rect 8585 2873 8619 2907
rect 4261 2805 4295 2839
rect 5089 2805 5123 2839
rect 8217 2805 8251 2839
rect 12587 2805 12621 2839
rect 13277 2805 13311 2839
rect 1961 2601 1995 2635
rect 7757 2601 7791 2635
rect 10057 2601 10091 2635
rect 2329 2533 2363 2567
rect 2605 2533 2639 2567
rect 3157 2533 3191 2567
rect 3893 2533 3927 2567
rect 4439 2533 4473 2567
rect 5365 2533 5399 2567
rect 5963 2533 5997 2567
rect 7113 2533 7147 2567
rect 1476 2465 1510 2499
rect 3525 2465 3559 2499
rect 4077 2465 4111 2499
rect 5860 2465 5894 2499
rect 6285 2465 6319 2499
rect 8493 2465 8527 2499
rect 9045 2465 9079 2499
rect 9873 2465 9907 2499
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 12668 2465 12702 2499
rect 13093 2465 13127 2499
rect 2513 2397 2547 2431
rect 5733 2397 5767 2431
rect 7021 2397 7055 2431
rect 8033 2397 8067 2431
rect 12771 2397 12805 2431
rect 9505 2329 9539 2363
rect 11621 2329 11655 2363
rect 1547 2261 1581 2295
rect 4997 2261 5031 2295
rect 6653 2261 6687 2295
rect 8309 2261 8343 2295
rect 8677 2261 8711 2295
<< metal1 >>
rect 6178 39760 6184 39772
rect 4126 39732 6184 39760
rect 382 39652 388 39704
rect 440 39692 446 39704
rect 4126 39692 4154 39732
rect 6178 39720 6184 39732
rect 6236 39720 6242 39772
rect 440 39664 4154 39692
rect 440 39652 446 39664
rect 5534 39652 5540 39704
rect 5592 39692 5598 39704
rect 6546 39692 6552 39704
rect 5592 39664 6552 39692
rect 5592 39652 5598 39664
rect 6546 39652 6552 39664
rect 6604 39652 6610 39704
rect 1486 39584 1492 39636
rect 1544 39624 1550 39636
rect 2130 39624 2136 39636
rect 1544 39596 2136 39624
rect 1544 39584 1550 39596
rect 2130 39584 2136 39596
rect 2188 39584 2194 39636
rect 3050 39584 3056 39636
rect 3108 39584 3114 39636
rect 3878 39584 3884 39636
rect 3936 39624 3942 39636
rect 3936 39596 4154 39624
rect 3936 39584 3942 39596
rect 3068 39488 3096 39584
rect 4126 39556 4154 39596
rect 5074 39584 5080 39636
rect 5132 39624 5138 39636
rect 5718 39624 5724 39636
rect 5132 39596 5724 39624
rect 5132 39584 5138 39596
rect 5718 39584 5724 39596
rect 5776 39584 5782 39636
rect 7466 39584 7472 39636
rect 7524 39624 7530 39636
rect 8018 39624 8024 39636
rect 7524 39596 8024 39624
rect 7524 39584 7530 39596
rect 8018 39584 8024 39596
rect 8076 39584 8082 39636
rect 13814 39584 13820 39636
rect 13872 39624 13878 39636
rect 15470 39624 15476 39636
rect 13872 39596 15476 39624
rect 13872 39584 13878 39596
rect 15470 39584 15476 39596
rect 15528 39584 15534 39636
rect 9398 39556 9404 39568
rect 4126 39528 9404 39556
rect 9398 39516 9404 39528
rect 9456 39516 9462 39568
rect 5810 39488 5816 39500
rect 3068 39460 5816 39488
rect 5810 39448 5816 39460
rect 5868 39448 5874 39500
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 7837 35275 7895 35281
rect 7837 35241 7849 35275
rect 7883 35272 7895 35275
rect 8110 35272 8116 35284
rect 7883 35244 8116 35272
rect 7883 35241 7895 35244
rect 7837 35235 7895 35241
rect 8110 35232 8116 35244
rect 8168 35232 8174 35284
rect 7650 35136 7656 35148
rect 7611 35108 7656 35136
rect 7650 35096 7656 35108
rect 7708 35096 7714 35148
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 8481 34731 8539 34737
rect 8481 34697 8493 34731
rect 8527 34728 8539 34731
rect 9766 34728 9772 34740
rect 8527 34700 9772 34728
rect 8527 34697 8539 34700
rect 8481 34691 8539 34697
rect 9766 34688 9772 34700
rect 9824 34688 9830 34740
rect 9861 34731 9919 34737
rect 9861 34697 9873 34731
rect 9907 34728 9919 34731
rect 10686 34728 10692 34740
rect 9907 34700 10692 34728
rect 9907 34697 9919 34700
rect 9861 34691 9919 34697
rect 10686 34688 10692 34700
rect 10744 34688 10750 34740
rect 13357 34731 13415 34737
rect 13357 34697 13369 34731
rect 13403 34728 13415 34731
rect 14642 34728 14648 34740
rect 13403 34700 14648 34728
rect 13403 34697 13415 34700
rect 13357 34691 13415 34697
rect 14642 34688 14648 34700
rect 14700 34688 14706 34740
rect 4709 34663 4767 34669
rect 4709 34629 4721 34663
rect 4755 34660 4767 34663
rect 7009 34663 7067 34669
rect 4755 34632 6868 34660
rect 4755 34629 4767 34632
rect 4709 34623 4767 34629
rect 4614 34552 4620 34604
rect 4672 34592 4678 34604
rect 6549 34595 6607 34601
rect 6549 34592 6561 34595
rect 4672 34564 6561 34592
rect 4672 34552 4678 34564
rect 6549 34561 6561 34564
rect 6595 34561 6607 34595
rect 6840 34592 6868 34632
rect 7009 34629 7021 34663
rect 7055 34660 7067 34663
rect 13446 34660 13452 34672
rect 7055 34632 13452 34660
rect 7055 34629 7067 34632
rect 7009 34623 7067 34629
rect 13446 34620 13452 34632
rect 13504 34620 13510 34672
rect 12526 34592 12532 34604
rect 6840 34564 12532 34592
rect 6549 34555 6607 34561
rect 4525 34527 4583 34533
rect 4525 34493 4537 34527
rect 4571 34524 4583 34527
rect 6564 34524 6592 34555
rect 12526 34552 12532 34564
rect 12584 34552 12590 34604
rect 6825 34527 6883 34533
rect 6825 34524 6837 34527
rect 4571 34496 5212 34524
rect 6564 34496 6837 34524
rect 4571 34493 4583 34496
rect 4525 34487 4583 34493
rect 5184 34397 5212 34496
rect 6825 34493 6837 34496
rect 6871 34493 6883 34527
rect 8294 34524 8300 34536
rect 8255 34496 8300 34524
rect 6825 34487 6883 34493
rect 8294 34484 8300 34496
rect 8352 34524 8358 34536
rect 8849 34527 8907 34533
rect 8849 34524 8861 34527
rect 8352 34496 8861 34524
rect 8352 34484 8358 34496
rect 8849 34493 8861 34496
rect 8895 34493 8907 34527
rect 8849 34487 8907 34493
rect 9306 34484 9312 34536
rect 9364 34524 9370 34536
rect 9677 34527 9735 34533
rect 9677 34524 9689 34527
rect 9364 34496 9689 34524
rect 9364 34484 9370 34496
rect 9677 34493 9689 34496
rect 9723 34524 9735 34527
rect 10229 34527 10287 34533
rect 10229 34524 10241 34527
rect 9723 34496 10241 34524
rect 9723 34493 9735 34496
rect 9677 34487 9735 34493
rect 10229 34493 10241 34496
rect 10275 34493 10287 34527
rect 10229 34487 10287 34493
rect 11974 34484 11980 34536
rect 12032 34524 12038 34536
rect 13173 34527 13231 34533
rect 13173 34524 13185 34527
rect 12032 34496 13185 34524
rect 12032 34484 12038 34496
rect 13173 34493 13185 34496
rect 13219 34524 13231 34527
rect 13725 34527 13783 34533
rect 13725 34524 13737 34527
rect 13219 34496 13737 34524
rect 13219 34493 13231 34496
rect 13173 34487 13231 34493
rect 13725 34493 13737 34496
rect 13771 34493 13783 34527
rect 13725 34487 13783 34493
rect 5169 34391 5227 34397
rect 5169 34357 5181 34391
rect 5215 34388 5227 34391
rect 5258 34388 5264 34400
rect 5215 34360 5264 34388
rect 5215 34357 5227 34360
rect 5169 34351 5227 34357
rect 5258 34348 5264 34360
rect 5316 34348 5322 34400
rect 7650 34348 7656 34400
rect 7708 34388 7714 34400
rect 7745 34391 7803 34397
rect 7745 34388 7757 34391
rect 7708 34360 7757 34388
rect 7708 34348 7714 34360
rect 7745 34357 7757 34360
rect 7791 34388 7803 34391
rect 10502 34388 10508 34400
rect 7791 34360 10508 34388
rect 7791 34357 7803 34360
rect 7745 34351 7803 34357
rect 10502 34348 10508 34360
rect 10560 34348 10566 34400
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 8297 34187 8355 34193
rect 8297 34153 8309 34187
rect 8343 34184 8355 34187
rect 8846 34184 8852 34196
rect 8343 34156 8852 34184
rect 8343 34153 8355 34156
rect 8297 34147 8355 34153
rect 8846 34144 8852 34156
rect 8904 34144 8910 34196
rect 8110 34048 8116 34060
rect 8071 34020 8116 34048
rect 8110 34008 8116 34020
rect 8168 34008 8174 34060
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 5626 33260 5632 33312
rect 5684 33300 5690 33312
rect 8110 33300 8116 33312
rect 5684 33272 8116 33300
rect 5684 33260 5690 33272
rect 8110 33260 8116 33272
rect 8168 33260 8174 33312
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 1026 30336 1032 30388
rect 1084 30376 1090 30388
rect 1535 30379 1593 30385
rect 1535 30376 1547 30379
rect 1084 30348 1547 30376
rect 1084 30336 1090 30348
rect 1535 30345 1547 30348
rect 1581 30345 1593 30379
rect 1535 30339 1593 30345
rect 1464 30175 1522 30181
rect 1464 30141 1476 30175
rect 1510 30172 1522 30175
rect 1510 30144 1992 30172
rect 1510 30141 1522 30144
rect 1464 30135 1522 30141
rect 1964 30045 1992 30144
rect 1949 30039 2007 30045
rect 1949 30005 1961 30039
rect 1995 30036 2007 30039
rect 3142 30036 3148 30048
rect 1995 30008 3148 30036
rect 1995 30005 2007 30008
rect 1949 29999 2007 30005
rect 3142 29996 3148 30008
rect 3200 29996 3206 30048
rect 7285 30039 7343 30045
rect 7285 30005 7297 30039
rect 7331 30036 7343 30039
rect 10042 30036 10048 30048
rect 7331 30008 10048 30036
rect 7331 30005 7343 30008
rect 7285 29999 7343 30005
rect 10042 29996 10048 30008
rect 10100 29996 10106 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 7098 29792 7104 29844
rect 7156 29832 7162 29844
rect 7607 29835 7665 29841
rect 7607 29832 7619 29835
rect 7156 29804 7619 29832
rect 7156 29792 7162 29804
rect 7607 29801 7619 29804
rect 7653 29801 7665 29835
rect 7607 29795 7665 29801
rect 6086 29764 6092 29776
rect 6047 29736 6092 29764
rect 6086 29724 6092 29736
rect 6144 29724 6150 29776
rect 7536 29699 7594 29705
rect 7536 29665 7548 29699
rect 7582 29696 7594 29699
rect 7834 29696 7840 29708
rect 7582 29668 7840 29696
rect 7582 29665 7594 29668
rect 7536 29659 7594 29665
rect 7834 29656 7840 29668
rect 7892 29656 7898 29708
rect 5994 29628 6000 29640
rect 5955 29600 6000 29628
rect 5994 29588 6000 29600
rect 6052 29588 6058 29640
rect 6641 29631 6699 29637
rect 6641 29597 6653 29631
rect 6687 29628 6699 29631
rect 7190 29628 7196 29640
rect 6687 29600 7196 29628
rect 6687 29597 6699 29600
rect 6641 29591 6699 29597
rect 7190 29588 7196 29600
rect 7248 29588 7254 29640
rect 6270 29452 6276 29504
rect 6328 29492 6334 29504
rect 8294 29492 8300 29504
rect 6328 29464 8300 29492
rect 6328 29452 6334 29464
rect 8294 29452 8300 29464
rect 8352 29452 8358 29504
rect 8478 29492 8484 29504
rect 8439 29464 8484 29492
rect 8478 29452 8484 29464
rect 8536 29452 8542 29504
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 5902 29248 5908 29300
rect 5960 29288 5966 29300
rect 6270 29288 6276 29300
rect 5960 29260 6276 29288
rect 5960 29248 5966 29260
rect 6270 29248 6276 29260
rect 6328 29248 6334 29300
rect 7834 29288 7840 29300
rect 7795 29260 7840 29288
rect 7834 29248 7840 29260
rect 7892 29248 7898 29300
rect 6178 29180 6184 29232
rect 6236 29220 6242 29232
rect 7098 29220 7104 29232
rect 6236 29192 7104 29220
rect 6236 29180 6242 29192
rect 7098 29180 7104 29192
rect 7156 29180 7162 29232
rect 4847 29155 4905 29161
rect 4847 29121 4859 29155
rect 4893 29152 4905 29155
rect 7282 29152 7288 29164
rect 4893 29124 7288 29152
rect 4893 29121 4905 29124
rect 4847 29115 4905 29121
rect 7282 29112 7288 29124
rect 7340 29112 7346 29164
rect 7852 29152 7880 29248
rect 8757 29155 8815 29161
rect 8757 29152 8769 29155
rect 7852 29124 8769 29152
rect 8757 29121 8769 29124
rect 8803 29152 8815 29155
rect 10594 29152 10600 29164
rect 8803 29124 10600 29152
rect 8803 29121 8815 29124
rect 8757 29115 8815 29121
rect 10594 29112 10600 29124
rect 10652 29112 10658 29164
rect 4760 29087 4818 29093
rect 4760 29053 4772 29087
rect 4806 29084 4818 29087
rect 5772 29087 5830 29093
rect 4806 29056 5120 29084
rect 4806 29053 4818 29056
rect 4760 29047 4818 29053
rect 5092 28960 5120 29056
rect 5772 29053 5784 29087
rect 5818 29084 5830 29087
rect 6270 29084 6276 29096
rect 5818 29056 6276 29084
rect 5818 29053 5830 29056
rect 5772 29047 5830 29053
rect 6270 29044 6276 29056
rect 6328 29044 6334 29096
rect 5859 29019 5917 29025
rect 5859 28985 5871 29019
rect 5905 29016 5917 29019
rect 6914 29016 6920 29028
rect 5905 28988 6920 29016
rect 5905 28985 5917 28988
rect 5859 28979 5917 28985
rect 6914 28976 6920 28988
rect 6972 28976 6978 29028
rect 7009 29019 7067 29025
rect 7009 28985 7021 29019
rect 7055 28985 7067 29019
rect 7009 28979 7067 28985
rect 5074 28908 5080 28960
rect 5132 28948 5138 28960
rect 5169 28951 5227 28957
rect 5169 28948 5181 28951
rect 5132 28920 5181 28948
rect 5132 28908 5138 28920
rect 5169 28917 5181 28920
rect 5215 28917 5227 28951
rect 5169 28911 5227 28917
rect 5629 28951 5687 28957
rect 5629 28917 5641 28951
rect 5675 28948 5687 28951
rect 6086 28948 6092 28960
rect 5675 28920 6092 28948
rect 5675 28917 5687 28920
rect 5629 28911 5687 28917
rect 6086 28908 6092 28920
rect 6144 28908 6150 28960
rect 6638 28948 6644 28960
rect 6599 28920 6644 28948
rect 6638 28908 6644 28920
rect 6696 28948 6702 28960
rect 7024 28948 7052 28979
rect 7190 28976 7196 29028
rect 7248 29016 7254 29028
rect 7561 29019 7619 29025
rect 7561 29016 7573 29019
rect 7248 28988 7573 29016
rect 7248 28976 7254 28988
rect 7561 28985 7573 28988
rect 7607 28985 7619 29019
rect 8478 29016 8484 29028
rect 8439 28988 8484 29016
rect 7561 28979 7619 28985
rect 8478 28976 8484 28988
rect 8536 28976 8542 29028
rect 8570 28976 8576 29028
rect 8628 29016 8634 29028
rect 8628 28988 8673 29016
rect 8628 28976 8634 28988
rect 7650 28948 7656 28960
rect 6696 28920 7656 28948
rect 6696 28908 6702 28920
rect 7650 28908 7656 28920
rect 7708 28908 7714 28960
rect 8297 28951 8355 28957
rect 8297 28917 8309 28951
rect 8343 28948 8355 28951
rect 8588 28948 8616 28976
rect 8343 28920 8616 28948
rect 8343 28917 8355 28920
rect 8297 28911 8355 28917
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 5031 28747 5089 28753
rect 5031 28713 5043 28747
rect 5077 28744 5089 28747
rect 5813 28747 5871 28753
rect 5813 28744 5825 28747
rect 5077 28716 5825 28744
rect 5077 28713 5089 28716
rect 5031 28707 5089 28713
rect 5813 28713 5825 28716
rect 5859 28744 5871 28747
rect 5994 28744 6000 28756
rect 5859 28716 6000 28744
rect 5859 28713 5871 28716
rect 5813 28707 5871 28713
rect 5994 28704 6000 28716
rect 6052 28704 6058 28756
rect 6914 28744 6920 28756
rect 6875 28716 6920 28744
rect 6914 28704 6920 28716
rect 6972 28704 6978 28756
rect 7282 28744 7288 28756
rect 7243 28716 7288 28744
rect 7282 28704 7288 28716
rect 7340 28744 7346 28756
rect 7340 28716 7604 28744
rect 7340 28704 7346 28716
rect 6086 28676 6092 28688
rect 6047 28648 6092 28676
rect 6086 28636 6092 28648
rect 6144 28636 6150 28688
rect 7576 28685 7604 28716
rect 7561 28679 7619 28685
rect 7561 28645 7573 28679
rect 7607 28645 7619 28679
rect 7561 28639 7619 28645
rect 7650 28636 7656 28688
rect 7708 28676 7714 28688
rect 7708 28648 7753 28676
rect 7708 28636 7714 28648
rect 1486 28568 1492 28620
rect 1544 28608 1550 28620
rect 4982 28617 4988 28620
rect 4928 28611 4988 28617
rect 4928 28608 4940 28611
rect 1544 28580 4940 28608
rect 1544 28568 1550 28580
rect 4928 28577 4940 28580
rect 4974 28577 4988 28611
rect 4928 28571 4988 28577
rect 4982 28568 4988 28571
rect 5040 28568 5046 28620
rect 9582 28608 9588 28620
rect 9543 28580 9588 28608
rect 9582 28568 9588 28580
rect 9640 28568 9646 28620
rect 4430 28500 4436 28552
rect 4488 28540 4494 28552
rect 5994 28540 6000 28552
rect 4488 28512 6000 28540
rect 4488 28500 4494 28512
rect 5994 28500 6000 28512
rect 6052 28500 6058 28552
rect 6641 28543 6699 28549
rect 6641 28509 6653 28543
rect 6687 28540 6699 28543
rect 7006 28540 7012 28552
rect 6687 28512 7012 28540
rect 6687 28509 6699 28512
rect 6641 28503 6699 28509
rect 7006 28500 7012 28512
rect 7064 28540 7070 28552
rect 7837 28543 7895 28549
rect 7837 28540 7849 28543
rect 7064 28512 7849 28540
rect 7064 28500 7070 28512
rect 7837 28509 7849 28512
rect 7883 28509 7895 28543
rect 7837 28503 7895 28509
rect 5350 28404 5356 28416
rect 5311 28376 5356 28404
rect 5350 28364 5356 28376
rect 5408 28364 5414 28416
rect 8202 28364 8208 28416
rect 8260 28404 8266 28416
rect 9306 28404 9312 28416
rect 8260 28376 9312 28404
rect 8260 28364 8266 28376
rect 9306 28364 9312 28376
rect 9364 28364 9370 28416
rect 9674 28364 9680 28416
rect 9732 28404 9738 28416
rect 9815 28407 9873 28413
rect 9815 28404 9827 28407
rect 9732 28376 9827 28404
rect 9732 28364 9738 28376
rect 9815 28373 9827 28376
rect 9861 28373 9873 28407
rect 9815 28367 9873 28373
rect 10321 28407 10379 28413
rect 10321 28373 10333 28407
rect 10367 28404 10379 28407
rect 10410 28404 10416 28416
rect 10367 28376 10416 28404
rect 10367 28373 10379 28376
rect 10321 28367 10379 28373
rect 10410 28364 10416 28376
rect 10468 28364 10474 28416
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 3283 28203 3341 28209
rect 3283 28169 3295 28203
rect 3329 28200 3341 28203
rect 4430 28200 4436 28212
rect 3329 28172 4436 28200
rect 3329 28169 3341 28172
rect 3283 28163 3341 28169
rect 4430 28160 4436 28172
rect 4488 28160 4494 28212
rect 4614 28200 4620 28212
rect 4575 28172 4620 28200
rect 4614 28160 4620 28172
rect 4672 28160 4678 28212
rect 4982 28200 4988 28212
rect 4943 28172 4988 28200
rect 4982 28160 4988 28172
rect 5040 28160 5046 28212
rect 7650 28160 7656 28212
rect 7708 28200 7714 28212
rect 8113 28203 8171 28209
rect 8113 28200 8125 28203
rect 7708 28172 8125 28200
rect 7708 28160 7714 28172
rect 8113 28169 8125 28172
rect 8159 28169 8171 28203
rect 10042 28200 10048 28212
rect 10003 28172 10048 28200
rect 8113 28163 8171 28169
rect 10042 28160 10048 28172
rect 10100 28160 10106 28212
rect 3697 28135 3755 28141
rect 3697 28101 3709 28135
rect 3743 28132 3755 28135
rect 3970 28132 3976 28144
rect 3743 28104 3976 28132
rect 3743 28101 3755 28104
rect 3697 28095 3755 28101
rect 3212 27999 3270 28005
rect 3212 27965 3224 27999
rect 3258 27996 3270 27999
rect 3712 27996 3740 28095
rect 3970 28092 3976 28104
rect 4028 28092 4034 28144
rect 5534 28092 5540 28144
rect 5592 28132 5598 28144
rect 5718 28132 5724 28144
rect 5592 28104 5724 28132
rect 5592 28092 5598 28104
rect 5718 28092 5724 28104
rect 5776 28092 5782 28144
rect 7837 28135 7895 28141
rect 7837 28101 7849 28135
rect 7883 28132 7895 28135
rect 10410 28132 10416 28144
rect 7883 28104 10416 28132
rect 7883 28101 7895 28104
rect 7837 28095 7895 28101
rect 10410 28092 10416 28104
rect 10468 28092 10474 28144
rect 10042 28024 10048 28076
rect 10100 28064 10106 28076
rect 10321 28067 10379 28073
rect 10321 28064 10333 28067
rect 10100 28036 10333 28064
rect 10100 28024 10106 28036
rect 10321 28033 10333 28036
rect 10367 28033 10379 28067
rect 10594 28064 10600 28076
rect 10555 28036 10600 28064
rect 10321 28027 10379 28033
rect 10594 28024 10600 28036
rect 10652 28024 10658 28076
rect 3258 27968 3740 27996
rect 4203 27999 4261 28005
rect 3258 27965 3270 27968
rect 3212 27959 3270 27965
rect 4203 27965 4215 27999
rect 4249 27965 4261 27999
rect 6914 27996 6920 28008
rect 6875 27968 6920 27996
rect 4203 27959 4261 27965
rect 3326 27888 3332 27940
rect 3384 27928 3390 27940
rect 4218 27928 4246 27959
rect 6914 27956 6920 27968
rect 6972 27956 6978 28008
rect 4614 27928 4620 27940
rect 3384 27900 4620 27928
rect 3384 27888 3390 27900
rect 4614 27888 4620 27900
rect 4672 27888 4678 27940
rect 4982 27888 4988 27940
rect 5040 27928 5046 27940
rect 5261 27931 5319 27937
rect 5261 27928 5273 27931
rect 5040 27900 5273 27928
rect 5040 27888 5046 27900
rect 5261 27897 5273 27900
rect 5307 27897 5319 27931
rect 5261 27891 5319 27897
rect 5350 27888 5356 27940
rect 5408 27928 5414 27940
rect 5905 27931 5963 27937
rect 5408 27900 5453 27928
rect 5408 27888 5414 27900
rect 5905 27897 5917 27931
rect 5951 27928 5963 27931
rect 7006 27928 7012 27940
rect 5951 27900 7012 27928
rect 5951 27897 5963 27900
rect 5905 27891 5963 27897
rect 7006 27888 7012 27900
rect 7064 27888 7070 27940
rect 7238 27931 7296 27937
rect 7238 27897 7250 27931
rect 7284 27897 7296 27931
rect 8754 27928 8760 27940
rect 8715 27900 8760 27928
rect 7238 27891 7296 27897
rect 4295 27863 4353 27869
rect 4295 27829 4307 27863
rect 4341 27860 4353 27863
rect 5534 27860 5540 27872
rect 4341 27832 5540 27860
rect 4341 27829 4353 27832
rect 4295 27823 4353 27829
rect 5534 27820 5540 27832
rect 5592 27820 5598 27872
rect 6086 27820 6092 27872
rect 6144 27860 6150 27872
rect 6181 27863 6239 27869
rect 6181 27860 6193 27863
rect 6144 27832 6193 27860
rect 6144 27820 6150 27832
rect 6181 27829 6193 27832
rect 6227 27829 6239 27863
rect 6181 27823 6239 27829
rect 6641 27863 6699 27869
rect 6641 27829 6653 27863
rect 6687 27860 6699 27863
rect 6730 27860 6736 27872
rect 6687 27832 6736 27860
rect 6687 27829 6699 27832
rect 6641 27823 6699 27829
rect 6730 27820 6736 27832
rect 6788 27860 6794 27872
rect 7253 27860 7281 27891
rect 8754 27888 8760 27900
rect 8812 27888 8818 27940
rect 8849 27931 8907 27937
rect 8849 27897 8861 27931
rect 8895 27897 8907 27931
rect 9398 27928 9404 27940
rect 9359 27900 9404 27928
rect 8849 27891 8907 27897
rect 6788 27832 7281 27860
rect 6788 27820 6794 27832
rect 8294 27820 8300 27872
rect 8352 27860 8358 27872
rect 8573 27863 8631 27869
rect 8573 27860 8585 27863
rect 8352 27832 8585 27860
rect 8352 27820 8358 27832
rect 8573 27829 8585 27832
rect 8619 27860 8631 27863
rect 8864 27860 8892 27891
rect 9398 27888 9404 27900
rect 9456 27888 9462 27940
rect 9858 27928 9864 27940
rect 9508 27900 9864 27928
rect 9508 27860 9536 27900
rect 9858 27888 9864 27900
rect 9916 27888 9922 27940
rect 10410 27888 10416 27940
rect 10468 27928 10474 27940
rect 10468 27900 10513 27928
rect 10468 27888 10474 27900
rect 8619 27832 9536 27860
rect 8619 27829 8631 27832
rect 8573 27823 8631 27829
rect 9582 27820 9588 27872
rect 9640 27860 9646 27872
rect 9769 27863 9827 27869
rect 9769 27860 9781 27863
rect 9640 27832 9781 27860
rect 9640 27820 9646 27832
rect 9769 27829 9781 27832
rect 9815 27860 9827 27863
rect 12066 27860 12072 27872
rect 9815 27832 12072 27860
rect 9815 27829 9827 27832
rect 9769 27823 9827 27829
rect 12066 27820 12072 27832
rect 12124 27820 12130 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 4982 27656 4988 27668
rect 4943 27628 4988 27656
rect 4982 27616 4988 27628
rect 5040 27616 5046 27668
rect 5994 27616 6000 27668
rect 6052 27656 6058 27668
rect 6273 27659 6331 27665
rect 6273 27656 6285 27659
rect 6052 27628 6285 27656
rect 6052 27616 6058 27628
rect 6273 27625 6285 27628
rect 6319 27625 6331 27659
rect 8294 27656 8300 27668
rect 8255 27628 8300 27656
rect 6273 27619 6331 27625
rect 8294 27616 8300 27628
rect 8352 27616 8358 27668
rect 9674 27616 9680 27668
rect 9732 27656 9738 27668
rect 9732 27628 9812 27656
rect 9732 27616 9738 27628
rect 5166 27548 5172 27600
rect 5224 27588 5230 27600
rect 5398 27591 5456 27597
rect 5398 27588 5410 27591
rect 5224 27560 5410 27588
rect 5224 27548 5230 27560
rect 5398 27557 5410 27560
rect 5444 27557 5456 27591
rect 5398 27551 5456 27557
rect 7739 27591 7797 27597
rect 7739 27557 7751 27591
rect 7785 27588 7797 27591
rect 8110 27588 8116 27600
rect 7785 27560 8116 27588
rect 7785 27557 7797 27560
rect 7739 27551 7797 27557
rect 8110 27548 8116 27560
rect 8168 27548 8174 27600
rect 9784 27597 9812 27628
rect 9769 27591 9827 27597
rect 9769 27557 9781 27591
rect 9815 27557 9827 27591
rect 9769 27551 9827 27557
rect 9858 27548 9864 27600
rect 9916 27588 9922 27600
rect 9916 27560 9961 27588
rect 9916 27548 9922 27560
rect 3012 27523 3070 27529
rect 3012 27489 3024 27523
rect 3058 27520 3070 27523
rect 3234 27520 3240 27532
rect 3058 27492 3240 27520
rect 3058 27489 3070 27492
rect 3012 27483 3070 27489
rect 3234 27480 3240 27492
rect 3292 27480 3298 27532
rect 4132 27523 4190 27529
rect 4132 27489 4144 27523
rect 4178 27520 4190 27523
rect 4338 27520 4344 27532
rect 4178 27492 4344 27520
rect 4178 27489 4190 27492
rect 4132 27483 4190 27489
rect 4338 27480 4344 27492
rect 4396 27480 4402 27532
rect 5997 27523 6055 27529
rect 5997 27489 6009 27523
rect 6043 27520 6055 27523
rect 6638 27520 6644 27532
rect 6043 27492 6644 27520
rect 6043 27489 6055 27492
rect 5997 27483 6055 27489
rect 6638 27480 6644 27492
rect 6696 27480 6702 27532
rect 10502 27480 10508 27532
rect 10560 27520 10566 27532
rect 11238 27520 11244 27532
rect 11296 27529 11302 27532
rect 11296 27523 11334 27529
rect 10560 27492 11244 27520
rect 10560 27480 10566 27492
rect 11238 27480 11244 27492
rect 11322 27489 11334 27523
rect 11296 27483 11334 27489
rect 11296 27480 11302 27483
rect 3099 27455 3157 27461
rect 3099 27421 3111 27455
rect 3145 27452 3157 27455
rect 4982 27452 4988 27464
rect 3145 27424 4988 27452
rect 3145 27421 3157 27424
rect 3099 27415 3157 27421
rect 4982 27412 4988 27424
rect 5040 27412 5046 27464
rect 5077 27455 5135 27461
rect 5077 27421 5089 27455
rect 5123 27421 5135 27455
rect 7374 27452 7380 27464
rect 7335 27424 7380 27452
rect 5077 27415 5135 27421
rect 2958 27344 2964 27396
rect 3016 27384 3022 27396
rect 5092 27384 5120 27415
rect 7374 27412 7380 27424
rect 7432 27412 7438 27464
rect 8754 27452 8760 27464
rect 8667 27424 8760 27452
rect 8754 27412 8760 27424
rect 8812 27452 8818 27464
rect 11379 27455 11437 27461
rect 11379 27452 11391 27455
rect 8812 27424 11391 27452
rect 8812 27412 8818 27424
rect 11379 27421 11391 27424
rect 11425 27421 11437 27455
rect 11379 27415 11437 27421
rect 6178 27384 6184 27396
rect 3016 27356 6184 27384
rect 3016 27344 3022 27356
rect 6178 27344 6184 27356
rect 6236 27344 6242 27396
rect 8478 27344 8484 27396
rect 8536 27384 8542 27396
rect 9950 27384 9956 27396
rect 8536 27356 9956 27384
rect 8536 27344 8542 27356
rect 9950 27344 9956 27356
rect 10008 27384 10014 27396
rect 10321 27387 10379 27393
rect 10321 27384 10333 27387
rect 10008 27356 10333 27384
rect 10008 27344 10014 27356
rect 10321 27353 10333 27356
rect 10367 27353 10379 27387
rect 10321 27347 10379 27353
rect 3510 27316 3516 27328
rect 3471 27288 3516 27316
rect 3510 27276 3516 27288
rect 3568 27276 3574 27328
rect 4062 27276 4068 27328
rect 4120 27316 4126 27328
rect 4203 27319 4261 27325
rect 4203 27316 4215 27319
rect 4120 27288 4215 27316
rect 4120 27276 4126 27288
rect 4203 27285 4215 27288
rect 4249 27285 4261 27319
rect 4203 27279 4261 27285
rect 6914 27276 6920 27328
rect 6972 27316 6978 27328
rect 7009 27319 7067 27325
rect 7009 27316 7021 27319
rect 6972 27288 7021 27316
rect 6972 27276 6978 27288
rect 7009 27285 7021 27288
rect 7055 27316 7067 27319
rect 7558 27316 7564 27328
rect 7055 27288 7564 27316
rect 7055 27285 7067 27288
rect 7009 27279 7067 27285
rect 7558 27276 7564 27288
rect 7616 27276 7622 27328
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 3234 27112 3240 27124
rect 3195 27084 3240 27112
rect 3234 27072 3240 27084
rect 3292 27112 3298 27124
rect 3292 27084 4154 27112
rect 3292 27072 3298 27084
rect 4126 27044 4154 27084
rect 4338 27072 4344 27124
rect 4396 27112 4402 27124
rect 4433 27115 4491 27121
rect 4433 27112 4445 27115
rect 4396 27084 4445 27112
rect 4396 27072 4402 27084
rect 4433 27081 4445 27084
rect 4479 27081 4491 27115
rect 4433 27075 4491 27081
rect 5905 27115 5963 27121
rect 5905 27081 5917 27115
rect 5951 27112 5963 27115
rect 6086 27112 6092 27124
rect 5951 27084 6092 27112
rect 5951 27081 5963 27084
rect 5905 27075 5963 27081
rect 6086 27072 6092 27084
rect 6144 27072 6150 27124
rect 9858 27072 9864 27124
rect 9916 27112 9922 27124
rect 10321 27115 10379 27121
rect 10321 27112 10333 27115
rect 9916 27084 10333 27112
rect 9916 27072 9922 27084
rect 10321 27081 10333 27084
rect 10367 27081 10379 27115
rect 11238 27112 11244 27124
rect 11199 27084 11244 27112
rect 10321 27075 10379 27081
rect 11238 27072 11244 27084
rect 11296 27112 11302 27124
rect 12342 27112 12348 27124
rect 11296 27084 12348 27112
rect 11296 27072 11302 27084
rect 12342 27072 12348 27084
rect 12400 27072 12406 27124
rect 5718 27044 5724 27056
rect 4126 27016 5724 27044
rect 5718 27004 5724 27016
rect 5776 27044 5782 27056
rect 10410 27044 10416 27056
rect 5776 27016 10416 27044
rect 5776 27004 5782 27016
rect 10410 27004 10416 27016
rect 10468 27004 10474 27056
rect 3510 26976 3516 26988
rect 3471 26948 3516 26976
rect 3510 26936 3516 26948
rect 3568 26936 3574 26988
rect 6178 26976 6184 26988
rect 6139 26948 6184 26976
rect 6178 26936 6184 26948
rect 6236 26936 6242 26988
rect 6730 26936 6736 26988
rect 6788 26976 6794 26988
rect 7101 26979 7159 26985
rect 7101 26976 7113 26979
rect 6788 26948 7113 26976
rect 6788 26936 6794 26948
rect 7101 26945 7113 26948
rect 7147 26976 7159 26979
rect 7377 26979 7435 26985
rect 7377 26976 7389 26979
rect 7147 26948 7389 26976
rect 7147 26945 7159 26948
rect 7101 26939 7159 26945
rect 7377 26945 7389 26948
rect 7423 26976 7435 26979
rect 8110 26976 8116 26988
rect 7423 26948 8116 26976
rect 7423 26945 7435 26948
rect 7377 26939 7435 26945
rect 2476 26911 2534 26917
rect 2476 26877 2488 26911
rect 2522 26908 2534 26911
rect 4985 26911 5043 26917
rect 2522 26880 3004 26908
rect 2522 26877 2534 26880
rect 2476 26871 2534 26877
rect 2406 26732 2412 26784
rect 2464 26772 2470 26784
rect 2976 26781 3004 26880
rect 4985 26877 4997 26911
rect 5031 26908 5043 26911
rect 7561 26911 7619 26917
rect 5031 26880 6684 26908
rect 5031 26877 5043 26880
rect 4985 26871 5043 26877
rect 3602 26840 3608 26852
rect 3563 26812 3608 26840
rect 3602 26800 3608 26812
rect 3660 26800 3666 26852
rect 4157 26843 4215 26849
rect 4157 26809 4169 26843
rect 4203 26840 4215 26843
rect 4890 26840 4896 26852
rect 4203 26812 4896 26840
rect 4203 26809 4215 26812
rect 4157 26803 4215 26809
rect 4890 26800 4896 26812
rect 4948 26800 4954 26852
rect 5166 26840 5172 26852
rect 5000 26812 5172 26840
rect 5000 26784 5028 26812
rect 5166 26800 5172 26812
rect 5224 26840 5230 26852
rect 5306 26843 5364 26849
rect 5306 26840 5318 26843
rect 5224 26812 5318 26840
rect 5224 26800 5230 26812
rect 5306 26809 5318 26812
rect 5352 26809 5364 26843
rect 5306 26803 5364 26809
rect 2547 26775 2605 26781
rect 2547 26772 2559 26775
rect 2464 26744 2559 26772
rect 2464 26732 2470 26744
rect 2547 26741 2559 26744
rect 2593 26741 2605 26775
rect 2547 26735 2605 26741
rect 2961 26775 3019 26781
rect 2961 26741 2973 26775
rect 3007 26772 3019 26775
rect 3326 26772 3332 26784
rect 3007 26744 3332 26772
rect 3007 26741 3019 26744
rect 2961 26735 3019 26741
rect 3326 26732 3332 26744
rect 3384 26732 3390 26784
rect 4801 26775 4859 26781
rect 4801 26741 4813 26775
rect 4847 26772 4859 26775
rect 4982 26772 4988 26784
rect 4847 26744 4988 26772
rect 4847 26741 4859 26744
rect 4801 26735 4859 26741
rect 4982 26732 4988 26744
rect 5040 26732 5046 26784
rect 6656 26781 6684 26880
rect 7561 26877 7573 26911
rect 7607 26908 7619 26911
rect 7607 26880 7788 26908
rect 7607 26877 7619 26880
rect 7561 26871 7619 26877
rect 6641 26775 6699 26781
rect 6641 26741 6653 26775
rect 6687 26772 6699 26775
rect 6914 26772 6920 26784
rect 6687 26744 6920 26772
rect 6687 26741 6699 26744
rect 6641 26735 6699 26741
rect 6914 26732 6920 26744
rect 6972 26732 6978 26784
rect 7760 26772 7788 26880
rect 7897 26849 7925 26948
rect 8110 26936 8116 26948
rect 8168 26936 8174 26988
rect 10045 26979 10103 26985
rect 10045 26945 10057 26979
rect 10091 26976 10103 26979
rect 10594 26976 10600 26988
rect 10091 26948 10600 26976
rect 10091 26945 10103 26948
rect 10045 26939 10103 26945
rect 10594 26936 10600 26948
rect 10652 26936 10658 26988
rect 8481 26911 8539 26917
rect 8481 26877 8493 26911
rect 8527 26908 8539 26911
rect 9125 26911 9183 26917
rect 9125 26908 9137 26911
rect 8527 26880 9137 26908
rect 8527 26877 8539 26880
rect 8481 26871 8539 26877
rect 9125 26877 9137 26880
rect 9171 26877 9183 26911
rect 9125 26871 9183 26877
rect 7882 26843 7940 26849
rect 7882 26809 7894 26843
rect 7928 26809 7940 26843
rect 7882 26803 7940 26809
rect 8754 26772 8760 26784
rect 7760 26744 8760 26772
rect 8754 26732 8760 26744
rect 8812 26732 8818 26784
rect 9140 26772 9168 26871
rect 9398 26840 9404 26852
rect 9359 26812 9404 26840
rect 9398 26800 9404 26812
rect 9456 26800 9462 26852
rect 9493 26843 9551 26849
rect 9493 26809 9505 26843
rect 9539 26809 9551 26843
rect 9493 26803 9551 26809
rect 9508 26772 9536 26803
rect 9140 26744 9536 26772
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 2317 26571 2375 26577
rect 2317 26537 2329 26571
rect 2363 26568 2375 26571
rect 2406 26568 2412 26580
rect 2363 26540 2412 26568
rect 2363 26537 2375 26540
rect 2317 26531 2375 26537
rect 2406 26528 2412 26540
rect 2464 26568 2470 26580
rect 2464 26540 2544 26568
rect 2464 26528 2470 26540
rect 2516 26509 2544 26540
rect 3510 26528 3516 26580
rect 3568 26568 3574 26580
rect 4203 26571 4261 26577
rect 4203 26568 4215 26571
rect 3568 26540 4215 26568
rect 3568 26528 3574 26540
rect 4203 26537 4215 26540
rect 4249 26537 4261 26571
rect 4203 26531 4261 26537
rect 5350 26528 5356 26580
rect 5408 26568 5414 26580
rect 6273 26571 6331 26577
rect 6273 26568 6285 26571
rect 5408 26540 6285 26568
rect 5408 26528 5414 26540
rect 6273 26537 6285 26540
rect 6319 26568 6331 26571
rect 6638 26568 6644 26580
rect 6319 26540 6644 26568
rect 6319 26537 6331 26540
rect 6273 26531 6331 26537
rect 6638 26528 6644 26540
rect 6696 26528 6702 26580
rect 8481 26571 8539 26577
rect 8481 26537 8493 26571
rect 8527 26568 8539 26571
rect 8570 26568 8576 26580
rect 8527 26540 8576 26568
rect 8527 26537 8539 26540
rect 8481 26531 8539 26537
rect 8570 26528 8576 26540
rect 8628 26528 8634 26580
rect 9674 26528 9680 26580
rect 9732 26568 9738 26580
rect 9861 26571 9919 26577
rect 9861 26568 9873 26571
rect 9732 26540 9873 26568
rect 9732 26528 9738 26540
rect 9861 26537 9873 26540
rect 9907 26537 9919 26571
rect 9861 26531 9919 26537
rect 2501 26503 2559 26509
rect 2501 26469 2513 26503
rect 2547 26469 2559 26503
rect 2501 26463 2559 26469
rect 2593 26503 2651 26509
rect 2593 26469 2605 26503
rect 2639 26500 2651 26503
rect 3142 26500 3148 26512
rect 2639 26472 3148 26500
rect 2639 26469 2651 26472
rect 2593 26463 2651 26469
rect 3142 26460 3148 26472
rect 3200 26460 3206 26512
rect 4982 26460 4988 26512
rect 5040 26500 5046 26512
rect 5674 26503 5732 26509
rect 5674 26500 5686 26503
rect 5040 26472 5686 26500
rect 5040 26460 5046 26472
rect 5674 26469 5686 26472
rect 5720 26469 5732 26503
rect 5674 26463 5732 26469
rect 7923 26503 7981 26509
rect 7923 26469 7935 26503
rect 7969 26500 7981 26503
rect 8110 26500 8116 26512
rect 7969 26472 8116 26500
rect 7969 26469 7981 26472
rect 7923 26463 7981 26469
rect 8110 26460 8116 26472
rect 8168 26460 8174 26512
rect 4154 26441 4160 26444
rect 4132 26435 4160 26441
rect 4132 26401 4144 26435
rect 4132 26395 4160 26401
rect 4154 26392 4160 26395
rect 4212 26392 4218 26444
rect 5534 26392 5540 26444
rect 5592 26432 5598 26444
rect 6641 26435 6699 26441
rect 6641 26432 6653 26435
rect 5592 26404 6653 26432
rect 5592 26392 5598 26404
rect 6641 26401 6653 26404
rect 6687 26432 6699 26435
rect 6730 26432 6736 26444
rect 6687 26404 6736 26432
rect 6687 26401 6699 26404
rect 6641 26395 6699 26401
rect 6730 26392 6736 26404
rect 6788 26392 6794 26444
rect 3145 26367 3203 26373
rect 3145 26333 3157 26367
rect 3191 26364 3203 26367
rect 4430 26364 4436 26376
rect 3191 26336 4436 26364
rect 3191 26333 3203 26336
rect 3145 26327 3203 26333
rect 4430 26324 4436 26336
rect 4488 26324 4494 26376
rect 5353 26367 5411 26373
rect 5353 26333 5365 26367
rect 5399 26364 5411 26367
rect 5994 26364 6000 26376
rect 5399 26336 6000 26364
rect 5399 26333 5411 26336
rect 5353 26327 5411 26333
rect 5994 26324 6000 26336
rect 6052 26324 6058 26376
rect 7101 26367 7159 26373
rect 7101 26333 7113 26367
rect 7147 26364 7159 26367
rect 7561 26367 7619 26373
rect 7561 26364 7573 26367
rect 7147 26336 7573 26364
rect 7147 26333 7159 26336
rect 7101 26327 7159 26333
rect 7561 26333 7573 26336
rect 7607 26364 7619 26367
rect 9306 26364 9312 26376
rect 7607 26336 9312 26364
rect 7607 26333 7619 26336
rect 7561 26327 7619 26333
rect 9306 26324 9312 26336
rect 9364 26324 9370 26376
rect 3510 26228 3516 26240
rect 3471 26200 3516 26228
rect 3510 26188 3516 26200
rect 3568 26188 3574 26240
rect 4617 26231 4675 26237
rect 4617 26197 4629 26231
rect 4663 26228 4675 26231
rect 4706 26228 4712 26240
rect 4663 26200 4712 26228
rect 4663 26197 4675 26200
rect 4617 26191 4675 26197
rect 4706 26188 4712 26200
rect 4764 26188 4770 26240
rect 4982 26188 4988 26240
rect 5040 26228 5046 26240
rect 5077 26231 5135 26237
rect 5077 26228 5089 26231
rect 5040 26200 5089 26228
rect 5040 26188 5046 26200
rect 5077 26197 5089 26200
rect 5123 26197 5135 26231
rect 5077 26191 5135 26197
rect 7374 26188 7380 26240
rect 7432 26228 7438 26240
rect 7469 26231 7527 26237
rect 7469 26228 7481 26231
rect 7432 26200 7481 26228
rect 7432 26188 7438 26200
rect 7469 26197 7481 26200
rect 7515 26228 7527 26231
rect 8478 26228 8484 26240
rect 7515 26200 8484 26228
rect 7515 26197 7527 26200
rect 7469 26191 7527 26197
rect 8478 26188 8484 26200
rect 8536 26188 8542 26240
rect 9398 26228 9404 26240
rect 9311 26200 9404 26228
rect 9398 26188 9404 26200
rect 9456 26228 9462 26240
rect 10686 26228 10692 26240
rect 9456 26200 10692 26228
rect 9456 26188 9462 26200
rect 10686 26188 10692 26200
rect 10744 26188 10750 26240
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 4154 25984 4160 26036
rect 4212 26024 4218 26036
rect 5166 26024 5172 26036
rect 4212 25996 5172 26024
rect 4212 25984 4218 25996
rect 5166 25984 5172 25996
rect 5224 26024 5230 26036
rect 5626 26024 5632 26036
rect 5224 25996 5632 26024
rect 5224 25984 5230 25996
rect 5626 25984 5632 25996
rect 5684 25984 5690 26036
rect 6638 26024 6644 26036
rect 6599 25996 6644 26024
rect 6638 25984 6644 25996
rect 6696 25984 6702 26036
rect 1673 25959 1731 25965
rect 1673 25925 1685 25959
rect 1719 25956 1731 25959
rect 3142 25956 3148 25968
rect 1719 25928 3148 25956
rect 1719 25925 1731 25928
rect 1673 25919 1731 25925
rect 3142 25916 3148 25928
rect 3200 25916 3206 25968
rect 1903 25891 1961 25897
rect 1903 25857 1915 25891
rect 1949 25888 1961 25891
rect 4890 25888 4896 25900
rect 1949 25860 4476 25888
rect 4851 25860 4896 25888
rect 1949 25857 1961 25860
rect 1903 25851 1961 25857
rect 1302 25780 1308 25832
rect 1360 25820 1366 25832
rect 1800 25823 1858 25829
rect 1800 25820 1812 25823
rect 1360 25792 1812 25820
rect 1360 25780 1366 25792
rect 1800 25789 1812 25792
rect 1846 25820 1858 25823
rect 2225 25823 2283 25829
rect 2225 25820 2237 25823
rect 1846 25792 2237 25820
rect 1846 25789 1858 25792
rect 1800 25783 1858 25789
rect 2225 25789 2237 25792
rect 2271 25820 2283 25823
rect 2314 25820 2320 25832
rect 2271 25792 2320 25820
rect 2271 25789 2283 25792
rect 2225 25783 2283 25789
rect 2314 25780 2320 25792
rect 2372 25780 2378 25832
rect 2777 25823 2835 25829
rect 2777 25789 2789 25823
rect 2823 25820 2835 25823
rect 3418 25820 3424 25832
rect 2823 25792 3424 25820
rect 2823 25789 2835 25792
rect 2777 25783 2835 25789
rect 3418 25780 3424 25792
rect 3476 25780 3482 25832
rect 3510 25780 3516 25832
rect 3568 25820 3574 25832
rect 3697 25823 3755 25829
rect 3697 25820 3709 25823
rect 3568 25792 3709 25820
rect 3568 25780 3574 25792
rect 3697 25789 3709 25792
rect 3743 25820 3755 25823
rect 4246 25820 4252 25832
rect 3743 25792 4252 25820
rect 3743 25789 3755 25792
rect 3697 25783 3755 25789
rect 4246 25780 4252 25792
rect 4304 25780 4310 25832
rect 3099 25755 3157 25761
rect 3099 25721 3111 25755
rect 3145 25721 3157 25755
rect 4448 25752 4476 25860
rect 4890 25848 4896 25860
rect 4948 25848 4954 25900
rect 6730 25848 6736 25900
rect 6788 25888 6794 25900
rect 6917 25891 6975 25897
rect 6917 25888 6929 25891
rect 6788 25860 6929 25888
rect 6788 25848 6794 25860
rect 6917 25857 6929 25860
rect 6963 25857 6975 25891
rect 6917 25851 6975 25857
rect 7190 25848 7196 25900
rect 7248 25888 7254 25900
rect 7285 25891 7343 25897
rect 7285 25888 7297 25891
rect 7248 25860 7297 25888
rect 7248 25848 7254 25860
rect 7285 25857 7297 25860
rect 7331 25857 7343 25891
rect 7285 25851 7343 25857
rect 8573 25891 8631 25897
rect 8573 25857 8585 25891
rect 8619 25888 8631 25891
rect 8846 25888 8852 25900
rect 8619 25860 8852 25888
rect 8619 25857 8631 25860
rect 8573 25851 8631 25857
rect 8846 25848 8852 25860
rect 8904 25848 8910 25900
rect 4614 25752 4620 25764
rect 4448 25724 4620 25752
rect 3099 25715 3157 25721
rect 2590 25684 2596 25696
rect 2551 25656 2596 25684
rect 2590 25644 2596 25656
rect 2648 25684 2654 25696
rect 3114 25684 3142 25715
rect 4614 25712 4620 25724
rect 4672 25712 4678 25764
rect 4706 25712 4712 25764
rect 4764 25752 4770 25764
rect 7009 25755 7067 25761
rect 4764 25724 4809 25752
rect 4764 25712 4770 25724
rect 7009 25721 7021 25755
rect 7055 25721 7067 25755
rect 7009 25715 7067 25721
rect 8389 25755 8447 25761
rect 8389 25721 8401 25755
rect 8435 25752 8447 25755
rect 8662 25752 8668 25764
rect 8435 25724 8668 25752
rect 8435 25721 8447 25724
rect 8389 25715 8447 25721
rect 4982 25684 4988 25696
rect 2648 25656 4988 25684
rect 2648 25644 2654 25656
rect 4982 25644 4988 25656
rect 5040 25684 5046 25696
rect 5537 25687 5595 25693
rect 5537 25684 5549 25687
rect 5040 25656 5549 25684
rect 5040 25644 5046 25656
rect 5537 25653 5549 25656
rect 5583 25653 5595 25687
rect 5994 25684 6000 25696
rect 5955 25656 6000 25684
rect 5537 25647 5595 25653
rect 5994 25644 6000 25656
rect 6052 25644 6058 25696
rect 6638 25644 6644 25696
rect 6696 25684 6702 25696
rect 7024 25684 7052 25715
rect 8662 25712 8668 25724
rect 8720 25712 8726 25764
rect 9217 25755 9275 25761
rect 9217 25721 9229 25755
rect 9263 25752 9275 25755
rect 9858 25752 9864 25764
rect 9263 25724 9864 25752
rect 9263 25721 9275 25724
rect 9217 25715 9275 25721
rect 9858 25712 9864 25724
rect 9916 25712 9922 25764
rect 6696 25656 7052 25684
rect 7929 25687 7987 25693
rect 6696 25644 6702 25656
rect 7929 25653 7941 25687
rect 7975 25684 7987 25687
rect 8110 25684 8116 25696
rect 7975 25656 8116 25684
rect 7975 25653 7987 25656
rect 7929 25647 7987 25653
rect 8110 25644 8116 25656
rect 8168 25644 8174 25696
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 2590 25480 2596 25492
rect 2551 25452 2596 25480
rect 2590 25440 2596 25452
rect 2648 25440 2654 25492
rect 4614 25440 4620 25492
rect 4672 25480 4678 25492
rect 5077 25483 5135 25489
rect 5077 25480 5089 25483
rect 4672 25452 5089 25480
rect 4672 25440 4678 25452
rect 5077 25449 5089 25452
rect 5123 25449 5135 25483
rect 5077 25443 5135 25449
rect 5994 25440 6000 25492
rect 6052 25480 6058 25492
rect 7285 25483 7343 25489
rect 7285 25480 7297 25483
rect 6052 25452 7297 25480
rect 6052 25440 6058 25452
rect 7285 25449 7297 25452
rect 7331 25449 7343 25483
rect 7285 25443 7343 25449
rect 10321 25483 10379 25489
rect 10321 25449 10333 25483
rect 10367 25480 10379 25483
rect 13814 25480 13820 25492
rect 10367 25452 13820 25480
rect 10367 25449 10379 25452
rect 10321 25443 10379 25449
rect 13814 25440 13820 25452
rect 13872 25440 13878 25492
rect 4246 25372 4252 25424
rect 4304 25412 4310 25424
rect 4982 25412 4988 25424
rect 4304 25384 4988 25412
rect 4304 25372 4310 25384
rect 4982 25372 4988 25384
rect 5040 25372 5046 25424
rect 5442 25372 5448 25424
rect 5500 25412 5506 25424
rect 5813 25415 5871 25421
rect 5813 25412 5825 25415
rect 5500 25384 5825 25412
rect 5500 25372 5506 25384
rect 5813 25381 5825 25384
rect 5859 25381 5871 25415
rect 5813 25375 5871 25381
rect 7469 25347 7527 25353
rect 7469 25313 7481 25347
rect 7515 25313 7527 25347
rect 7650 25344 7656 25356
rect 7611 25316 7656 25344
rect 7469 25307 7527 25313
rect 2222 25276 2228 25288
rect 2183 25248 2228 25276
rect 2222 25236 2228 25248
rect 2280 25236 2286 25288
rect 3881 25279 3939 25285
rect 3881 25245 3893 25279
rect 3927 25276 3939 25279
rect 4154 25276 4160 25288
rect 3927 25248 4160 25276
rect 3927 25245 3939 25248
rect 3881 25239 3939 25245
rect 4154 25236 4160 25248
rect 4212 25236 4218 25288
rect 4430 25276 4436 25288
rect 4391 25248 4436 25276
rect 4430 25236 4436 25248
rect 4488 25276 4494 25288
rect 4488 25248 4752 25276
rect 4488 25236 4494 25248
rect 3142 25208 3148 25220
rect 3055 25180 3148 25208
rect 3142 25168 3148 25180
rect 3200 25208 3206 25220
rect 4614 25208 4620 25220
rect 3200 25180 4620 25208
rect 3200 25168 3206 25180
rect 4614 25168 4620 25180
rect 4672 25168 4678 25220
rect 4724 25208 4752 25248
rect 5534 25236 5540 25288
rect 5592 25276 5598 25288
rect 5721 25279 5779 25285
rect 5721 25276 5733 25279
rect 5592 25248 5733 25276
rect 5592 25236 5598 25248
rect 5721 25245 5733 25248
rect 5767 25245 5779 25279
rect 5721 25239 5779 25245
rect 5997 25279 6055 25285
rect 5997 25245 6009 25279
rect 6043 25245 6055 25279
rect 7484 25276 7512 25307
rect 7650 25304 7656 25316
rect 7708 25304 7714 25356
rect 8386 25304 8392 25356
rect 8444 25344 8450 25356
rect 10137 25347 10195 25353
rect 10137 25344 10149 25347
rect 8444 25316 10149 25344
rect 8444 25304 8450 25316
rect 10137 25313 10149 25316
rect 10183 25344 10195 25347
rect 10962 25344 10968 25356
rect 10183 25316 10968 25344
rect 10183 25313 10195 25316
rect 10137 25307 10195 25313
rect 10962 25304 10968 25316
rect 11020 25304 11026 25356
rect 7834 25276 7840 25288
rect 7484 25248 7840 25276
rect 5997 25239 6055 25245
rect 6012 25208 6040 25239
rect 7834 25236 7840 25248
rect 7892 25236 7898 25288
rect 4724 25180 6040 25208
rect 3418 25140 3424 25152
rect 3379 25112 3424 25140
rect 3418 25100 3424 25112
rect 3476 25100 3482 25152
rect 3510 25100 3516 25152
rect 3568 25140 3574 25152
rect 6825 25143 6883 25149
rect 6825 25140 6837 25143
rect 3568 25112 6837 25140
rect 3568 25100 3574 25112
rect 6825 25109 6837 25112
rect 6871 25140 6883 25143
rect 7282 25140 7288 25152
rect 6871 25112 7288 25140
rect 6871 25109 6883 25112
rect 6825 25103 6883 25109
rect 7282 25100 7288 25112
rect 7340 25140 7346 25152
rect 7650 25140 7656 25152
rect 7340 25112 7656 25140
rect 7340 25100 7346 25112
rect 7650 25100 7656 25112
rect 7708 25100 7714 25152
rect 8294 25100 8300 25152
rect 8352 25140 8358 25152
rect 8389 25143 8447 25149
rect 8389 25140 8401 25143
rect 8352 25112 8401 25140
rect 8352 25100 8358 25112
rect 8389 25109 8401 25112
rect 8435 25109 8447 25143
rect 8846 25140 8852 25152
rect 8807 25112 8852 25140
rect 8389 25103 8447 25109
rect 8846 25100 8852 25112
rect 8904 25100 8910 25152
rect 10042 25140 10048 25152
rect 10003 25112 10048 25140
rect 10042 25100 10048 25112
rect 10100 25100 10106 25152
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 3329 24939 3387 24945
rect 3329 24905 3341 24939
rect 3375 24936 3387 24939
rect 3510 24936 3516 24948
rect 3375 24908 3516 24936
rect 3375 24905 3387 24908
rect 3329 24899 3387 24905
rect 2958 24800 2964 24812
rect 2919 24772 2964 24800
rect 2958 24760 2964 24772
rect 3016 24760 3022 24812
rect 1765 24735 1823 24741
rect 1765 24701 1777 24735
rect 1811 24732 1823 24735
rect 1946 24732 1952 24744
rect 1811 24704 1952 24732
rect 1811 24701 1823 24704
rect 1765 24695 1823 24701
rect 1946 24692 1952 24704
rect 2004 24732 2010 24744
rect 2225 24735 2283 24741
rect 2225 24732 2237 24735
rect 2004 24704 2237 24732
rect 2004 24692 2010 24704
rect 2225 24701 2237 24704
rect 2271 24701 2283 24735
rect 2225 24695 2283 24701
rect 2777 24735 2835 24741
rect 2777 24701 2789 24735
rect 2823 24732 2835 24735
rect 3344 24732 3372 24899
rect 3510 24896 3516 24908
rect 3568 24896 3574 24948
rect 4982 24936 4988 24948
rect 4943 24908 4988 24936
rect 4982 24896 4988 24908
rect 5040 24896 5046 24948
rect 5442 24936 5448 24948
rect 5403 24908 5448 24936
rect 5442 24896 5448 24908
rect 5500 24896 5506 24948
rect 10962 24936 10968 24948
rect 10923 24908 10968 24936
rect 10962 24896 10968 24908
rect 11020 24896 11026 24948
rect 4246 24828 4252 24880
rect 4304 24868 4310 24880
rect 4709 24871 4767 24877
rect 4709 24868 4721 24871
rect 4304 24840 4721 24868
rect 4304 24828 4310 24840
rect 4709 24837 4721 24840
rect 4755 24868 4767 24871
rect 5460 24868 5488 24896
rect 4755 24840 5488 24868
rect 4755 24837 4767 24840
rect 4709 24831 4767 24837
rect 4338 24760 4344 24812
rect 4396 24800 4402 24812
rect 4982 24800 4988 24812
rect 4396 24772 4988 24800
rect 4396 24760 4402 24772
rect 4982 24760 4988 24772
rect 5040 24760 5046 24812
rect 5258 24760 5264 24812
rect 5316 24800 5322 24812
rect 5997 24803 6055 24809
rect 5997 24800 6009 24803
rect 5316 24772 6009 24800
rect 5316 24760 5322 24772
rect 2823 24704 3372 24732
rect 3789 24735 3847 24741
rect 2823 24701 2835 24704
rect 2777 24695 2835 24701
rect 3789 24701 3801 24735
rect 3835 24732 3847 24735
rect 3878 24732 3884 24744
rect 3835 24704 3884 24732
rect 3835 24701 3847 24704
rect 3789 24695 3847 24701
rect 3878 24692 3884 24704
rect 3936 24692 3942 24744
rect 5619 24741 5647 24772
rect 5997 24769 6009 24772
rect 6043 24800 6055 24803
rect 6730 24800 6736 24812
rect 6043 24772 6736 24800
rect 6043 24769 6055 24772
rect 5997 24763 6055 24769
rect 6730 24760 6736 24772
rect 6788 24760 6794 24812
rect 10042 24800 10048 24812
rect 10003 24772 10048 24800
rect 10042 24760 10048 24772
rect 10100 24760 10106 24812
rect 5604 24735 5662 24741
rect 5604 24701 5616 24735
rect 5650 24701 5662 24735
rect 5604 24695 5662 24701
rect 6825 24735 6883 24741
rect 6825 24701 6837 24735
rect 6871 24701 6883 24735
rect 7282 24732 7288 24744
rect 7243 24704 7288 24732
rect 6825 24695 6883 24701
rect 4522 24624 4528 24676
rect 4580 24664 4586 24676
rect 6549 24667 6607 24673
rect 6549 24664 6561 24667
rect 4580 24636 6561 24664
rect 4580 24624 4586 24636
rect 6549 24633 6561 24636
rect 6595 24664 6607 24667
rect 6840 24664 6868 24695
rect 7282 24692 7288 24704
rect 7340 24692 7346 24744
rect 8294 24692 8300 24744
rect 8352 24732 8358 24744
rect 8389 24735 8447 24741
rect 8389 24732 8401 24735
rect 8352 24704 8401 24732
rect 8352 24692 8358 24704
rect 8389 24701 8401 24704
rect 8435 24701 8447 24735
rect 8389 24695 8447 24701
rect 8849 24735 8907 24741
rect 8849 24701 8861 24735
rect 8895 24701 8907 24735
rect 8849 24695 8907 24701
rect 8864 24664 8892 24695
rect 10137 24667 10195 24673
rect 10137 24664 10149 24667
rect 6595 24636 6868 24664
rect 8220 24636 8892 24664
rect 9784 24636 10149 24664
rect 6595 24633 6607 24636
rect 6549 24627 6607 24633
rect 2133 24599 2191 24605
rect 2133 24565 2145 24599
rect 2179 24596 2191 24599
rect 2590 24596 2596 24608
rect 2179 24568 2596 24596
rect 2179 24565 2191 24568
rect 2133 24559 2191 24565
rect 2590 24556 2596 24568
rect 2648 24596 2654 24608
rect 3697 24599 3755 24605
rect 3697 24596 3709 24599
rect 2648 24568 3709 24596
rect 2648 24556 2654 24568
rect 3697 24565 3709 24568
rect 3743 24596 3755 24599
rect 3970 24596 3976 24608
rect 3743 24568 3976 24596
rect 3743 24565 3755 24568
rect 3697 24559 3755 24565
rect 3970 24556 3976 24568
rect 4028 24556 4034 24608
rect 4154 24596 4160 24608
rect 4115 24568 4160 24596
rect 4154 24556 4160 24568
rect 4212 24556 4218 24608
rect 4338 24556 4344 24608
rect 4396 24596 4402 24608
rect 4798 24596 4804 24608
rect 4396 24568 4804 24596
rect 4396 24556 4402 24568
rect 4798 24556 4804 24568
rect 4856 24596 4862 24608
rect 5675 24599 5733 24605
rect 5675 24596 5687 24599
rect 4856 24568 5687 24596
rect 4856 24556 4862 24568
rect 5675 24565 5687 24568
rect 5721 24565 5733 24599
rect 6914 24596 6920 24608
rect 6875 24568 6920 24596
rect 5675 24559 5733 24565
rect 6914 24556 6920 24568
rect 6972 24556 6978 24608
rect 7834 24596 7840 24608
rect 7795 24568 7840 24596
rect 7834 24556 7840 24568
rect 7892 24556 7898 24608
rect 7926 24556 7932 24608
rect 7984 24596 7990 24608
rect 8220 24605 8248 24636
rect 8205 24599 8263 24605
rect 8205 24596 8217 24599
rect 7984 24568 8217 24596
rect 7984 24556 7990 24568
rect 8205 24565 8217 24568
rect 8251 24565 8263 24599
rect 8478 24596 8484 24608
rect 8439 24568 8484 24596
rect 8205 24559 8263 24565
rect 8478 24556 8484 24568
rect 8536 24556 8542 24608
rect 9582 24556 9588 24608
rect 9640 24596 9646 24608
rect 9784 24605 9812 24636
rect 10137 24633 10149 24636
rect 10183 24633 10195 24667
rect 10686 24664 10692 24676
rect 10647 24636 10692 24664
rect 10137 24627 10195 24633
rect 10686 24624 10692 24636
rect 10744 24624 10750 24676
rect 9769 24599 9827 24605
rect 9769 24596 9781 24599
rect 9640 24568 9781 24596
rect 9640 24556 9646 24568
rect 9769 24565 9781 24568
rect 9815 24565 9827 24599
rect 9769 24559 9827 24565
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 2133 24395 2191 24401
rect 2133 24361 2145 24395
rect 2179 24392 2191 24395
rect 2222 24392 2228 24404
rect 2179 24364 2228 24392
rect 2179 24361 2191 24364
rect 2133 24355 2191 24361
rect 2222 24352 2228 24364
rect 2280 24392 2286 24404
rect 2317 24395 2375 24401
rect 2317 24392 2329 24395
rect 2280 24364 2329 24392
rect 2280 24352 2286 24364
rect 2317 24361 2329 24364
rect 2363 24361 2375 24395
rect 2317 24355 2375 24361
rect 4706 24352 4712 24404
rect 4764 24352 4770 24404
rect 7282 24392 7288 24404
rect 7243 24364 7288 24392
rect 7282 24352 7288 24364
rect 7340 24352 7346 24404
rect 7558 24392 7564 24404
rect 7519 24364 7564 24392
rect 7558 24352 7564 24364
rect 7616 24352 7622 24404
rect 11425 24395 11483 24401
rect 11425 24361 11437 24395
rect 11471 24392 11483 24395
rect 11514 24392 11520 24404
rect 11471 24364 11520 24392
rect 11471 24361 11483 24364
rect 11425 24355 11483 24361
rect 11514 24352 11520 24364
rect 11572 24352 11578 24404
rect 4246 24324 4252 24336
rect 4207 24296 4252 24324
rect 4246 24284 4252 24296
rect 4304 24284 4310 24336
rect 4724 24324 4752 24352
rect 4801 24327 4859 24333
rect 4801 24324 4813 24327
rect 4724 24296 4813 24324
rect 4801 24293 4813 24296
rect 4847 24324 4859 24327
rect 4890 24324 4896 24336
rect 4847 24296 4896 24324
rect 4847 24293 4859 24296
rect 4801 24287 4859 24293
rect 4890 24284 4896 24296
rect 4948 24284 4954 24336
rect 6086 24324 6092 24336
rect 6047 24296 6092 24324
rect 6086 24284 6092 24296
rect 6144 24284 6150 24336
rect 9582 24284 9588 24336
rect 9640 24324 9646 24336
rect 9861 24327 9919 24333
rect 9861 24324 9873 24327
rect 9640 24296 9873 24324
rect 9640 24284 9646 24296
rect 9861 24293 9873 24296
rect 9907 24293 9919 24327
rect 9861 24287 9919 24293
rect 2501 24259 2559 24265
rect 2501 24225 2513 24259
rect 2547 24225 2559 24259
rect 2682 24256 2688 24268
rect 2643 24228 2688 24256
rect 2501 24219 2559 24225
rect 2516 24188 2544 24219
rect 2682 24216 2688 24228
rect 2740 24216 2746 24268
rect 7466 24256 7472 24268
rect 7427 24228 7472 24256
rect 7466 24216 7472 24228
rect 7524 24216 7530 24268
rect 7926 24256 7932 24268
rect 7887 24228 7932 24256
rect 7926 24216 7932 24228
rect 7984 24216 7990 24268
rect 11238 24256 11244 24268
rect 11199 24228 11244 24256
rect 11238 24216 11244 24228
rect 11296 24216 11302 24268
rect 3142 24188 3148 24200
rect 2516 24160 3148 24188
rect 3142 24148 3148 24160
rect 3200 24148 3206 24200
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 4338 24188 4344 24200
rect 4203 24160 4344 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4338 24148 4344 24160
rect 4396 24148 4402 24200
rect 5718 24148 5724 24200
rect 5776 24188 5782 24200
rect 5997 24191 6055 24197
rect 5997 24188 6009 24191
rect 5776 24160 6009 24188
rect 5776 24148 5782 24160
rect 5997 24157 6009 24160
rect 6043 24157 6055 24191
rect 5997 24151 6055 24157
rect 6641 24191 6699 24197
rect 6641 24157 6653 24191
rect 6687 24188 6699 24191
rect 7374 24188 7380 24200
rect 6687 24160 7380 24188
rect 6687 24157 6699 24160
rect 6641 24151 6699 24157
rect 7374 24148 7380 24160
rect 7432 24148 7438 24200
rect 9766 24188 9772 24200
rect 9727 24160 9772 24188
rect 9766 24148 9772 24160
rect 9824 24148 9830 24200
rect 9858 24148 9864 24200
rect 9916 24188 9922 24200
rect 10045 24191 10103 24197
rect 10045 24188 10057 24191
rect 9916 24160 10057 24188
rect 9916 24148 9922 24160
rect 10045 24157 10057 24160
rect 10091 24157 10103 24191
rect 10045 24151 10103 24157
rect 3160 24120 3188 24148
rect 4522 24120 4528 24132
rect 3160 24092 4528 24120
rect 4522 24080 4528 24092
rect 4580 24080 4586 24132
rect 5258 24080 5264 24132
rect 5316 24120 5322 24132
rect 7190 24120 7196 24132
rect 5316 24092 7196 24120
rect 5316 24080 5322 24092
rect 7190 24080 7196 24092
rect 7248 24080 7254 24132
rect 3881 24055 3939 24061
rect 3881 24021 3893 24055
rect 3927 24052 3939 24055
rect 3970 24052 3976 24064
rect 3927 24024 3976 24052
rect 3927 24021 3939 24024
rect 3881 24015 3939 24021
rect 3970 24012 3976 24024
rect 4028 24052 4034 24064
rect 4154 24052 4160 24064
rect 4028 24024 4160 24052
rect 4028 24012 4034 24024
rect 4154 24012 4160 24024
rect 4212 24012 4218 24064
rect 4614 24012 4620 24064
rect 4672 24052 4678 24064
rect 5534 24052 5540 24064
rect 4672 24024 5540 24052
rect 4672 24012 4678 24024
rect 5534 24012 5540 24024
rect 5592 24052 5598 24064
rect 5629 24055 5687 24061
rect 5629 24052 5641 24055
rect 5592 24024 5641 24052
rect 5592 24012 5598 24024
rect 5629 24021 5641 24024
rect 5675 24021 5687 24055
rect 8478 24052 8484 24064
rect 8439 24024 8484 24052
rect 5629 24015 5687 24021
rect 8478 24012 8484 24024
rect 8536 24012 8542 24064
rect 11514 24012 11520 24064
rect 11572 24052 11578 24064
rect 12710 24052 12716 24064
rect 11572 24024 12716 24052
rect 11572 24012 11578 24024
rect 12710 24012 12716 24024
rect 12768 24012 12774 24064
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 1946 23848 1952 23860
rect 1907 23820 1952 23848
rect 1946 23808 1952 23820
rect 2004 23808 2010 23860
rect 4246 23808 4252 23860
rect 4304 23848 4310 23860
rect 4617 23851 4675 23857
rect 4617 23848 4629 23851
rect 4304 23820 4629 23848
rect 4304 23808 4310 23820
rect 4617 23817 4629 23820
rect 4663 23817 4675 23851
rect 4617 23811 4675 23817
rect 6086 23808 6092 23860
rect 6144 23848 6150 23860
rect 6549 23851 6607 23857
rect 6549 23848 6561 23851
rect 6144 23820 6561 23848
rect 6144 23808 6150 23820
rect 6549 23817 6561 23820
rect 6595 23817 6607 23851
rect 6549 23811 6607 23817
rect 7285 23851 7343 23857
rect 7285 23817 7297 23851
rect 7331 23848 7343 23851
rect 7926 23848 7932 23860
rect 7331 23820 7932 23848
rect 7331 23817 7343 23820
rect 7285 23811 7343 23817
rect 7926 23808 7932 23820
rect 7984 23808 7990 23860
rect 8662 23848 8668 23860
rect 8623 23820 8668 23848
rect 8662 23808 8668 23820
rect 8720 23808 8726 23860
rect 9766 23808 9772 23860
rect 9824 23848 9830 23860
rect 10873 23851 10931 23857
rect 10873 23848 10885 23851
rect 9824 23820 10885 23848
rect 9824 23808 9830 23820
rect 10873 23817 10885 23820
rect 10919 23817 10931 23851
rect 10873 23811 10931 23817
rect 7834 23780 7840 23792
rect 3620 23752 7840 23780
rect 2777 23715 2835 23721
rect 2777 23681 2789 23715
rect 2823 23712 2835 23715
rect 3418 23712 3424 23724
rect 2823 23684 3424 23712
rect 2823 23681 2835 23684
rect 2777 23675 2835 23681
rect 3418 23672 3424 23684
rect 3476 23672 3482 23724
rect 1946 23604 1952 23656
rect 2004 23644 2010 23656
rect 2041 23647 2099 23653
rect 2041 23644 2053 23647
rect 2004 23616 2053 23644
rect 2004 23604 2010 23616
rect 2041 23613 2053 23616
rect 2087 23644 2099 23647
rect 2130 23644 2136 23656
rect 2087 23616 2136 23644
rect 2087 23613 2099 23616
rect 2041 23607 2099 23613
rect 2130 23604 2136 23616
rect 2188 23604 2194 23656
rect 2593 23647 2651 23653
rect 2593 23613 2605 23647
rect 2639 23644 2651 23647
rect 2682 23644 2688 23656
rect 2639 23616 2688 23644
rect 2639 23613 2651 23616
rect 2593 23607 2651 23613
rect 2682 23604 2688 23616
rect 2740 23604 2746 23656
rect 3620 23653 3648 23752
rect 7834 23740 7840 23752
rect 7892 23740 7898 23792
rect 7944 23780 7972 23808
rect 9309 23783 9367 23789
rect 9309 23780 9321 23783
rect 7944 23752 9321 23780
rect 9309 23749 9321 23752
rect 9355 23749 9367 23783
rect 9309 23743 9367 23749
rect 4154 23712 4160 23724
rect 4115 23684 4160 23712
rect 4154 23672 4160 23684
rect 4212 23672 4218 23724
rect 5077 23715 5135 23721
rect 5077 23681 5089 23715
rect 5123 23712 5135 23715
rect 5626 23712 5632 23724
rect 5123 23684 5632 23712
rect 5123 23681 5135 23684
rect 5077 23675 5135 23681
rect 5626 23672 5632 23684
rect 5684 23672 5690 23724
rect 7745 23715 7803 23721
rect 7745 23681 7757 23715
rect 7791 23712 7803 23715
rect 8478 23712 8484 23724
rect 7791 23684 8484 23712
rect 7791 23681 7803 23684
rect 7745 23675 7803 23681
rect 8478 23672 8484 23684
rect 8536 23672 8542 23724
rect 9324 23712 9352 23743
rect 9324 23684 9996 23712
rect 3605 23647 3663 23653
rect 3605 23613 3617 23647
rect 3651 23613 3663 23647
rect 3605 23607 3663 23613
rect 1578 23536 1584 23588
rect 1636 23576 1642 23588
rect 3421 23579 3479 23585
rect 3421 23576 3433 23579
rect 1636 23548 3433 23576
rect 1636 23536 1642 23548
rect 3421 23545 3433 23548
rect 3467 23576 3479 23579
rect 3620 23576 3648 23607
rect 3970 23604 3976 23656
rect 4028 23644 4034 23656
rect 9968 23653 9996 23684
rect 4065 23647 4123 23653
rect 4065 23644 4077 23647
rect 4028 23616 4077 23644
rect 4028 23604 4034 23616
rect 4065 23613 4077 23616
rect 4111 23613 4123 23647
rect 9493 23647 9551 23653
rect 9493 23644 9505 23647
rect 4065 23607 4123 23613
rect 8956 23616 9505 23644
rect 5258 23576 5264 23588
rect 3467 23548 3648 23576
rect 5219 23548 5264 23576
rect 3467 23545 3479 23548
rect 3421 23539 3479 23545
rect 5258 23536 5264 23548
rect 5316 23536 5322 23588
rect 5362 23579 5420 23585
rect 5362 23545 5374 23579
rect 5408 23576 5420 23579
rect 5626 23576 5632 23588
rect 5408 23548 5632 23576
rect 5408 23545 5420 23548
rect 5362 23539 5420 23545
rect 5626 23536 5632 23548
rect 5684 23536 5690 23588
rect 5905 23579 5963 23585
rect 5905 23545 5917 23579
rect 5951 23576 5963 23579
rect 5994 23576 6000 23588
rect 5951 23548 6000 23576
rect 5951 23545 5963 23548
rect 5905 23539 5963 23545
rect 5994 23536 6000 23548
rect 6052 23576 6058 23588
rect 7374 23576 7380 23588
rect 6052 23548 7380 23576
rect 6052 23536 6058 23548
rect 7374 23536 7380 23548
rect 7432 23536 7438 23588
rect 7653 23579 7711 23585
rect 7653 23545 7665 23579
rect 7699 23576 7711 23579
rect 7926 23576 7932 23588
rect 7699 23548 7932 23576
rect 7699 23545 7711 23548
rect 7653 23539 7711 23545
rect 7926 23536 7932 23548
rect 7984 23576 7990 23588
rect 8110 23585 8116 23588
rect 8066 23579 8116 23585
rect 8066 23576 8078 23579
rect 7984 23548 8078 23576
rect 7984 23536 7990 23548
rect 8066 23545 8078 23548
rect 8112 23545 8116 23579
rect 8066 23539 8116 23545
rect 8110 23536 8116 23539
rect 8168 23536 8174 23588
rect 3142 23508 3148 23520
rect 3103 23480 3148 23508
rect 3142 23468 3148 23480
rect 3200 23468 3206 23520
rect 5718 23468 5724 23520
rect 5776 23508 5782 23520
rect 6181 23511 6239 23517
rect 6181 23508 6193 23511
rect 5776 23480 6193 23508
rect 5776 23468 5782 23480
rect 6181 23477 6193 23480
rect 6227 23477 6239 23511
rect 6181 23471 6239 23477
rect 7742 23468 7748 23520
rect 7800 23508 7806 23520
rect 8956 23517 8984 23616
rect 9493 23613 9505 23616
rect 9539 23613 9551 23647
rect 9493 23607 9551 23613
rect 9953 23647 10011 23653
rect 9953 23613 9965 23647
rect 9999 23644 10011 23647
rect 10042 23644 10048 23656
rect 9999 23616 10048 23644
rect 9999 23613 10011 23616
rect 9953 23607 10011 23613
rect 10042 23604 10048 23616
rect 10100 23604 10106 23656
rect 11124 23647 11182 23653
rect 11124 23613 11136 23647
rect 11170 23644 11182 23647
rect 11238 23644 11244 23656
rect 11170 23616 11244 23644
rect 11170 23613 11182 23616
rect 11124 23607 11182 23613
rect 11238 23604 11244 23616
rect 11296 23644 11302 23656
rect 11296 23616 11652 23644
rect 11296 23604 11302 23616
rect 8941 23511 8999 23517
rect 8941 23508 8953 23511
rect 7800 23480 8953 23508
rect 7800 23468 7806 23480
rect 8941 23477 8953 23480
rect 8987 23477 8999 23511
rect 8941 23471 8999 23477
rect 9398 23468 9404 23520
rect 9456 23508 9462 23520
rect 9585 23511 9643 23517
rect 9585 23508 9597 23511
rect 9456 23480 9597 23508
rect 9456 23468 9462 23480
rect 9585 23477 9597 23480
rect 9631 23477 9643 23511
rect 9585 23471 9643 23477
rect 9674 23468 9680 23520
rect 9732 23508 9738 23520
rect 10505 23511 10563 23517
rect 10505 23508 10517 23511
rect 9732 23480 10517 23508
rect 9732 23468 9738 23480
rect 10505 23477 10517 23480
rect 10551 23477 10563 23511
rect 10505 23471 10563 23477
rect 10962 23468 10968 23520
rect 11020 23508 11026 23520
rect 11624 23517 11652 23616
rect 11195 23511 11253 23517
rect 11195 23508 11207 23511
rect 11020 23480 11207 23508
rect 11020 23468 11026 23480
rect 11195 23477 11207 23480
rect 11241 23477 11253 23511
rect 11195 23471 11253 23477
rect 11609 23511 11667 23517
rect 11609 23477 11621 23511
rect 11655 23508 11667 23511
rect 11977 23511 12035 23517
rect 11977 23508 11989 23511
rect 11655 23480 11989 23508
rect 11655 23477 11667 23480
rect 11609 23471 11667 23477
rect 11977 23477 11989 23480
rect 12023 23508 12035 23511
rect 12158 23508 12164 23520
rect 12023 23480 12164 23508
rect 12023 23477 12035 23480
rect 11977 23471 12035 23477
rect 12158 23468 12164 23480
rect 12216 23468 12222 23520
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 1118 23264 1124 23316
rect 1176 23304 1182 23316
rect 1535 23307 1593 23313
rect 1535 23304 1547 23307
rect 1176 23276 1547 23304
rect 1176 23264 1182 23276
rect 1535 23273 1547 23276
rect 1581 23273 1593 23307
rect 1535 23267 1593 23273
rect 4387 23307 4445 23313
rect 4387 23273 4399 23307
rect 4433 23304 4445 23307
rect 4614 23304 4620 23316
rect 4433 23276 4620 23304
rect 4433 23273 4445 23276
rect 4387 23267 4445 23273
rect 4614 23264 4620 23276
rect 4672 23264 4678 23316
rect 4798 23304 4804 23316
rect 4759 23276 4804 23304
rect 4798 23264 4804 23276
rect 4856 23264 4862 23316
rect 5258 23304 5264 23316
rect 5219 23276 5264 23304
rect 5258 23264 5264 23276
rect 5316 23264 5322 23316
rect 6086 23264 6092 23316
rect 6144 23304 6150 23316
rect 6365 23307 6423 23313
rect 6365 23304 6377 23307
rect 6144 23276 6377 23304
rect 6144 23264 6150 23276
rect 6365 23273 6377 23276
rect 6411 23273 6423 23307
rect 6365 23267 6423 23273
rect 6917 23307 6975 23313
rect 6917 23273 6929 23307
rect 6963 23304 6975 23307
rect 7006 23304 7012 23316
rect 6963 23276 7012 23304
rect 6963 23273 6975 23276
rect 6917 23267 6975 23273
rect 7006 23264 7012 23276
rect 7064 23264 7070 23316
rect 7466 23304 7472 23316
rect 7427 23276 7472 23304
rect 7466 23264 7472 23276
rect 7524 23264 7530 23316
rect 8665 23307 8723 23313
rect 8665 23273 8677 23307
rect 8711 23304 8723 23307
rect 9582 23304 9588 23316
rect 8711 23276 9588 23304
rect 8711 23273 8723 23276
rect 8665 23267 8723 23273
rect 9582 23264 9588 23276
rect 9640 23264 9646 23316
rect 10781 23307 10839 23313
rect 10781 23273 10793 23307
rect 10827 23304 10839 23307
rect 10962 23304 10968 23316
rect 10827 23276 10968 23304
rect 10827 23273 10839 23276
rect 10781 23267 10839 23273
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 4062 23196 4068 23248
rect 4120 23236 4126 23248
rect 5534 23236 5540 23248
rect 4120 23208 5540 23236
rect 4120 23196 4126 23208
rect 5534 23196 5540 23208
rect 5592 23236 5598 23248
rect 5766 23239 5824 23245
rect 5766 23236 5778 23239
rect 5592 23208 5778 23236
rect 5592 23196 5598 23208
rect 5766 23205 5778 23208
rect 5812 23205 5824 23239
rect 5766 23199 5824 23205
rect 7834 23196 7840 23248
rect 7892 23236 7898 23248
rect 8066 23239 8124 23245
rect 8066 23236 8078 23239
rect 7892 23208 8078 23236
rect 7892 23196 7898 23208
rect 8066 23205 8078 23208
rect 8112 23205 8124 23239
rect 8066 23199 8124 23205
rect 1464 23171 1522 23177
rect 1464 23137 1476 23171
rect 1510 23168 1522 23171
rect 2038 23168 2044 23180
rect 1510 23140 2044 23168
rect 1510 23137 1522 23140
rect 1464 23131 1522 23137
rect 2038 23128 2044 23140
rect 2096 23128 2102 23180
rect 2961 23171 3019 23177
rect 2961 23137 2973 23171
rect 3007 23168 3019 23171
rect 3050 23168 3056 23180
rect 3007 23140 3056 23168
rect 3007 23137 3019 23140
rect 2961 23131 3019 23137
rect 3050 23128 3056 23140
rect 3108 23168 3114 23180
rect 4316 23171 4374 23177
rect 3108 23140 4154 23168
rect 3108 23128 3114 23140
rect 2317 23103 2375 23109
rect 2317 23069 2329 23103
rect 2363 23100 2375 23103
rect 2590 23100 2596 23112
rect 2363 23072 2596 23100
rect 2363 23069 2375 23072
rect 2317 23063 2375 23069
rect 2590 23060 2596 23072
rect 2648 23100 2654 23112
rect 3605 23103 3663 23109
rect 3605 23100 3617 23103
rect 2648 23072 3617 23100
rect 2648 23060 2654 23072
rect 3605 23069 3617 23072
rect 3651 23100 3663 23103
rect 3970 23100 3976 23112
rect 3651 23072 3976 23100
rect 3651 23069 3663 23072
rect 3605 23063 3663 23069
rect 3970 23060 3976 23072
rect 4028 23060 4034 23112
rect 4126 23100 4154 23140
rect 4316 23137 4328 23171
rect 4362 23168 4374 23171
rect 5074 23168 5080 23180
rect 4362 23140 5080 23168
rect 4362 23137 4374 23140
rect 4316 23131 4374 23137
rect 5074 23128 5080 23140
rect 5132 23128 5138 23180
rect 8294 23168 8300 23180
rect 5368 23140 8300 23168
rect 5368 23100 5396 23140
rect 8294 23128 8300 23140
rect 8352 23168 8358 23180
rect 9398 23168 9404 23180
rect 8352 23140 9404 23168
rect 8352 23128 8358 23140
rect 9398 23128 9404 23140
rect 9456 23128 9462 23180
rect 9766 23168 9772 23180
rect 9727 23140 9772 23168
rect 9766 23128 9772 23140
rect 9824 23128 9830 23180
rect 10042 23128 10048 23180
rect 10100 23168 10106 23180
rect 10137 23171 10195 23177
rect 10137 23168 10149 23171
rect 10100 23140 10149 23168
rect 10100 23128 10106 23140
rect 10137 23137 10149 23140
rect 10183 23137 10195 23171
rect 10137 23131 10195 23137
rect 11241 23171 11299 23177
rect 11241 23137 11253 23171
rect 11287 23168 11299 23171
rect 11330 23168 11336 23180
rect 11287 23140 11336 23168
rect 11287 23137 11299 23140
rect 11241 23131 11299 23137
rect 11330 23128 11336 23140
rect 11388 23128 11394 23180
rect 4126 23072 5396 23100
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23100 5503 23103
rect 6638 23100 6644 23112
rect 5491 23072 6644 23100
rect 5491 23069 5503 23072
rect 5445 23063 5503 23069
rect 6638 23060 6644 23072
rect 6696 23060 6702 23112
rect 7742 23100 7748 23112
rect 7703 23072 7748 23100
rect 7742 23060 7748 23072
rect 7800 23060 7806 23112
rect 8570 23060 8576 23112
rect 8628 23100 8634 23112
rect 10229 23103 10287 23109
rect 10229 23100 10241 23103
rect 8628 23072 10241 23100
rect 8628 23060 8634 23072
rect 10229 23069 10241 23072
rect 10275 23069 10287 23103
rect 10229 23063 10287 23069
rect 2130 22992 2136 23044
rect 2188 23032 2194 23044
rect 2188 23004 2728 23032
rect 2188 22992 2194 23004
rect 2700 22976 2728 23004
rect 2774 22992 2780 23044
rect 2832 23032 2838 23044
rect 5994 23032 6000 23044
rect 2832 23004 6000 23032
rect 2832 22992 2838 23004
rect 5994 22992 6000 23004
rect 6052 22992 6058 23044
rect 8846 22992 8852 23044
rect 8904 23032 8910 23044
rect 11379 23035 11437 23041
rect 11379 23032 11391 23035
rect 8904 23004 11391 23032
rect 8904 22992 8910 23004
rect 11379 23001 11391 23004
rect 11425 23001 11437 23035
rect 11379 22995 11437 23001
rect 1762 22924 1768 22976
rect 1820 22964 1826 22976
rect 2041 22967 2099 22973
rect 2041 22964 2053 22967
rect 1820 22936 2053 22964
rect 1820 22924 1826 22936
rect 2041 22933 2053 22936
rect 2087 22964 2099 22967
rect 2317 22967 2375 22973
rect 2317 22964 2329 22967
rect 2087 22936 2329 22964
rect 2087 22933 2099 22936
rect 2041 22927 2099 22933
rect 2317 22933 2329 22936
rect 2363 22964 2375 22967
rect 2409 22967 2467 22973
rect 2409 22964 2421 22967
rect 2363 22936 2421 22964
rect 2363 22933 2375 22936
rect 2317 22927 2375 22933
rect 2409 22933 2421 22936
rect 2455 22933 2467 22967
rect 2409 22927 2467 22933
rect 2682 22924 2688 22976
rect 2740 22964 2746 22976
rect 3145 22967 3203 22973
rect 3145 22964 3157 22967
rect 2740 22936 3157 22964
rect 2740 22924 2746 22936
rect 3145 22933 3157 22936
rect 3191 22933 3203 22967
rect 3145 22927 3203 22933
rect 5810 22924 5816 22976
rect 5868 22964 5874 22976
rect 13262 22964 13268 22976
rect 5868 22936 13268 22964
rect 5868 22924 5874 22936
rect 13262 22924 13268 22936
rect 13320 22924 13326 22976
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 2038 22760 2044 22772
rect 1951 22732 2044 22760
rect 2038 22720 2044 22732
rect 2096 22760 2102 22772
rect 2774 22760 2780 22772
rect 2096 22732 2780 22760
rect 2096 22720 2102 22732
rect 2774 22720 2780 22732
rect 2832 22720 2838 22772
rect 3050 22760 3056 22772
rect 3011 22732 3056 22760
rect 3050 22720 3056 22732
rect 3108 22720 3114 22772
rect 3513 22763 3571 22769
rect 3513 22729 3525 22763
rect 3559 22760 3571 22763
rect 4062 22760 4068 22772
rect 3559 22732 4068 22760
rect 3559 22729 3571 22732
rect 3513 22723 3571 22729
rect 4062 22720 4068 22732
rect 4120 22760 4126 22772
rect 4430 22760 4436 22772
rect 4120 22732 4436 22760
rect 4120 22720 4126 22732
rect 4430 22720 4436 22732
rect 4488 22720 4494 22772
rect 5902 22720 5908 22772
rect 5960 22760 5966 22772
rect 7282 22760 7288 22772
rect 5960 22732 7288 22760
rect 5960 22720 5966 22732
rect 7282 22720 7288 22732
rect 7340 22720 7346 22772
rect 5534 22652 5540 22704
rect 5592 22692 5598 22704
rect 7834 22692 7840 22704
rect 5592 22664 7840 22692
rect 5592 22652 5598 22664
rect 7834 22652 7840 22664
rect 7892 22652 7898 22704
rect 10962 22692 10968 22704
rect 10060 22664 10968 22692
rect 4062 22584 4068 22636
rect 4120 22624 4126 22636
rect 4120 22596 4165 22624
rect 4120 22584 4126 22596
rect 4246 22584 4252 22636
rect 4304 22624 4310 22636
rect 4341 22627 4399 22633
rect 4341 22624 4353 22627
rect 4304 22596 4353 22624
rect 4304 22584 4310 22596
rect 4341 22593 4353 22596
rect 4387 22593 4399 22627
rect 5718 22624 5724 22636
rect 5679 22596 5724 22624
rect 4341 22587 4399 22593
rect 5718 22584 5724 22596
rect 5776 22584 5782 22636
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22624 6975 22627
rect 7006 22624 7012 22636
rect 6963 22596 7012 22624
rect 6963 22593 6975 22596
rect 6917 22587 6975 22593
rect 7006 22584 7012 22596
rect 7064 22584 7070 22636
rect 7374 22624 7380 22636
rect 7335 22596 7380 22624
rect 7374 22584 7380 22596
rect 7432 22584 7438 22636
rect 8754 22584 8760 22636
rect 8812 22624 8818 22636
rect 10060 22633 10088 22664
rect 10962 22652 10968 22664
rect 11020 22652 11026 22704
rect 8941 22627 8999 22633
rect 8941 22624 8953 22627
rect 8812 22596 8953 22624
rect 8812 22584 8818 22596
rect 8941 22593 8953 22596
rect 8987 22593 8999 22627
rect 8941 22587 8999 22593
rect 10045 22627 10103 22633
rect 10045 22593 10057 22627
rect 10091 22593 10103 22627
rect 10686 22624 10692 22636
rect 10647 22596 10692 22624
rect 10045 22587 10103 22593
rect 10686 22584 10692 22596
rect 10744 22584 10750 22636
rect 5074 22556 5080 22568
rect 4987 22528 5080 22556
rect 5074 22516 5080 22528
rect 5132 22556 5138 22568
rect 6086 22556 6092 22568
rect 5132 22528 6092 22556
rect 5132 22516 5138 22528
rect 6086 22516 6092 22528
rect 6144 22516 6150 22568
rect 8570 22556 8576 22568
rect 8531 22528 8576 22556
rect 8570 22516 8576 22528
rect 8628 22516 8634 22568
rect 8846 22556 8852 22568
rect 8807 22528 8852 22556
rect 8846 22516 8852 22528
rect 8904 22516 8910 22568
rect 4154 22488 4160 22500
rect 4126 22448 4160 22488
rect 4212 22488 4218 22500
rect 4212 22460 4257 22488
rect 4212 22448 4218 22460
rect 5902 22448 5908 22500
rect 5960 22488 5966 22500
rect 6549 22491 6607 22497
rect 6549 22488 6561 22491
rect 5960 22460 6561 22488
rect 5960 22448 5966 22460
rect 6549 22457 6561 22460
rect 6595 22488 6607 22491
rect 7009 22491 7067 22497
rect 7009 22488 7021 22491
rect 6595 22460 7021 22488
rect 6595 22457 6607 22460
rect 6549 22451 6607 22457
rect 7009 22457 7021 22460
rect 7055 22457 7067 22491
rect 7009 22451 7067 22457
rect 8662 22448 8668 22500
rect 8720 22488 8726 22500
rect 10137 22491 10195 22497
rect 10137 22488 10149 22491
rect 8720 22460 10149 22488
rect 8720 22448 8726 22460
rect 10137 22457 10149 22460
rect 10183 22488 10195 22491
rect 10502 22488 10508 22500
rect 10183 22460 10508 22488
rect 10183 22457 10195 22460
rect 10137 22451 10195 22457
rect 10502 22448 10508 22460
rect 10560 22448 10566 22500
rect 1670 22420 1676 22432
rect 1631 22392 1676 22420
rect 1670 22380 1676 22392
rect 1728 22380 1734 22432
rect 2222 22420 2228 22432
rect 2183 22392 2228 22420
rect 2222 22380 2228 22392
rect 2280 22380 2286 22432
rect 3881 22423 3939 22429
rect 3881 22389 3893 22423
rect 3927 22420 3939 22423
rect 4126 22420 4154 22448
rect 5534 22420 5540 22432
rect 3927 22392 4154 22420
rect 5495 22392 5540 22420
rect 3927 22389 3939 22392
rect 3881 22383 3939 22389
rect 5534 22380 5540 22392
rect 5592 22380 5598 22432
rect 6273 22423 6331 22429
rect 6273 22389 6285 22423
rect 6319 22420 6331 22423
rect 6638 22420 6644 22432
rect 6319 22392 6644 22420
rect 6319 22389 6331 22392
rect 6273 22383 6331 22389
rect 6638 22380 6644 22392
rect 6696 22380 6702 22432
rect 8297 22423 8355 22429
rect 8297 22389 8309 22423
rect 8343 22420 8355 22423
rect 8846 22420 8852 22432
rect 8343 22392 8852 22420
rect 8343 22389 8355 22392
rect 8297 22383 8355 22389
rect 8846 22380 8852 22392
rect 8904 22420 8910 22432
rect 9677 22423 9735 22429
rect 9677 22420 9689 22423
rect 8904 22392 9689 22420
rect 8904 22380 8910 22392
rect 9677 22389 9689 22392
rect 9723 22420 9735 22423
rect 10042 22420 10048 22432
rect 9723 22392 10048 22420
rect 9723 22389 9735 22392
rect 9677 22383 9735 22389
rect 10042 22380 10048 22392
rect 10100 22380 10106 22432
rect 11330 22420 11336 22432
rect 11243 22392 11336 22420
rect 11330 22380 11336 22392
rect 11388 22420 11394 22432
rect 12434 22420 12440 22432
rect 11388 22392 12440 22420
rect 11388 22380 11394 22392
rect 12434 22380 12440 22392
rect 12492 22380 12498 22432
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 2317 22219 2375 22225
rect 2317 22185 2329 22219
rect 2363 22216 2375 22219
rect 5534 22216 5540 22228
rect 2363 22188 2636 22216
rect 5495 22188 5540 22216
rect 2363 22185 2375 22188
rect 2317 22179 2375 22185
rect 2608 22160 2636 22188
rect 5534 22176 5540 22188
rect 5592 22176 5598 22228
rect 5626 22176 5632 22228
rect 5684 22216 5690 22228
rect 6089 22219 6147 22225
rect 6089 22216 6101 22219
rect 5684 22188 6101 22216
rect 5684 22176 5690 22188
rect 6089 22185 6101 22188
rect 6135 22185 6147 22219
rect 6089 22179 6147 22185
rect 6638 22176 6644 22228
rect 6696 22216 6702 22228
rect 7009 22219 7067 22225
rect 7009 22216 7021 22219
rect 6696 22188 7021 22216
rect 6696 22176 6702 22188
rect 7009 22185 7021 22188
rect 7055 22185 7067 22219
rect 7009 22179 7067 22185
rect 7098 22176 7104 22228
rect 7156 22216 7162 22228
rect 9815 22219 9873 22225
rect 7156 22188 8661 22216
rect 7156 22176 7162 22188
rect 1302 22108 1308 22160
rect 1360 22148 1366 22160
rect 1535 22151 1593 22157
rect 1535 22148 1547 22151
rect 1360 22120 1547 22148
rect 1360 22108 1366 22120
rect 1535 22117 1547 22120
rect 1581 22117 1593 22151
rect 1535 22111 1593 22117
rect 2222 22108 2228 22160
rect 2280 22148 2286 22160
rect 2501 22151 2559 22157
rect 2501 22148 2513 22151
rect 2280 22120 2513 22148
rect 2280 22108 2286 22120
rect 2501 22117 2513 22120
rect 2547 22117 2559 22151
rect 2501 22111 2559 22117
rect 2590 22108 2596 22160
rect 2648 22148 2654 22160
rect 7466 22148 7472 22160
rect 2648 22120 2693 22148
rect 7208 22120 7472 22148
rect 2648 22108 2654 22120
rect 1448 22083 1506 22089
rect 1448 22049 1460 22083
rect 1494 22049 1506 22083
rect 1448 22043 1506 22049
rect 4157 22083 4215 22089
rect 4157 22049 4169 22083
rect 4203 22080 4215 22083
rect 4338 22080 4344 22092
rect 4203 22052 4344 22080
rect 4203 22049 4215 22052
rect 4157 22043 4215 22049
rect 1463 22012 1491 22043
rect 4338 22040 4344 22052
rect 4396 22040 4402 22092
rect 7208 22089 7236 22120
rect 7466 22108 7472 22120
rect 7524 22108 7530 22160
rect 7193 22083 7251 22089
rect 7193 22049 7205 22083
rect 7239 22049 7251 22083
rect 7377 22083 7435 22089
rect 7377 22080 7389 22083
rect 7193 22043 7251 22049
rect 7300 22052 7389 22080
rect 1670 22012 1676 22024
rect 1463 21984 1676 22012
rect 1670 21972 1676 21984
rect 1728 22012 1734 22024
rect 3145 22015 3203 22021
rect 3145 22012 3157 22015
rect 1728 21984 3157 22012
rect 1728 21972 1734 21984
rect 3145 21981 3157 21984
rect 3191 22012 3203 22015
rect 4246 22012 4252 22024
rect 3191 21984 4252 22012
rect 3191 21981 3203 21984
rect 3145 21975 3203 21981
rect 4246 21972 4252 21984
rect 4304 21972 4310 22024
rect 5166 22012 5172 22024
rect 5127 21984 5172 22012
rect 5166 21972 5172 21984
rect 5224 21972 5230 22024
rect 7190 21904 7196 21956
rect 7248 21944 7254 21956
rect 7300 21944 7328 22052
rect 7377 22049 7389 22052
rect 7423 22049 7435 22083
rect 7377 22043 7435 22049
rect 8202 22040 8208 22092
rect 8260 22080 8266 22092
rect 8386 22080 8392 22092
rect 8260 22052 8392 22080
rect 8260 22040 8266 22052
rect 8386 22040 8392 22052
rect 8444 22080 8450 22092
rect 8516 22083 8574 22089
rect 8516 22080 8528 22083
rect 8444 22052 8528 22080
rect 8444 22040 8450 22052
rect 8516 22049 8528 22052
rect 8562 22049 8574 22083
rect 8633 22080 8661 22188
rect 9815 22185 9827 22219
rect 9861 22216 9873 22219
rect 9950 22216 9956 22228
rect 9861 22188 9956 22216
rect 9861 22185 9873 22188
rect 9815 22179 9873 22185
rect 9950 22176 9956 22188
rect 10008 22176 10014 22228
rect 10502 22216 10508 22228
rect 10463 22188 10508 22216
rect 10502 22176 10508 22188
rect 10560 22176 10566 22228
rect 9674 22080 9680 22092
rect 9732 22089 9738 22092
rect 9732 22083 9770 22089
rect 8633 22052 9680 22080
rect 8516 22043 8574 22049
rect 9674 22040 9680 22052
rect 9758 22049 9770 22083
rect 10686 22080 10692 22092
rect 10647 22052 10692 22080
rect 9732 22043 9770 22049
rect 9732 22040 9738 22043
rect 10686 22040 10692 22052
rect 10744 22040 10750 22092
rect 8619 22015 8677 22021
rect 8619 21981 8631 22015
rect 8665 22012 8677 22015
rect 9858 22012 9864 22024
rect 8665 21984 9864 22012
rect 8665 21981 8677 21984
rect 8619 21975 8677 21981
rect 9858 21972 9864 21984
rect 9916 21972 9922 22024
rect 7248 21916 7328 21944
rect 7248 21904 7254 21916
rect 10042 21904 10048 21956
rect 10100 21944 10106 21956
rect 10873 21947 10931 21953
rect 10873 21944 10885 21947
rect 10100 21916 10885 21944
rect 10100 21904 10106 21916
rect 10873 21913 10885 21916
rect 10919 21913 10931 21947
rect 10873 21907 10931 21913
rect 1762 21836 1768 21888
rect 1820 21876 1826 21888
rect 1857 21879 1915 21885
rect 1857 21876 1869 21879
rect 1820 21848 1869 21876
rect 1820 21836 1826 21848
rect 1857 21845 1869 21848
rect 1903 21845 1915 21879
rect 1857 21839 1915 21845
rect 3050 21836 3056 21888
rect 3108 21876 3114 21888
rect 4341 21879 4399 21885
rect 4341 21876 4353 21879
rect 3108 21848 4353 21876
rect 3108 21836 3114 21848
rect 4341 21845 4353 21848
rect 4387 21845 4399 21879
rect 5074 21876 5080 21888
rect 5035 21848 5080 21876
rect 4341 21839 4399 21845
rect 5074 21836 5080 21848
rect 5132 21836 5138 21888
rect 7742 21836 7748 21888
rect 7800 21876 7806 21888
rect 8021 21879 8079 21885
rect 8021 21876 8033 21879
rect 7800 21848 8033 21876
rect 7800 21836 7806 21848
rect 8021 21845 8033 21848
rect 8067 21876 8079 21879
rect 8478 21876 8484 21888
rect 8067 21848 8484 21876
rect 8067 21845 8079 21848
rect 8021 21839 8079 21845
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 8570 21836 8576 21888
rect 8628 21876 8634 21888
rect 9033 21879 9091 21885
rect 9033 21876 9045 21879
rect 8628 21848 9045 21876
rect 8628 21836 8634 21848
rect 9033 21845 9045 21848
rect 9079 21876 9091 21879
rect 9306 21876 9312 21888
rect 9079 21848 9312 21876
rect 9079 21845 9091 21848
rect 9033 21839 9091 21845
rect 9306 21836 9312 21848
rect 9364 21836 9370 21888
rect 9490 21836 9496 21888
rect 9548 21876 9554 21888
rect 9766 21876 9772 21888
rect 9548 21848 9772 21876
rect 9548 21836 9554 21848
rect 9766 21836 9772 21848
rect 9824 21876 9830 21888
rect 10137 21879 10195 21885
rect 10137 21876 10149 21879
rect 9824 21848 10149 21876
rect 9824 21836 9830 21848
rect 10137 21845 10149 21848
rect 10183 21845 10195 21879
rect 10137 21839 10195 21845
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 2222 21632 2228 21684
rect 2280 21672 2286 21684
rect 2409 21675 2467 21681
rect 2409 21672 2421 21675
rect 2280 21644 2421 21672
rect 2280 21632 2286 21644
rect 2409 21641 2421 21644
rect 2455 21641 2467 21675
rect 2409 21635 2467 21641
rect 4249 21675 4307 21681
rect 4249 21641 4261 21675
rect 4295 21672 4307 21675
rect 4338 21672 4344 21684
rect 4295 21644 4344 21672
rect 4295 21641 4307 21644
rect 4249 21635 4307 21641
rect 4338 21632 4344 21644
rect 4396 21632 4402 21684
rect 5902 21672 5908 21684
rect 5863 21644 5908 21672
rect 5902 21632 5908 21644
rect 5960 21632 5966 21684
rect 7650 21632 7656 21684
rect 7708 21672 7714 21684
rect 7837 21675 7895 21681
rect 7837 21672 7849 21675
rect 7708 21644 7849 21672
rect 7708 21632 7714 21644
rect 7837 21641 7849 21644
rect 7883 21641 7895 21675
rect 9674 21672 9680 21684
rect 9635 21644 9680 21672
rect 7837 21635 7895 21641
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 4356 21604 4384 21632
rect 7374 21604 7380 21616
rect 4356 21576 7380 21604
rect 7374 21564 7380 21576
rect 7432 21604 7438 21616
rect 7432 21576 8340 21604
rect 7432 21564 7438 21576
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 1688 21508 6561 21536
rect 1688 21480 1716 21508
rect 6549 21505 6561 21508
rect 6595 21536 6607 21539
rect 6595 21508 6868 21536
rect 6595 21505 6607 21508
rect 6549 21499 6607 21505
rect 1670 21468 1676 21480
rect 1583 21440 1676 21468
rect 1670 21428 1676 21440
rect 1728 21428 1734 21480
rect 1762 21428 1768 21480
rect 1820 21468 1826 21480
rect 1857 21471 1915 21477
rect 1857 21468 1869 21471
rect 1820 21440 1869 21468
rect 1820 21428 1826 21440
rect 1857 21437 1869 21440
rect 1903 21437 1915 21471
rect 1857 21431 1915 21437
rect 2133 21471 2191 21477
rect 2133 21437 2145 21471
rect 2179 21468 2191 21471
rect 2961 21471 3019 21477
rect 2961 21468 2973 21471
rect 2179 21440 2973 21468
rect 2179 21437 2191 21440
rect 2133 21431 2191 21437
rect 2961 21437 2973 21440
rect 3007 21468 3019 21471
rect 3142 21468 3148 21480
rect 3007 21440 3148 21468
rect 3007 21437 3019 21440
rect 2961 21431 3019 21437
rect 3142 21428 3148 21440
rect 3200 21428 3206 21480
rect 4985 21471 5043 21477
rect 4985 21437 4997 21471
rect 5031 21468 5043 21471
rect 5074 21468 5080 21480
rect 5031 21440 5080 21468
rect 5031 21437 5043 21440
rect 4985 21431 5043 21437
rect 5074 21428 5080 21440
rect 5132 21468 5138 21480
rect 5902 21468 5908 21480
rect 5132 21440 5908 21468
rect 5132 21428 5138 21440
rect 5902 21428 5908 21440
rect 5960 21428 5966 21480
rect 6840 21477 6868 21508
rect 6825 21471 6883 21477
rect 6825 21437 6837 21471
rect 6871 21437 6883 21471
rect 6825 21431 6883 21437
rect 7190 21428 7196 21480
rect 7248 21468 7254 21480
rect 7285 21471 7343 21477
rect 7285 21468 7297 21471
rect 7248 21440 7297 21468
rect 7248 21428 7254 21440
rect 7285 21437 7297 21440
rect 7331 21437 7343 21471
rect 8312 21468 8340 21576
rect 8570 21496 8576 21548
rect 8628 21536 8634 21548
rect 10686 21536 10692 21548
rect 8628 21508 10692 21536
rect 8628 21496 8634 21508
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 8389 21471 8447 21477
rect 8389 21468 8401 21471
rect 8312 21440 8401 21468
rect 7285 21431 7343 21437
rect 8389 21437 8401 21440
rect 8435 21468 8447 21471
rect 8662 21468 8668 21480
rect 8435 21440 8668 21468
rect 8435 21437 8447 21440
rect 8389 21431 8447 21437
rect 8662 21428 8668 21440
rect 8720 21428 8726 21480
rect 8846 21468 8852 21480
rect 8807 21440 8852 21468
rect 8846 21428 8852 21440
rect 8904 21428 8910 21480
rect 2866 21400 2872 21412
rect 2779 21372 2872 21400
rect 2866 21360 2872 21372
rect 2924 21400 2930 21412
rect 3323 21403 3381 21409
rect 3323 21400 3335 21403
rect 2924 21372 3335 21400
rect 2924 21360 2930 21372
rect 3323 21369 3335 21372
rect 3369 21400 3381 21403
rect 5306 21403 5364 21409
rect 3369 21372 4660 21400
rect 3369 21369 3381 21372
rect 3323 21363 3381 21369
rect 4632 21344 4660 21372
rect 5306 21369 5318 21403
rect 5352 21400 5364 21403
rect 5534 21400 5540 21412
rect 5352 21372 5540 21400
rect 5352 21369 5364 21372
rect 5306 21363 5364 21369
rect 3881 21335 3939 21341
rect 3881 21301 3893 21335
rect 3927 21332 3939 21335
rect 3970 21332 3976 21344
rect 3927 21304 3976 21332
rect 3927 21301 3939 21304
rect 3881 21295 3939 21301
rect 3970 21292 3976 21304
rect 4028 21292 4034 21344
rect 4614 21292 4620 21344
rect 4672 21332 4678 21344
rect 4801 21335 4859 21341
rect 4801 21332 4813 21335
rect 4672 21304 4813 21332
rect 4672 21292 4678 21304
rect 4801 21301 4813 21304
rect 4847 21332 4859 21335
rect 5321 21332 5349 21363
rect 5534 21360 5540 21372
rect 5592 21360 5598 21412
rect 5994 21360 6000 21412
rect 6052 21400 6058 21412
rect 9953 21403 10011 21409
rect 9953 21400 9965 21403
rect 6052 21372 9965 21400
rect 6052 21360 6058 21372
rect 9953 21369 9965 21372
rect 9999 21369 10011 21403
rect 9953 21363 10011 21369
rect 6178 21332 6184 21344
rect 4847 21304 5349 21332
rect 6139 21304 6184 21332
rect 4847 21301 4859 21304
rect 4801 21295 4859 21301
rect 6178 21292 6184 21304
rect 6236 21292 6242 21344
rect 6914 21332 6920 21344
rect 6875 21304 6920 21332
rect 6914 21292 6920 21304
rect 6972 21292 6978 21344
rect 8202 21332 8208 21344
rect 8163 21304 8208 21332
rect 8202 21292 8208 21304
rect 8260 21292 8266 21344
rect 8478 21332 8484 21344
rect 8439 21304 8484 21332
rect 8478 21292 8484 21304
rect 8536 21292 8542 21344
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 1670 21128 1676 21140
rect 1631 21100 1676 21128
rect 1670 21088 1676 21100
rect 1728 21088 1734 21140
rect 2590 21088 2596 21140
rect 2648 21128 2654 21140
rect 2961 21131 3019 21137
rect 2961 21128 2973 21131
rect 2648 21100 2973 21128
rect 2648 21088 2654 21100
rect 2961 21097 2973 21100
rect 3007 21097 3019 21131
rect 2961 21091 3019 21097
rect 3142 21088 3148 21140
rect 3200 21128 3206 21140
rect 3237 21131 3295 21137
rect 3237 21128 3249 21131
rect 3200 21100 3249 21128
rect 3200 21088 3206 21100
rect 3237 21097 3249 21100
rect 3283 21097 3295 21131
rect 3237 21091 3295 21097
rect 4154 21088 4160 21140
rect 4212 21128 4218 21140
rect 4985 21131 5043 21137
rect 4985 21128 4997 21131
rect 4212 21100 4997 21128
rect 4212 21088 4218 21100
rect 4985 21097 4997 21100
rect 5031 21097 5043 21131
rect 5902 21128 5908 21140
rect 5863 21100 5908 21128
rect 4985 21091 5043 21097
rect 5902 21088 5908 21100
rect 5960 21088 5966 21140
rect 7285 21131 7343 21137
rect 7285 21097 7297 21131
rect 7331 21128 7343 21131
rect 7466 21128 7472 21140
rect 7331 21100 7472 21128
rect 7331 21097 7343 21100
rect 7285 21091 7343 21097
rect 7466 21088 7472 21100
rect 7524 21088 7530 21140
rect 8481 21131 8539 21137
rect 8481 21097 8493 21131
rect 8527 21128 8539 21131
rect 8846 21128 8852 21140
rect 8527 21100 8852 21128
rect 8527 21097 8539 21100
rect 8481 21091 8539 21097
rect 8846 21088 8852 21100
rect 8904 21088 8910 21140
rect 2403 21063 2461 21069
rect 2403 21029 2415 21063
rect 2449 21060 2461 21063
rect 2866 21060 2872 21072
rect 2449 21032 2872 21060
rect 2449 21029 2461 21032
rect 2403 21023 2461 21029
rect 2866 21020 2872 21032
rect 2924 21020 2930 21072
rect 3789 21063 3847 21069
rect 3789 21029 3801 21063
rect 3835 21060 3847 21063
rect 4427 21063 4485 21069
rect 3835 21032 4154 21060
rect 3835 21029 3847 21032
rect 3789 21023 3847 21029
rect 4126 21004 4154 21032
rect 4427 21029 4439 21063
rect 4473 21060 4485 21063
rect 4614 21060 4620 21072
rect 4473 21032 4620 21060
rect 4473 21029 4485 21032
rect 4427 21023 4485 21029
rect 4614 21020 4620 21032
rect 4672 21020 4678 21072
rect 5166 21020 5172 21072
rect 5224 21060 5230 21072
rect 5721 21063 5779 21069
rect 5721 21060 5733 21063
rect 5224 21032 5733 21060
rect 5224 21020 5230 21032
rect 5721 21029 5733 21032
rect 5767 21060 5779 21063
rect 6914 21060 6920 21072
rect 5767 21032 6920 21060
rect 5767 21029 5779 21032
rect 5721 21023 5779 21029
rect 6914 21020 6920 21032
rect 6972 21020 6978 21072
rect 8662 21020 8668 21072
rect 8720 21060 8726 21072
rect 8757 21063 8815 21069
rect 8757 21060 8769 21063
rect 8720 21032 8769 21060
rect 8720 21020 8726 21032
rect 8757 21029 8769 21032
rect 8803 21029 8815 21063
rect 9858 21060 9864 21072
rect 9819 21032 9864 21060
rect 8757 21023 8815 21029
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 4126 20964 4160 21004
rect 4154 20952 4160 20964
rect 4212 20992 4218 21004
rect 4706 20992 4712 21004
rect 4212 20964 4712 20992
rect 4212 20952 4218 20964
rect 4706 20952 4712 20964
rect 4764 20952 4770 21004
rect 5810 20992 5816 21004
rect 5771 20964 5816 20992
rect 5810 20952 5816 20964
rect 5868 20952 5874 21004
rect 6178 20952 6184 21004
rect 6236 20992 6242 21004
rect 6365 20995 6423 21001
rect 6365 20992 6377 20995
rect 6236 20964 6377 20992
rect 6236 20952 6242 20964
rect 6365 20961 6377 20964
rect 6411 20992 6423 20995
rect 7190 20992 7196 21004
rect 6411 20964 7196 20992
rect 6411 20961 6423 20964
rect 6365 20955 6423 20961
rect 2041 20927 2099 20933
rect 2041 20893 2053 20927
rect 2087 20924 2099 20927
rect 2590 20924 2596 20936
rect 2087 20896 2596 20924
rect 2087 20893 2099 20896
rect 2041 20887 2099 20893
rect 2590 20884 2596 20896
rect 2648 20884 2654 20936
rect 4062 20924 4068 20936
rect 4023 20896 4068 20924
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 6932 20800 6960 20964
rect 7190 20952 7196 20964
rect 7248 20952 7254 21004
rect 7650 20992 7656 21004
rect 7611 20964 7656 20992
rect 7650 20952 7656 20964
rect 7708 20952 7714 21004
rect 7742 20952 7748 21004
rect 7800 20992 7806 21004
rect 7837 20995 7895 21001
rect 7837 20992 7849 20995
rect 7800 20964 7849 20992
rect 7800 20952 7806 20964
rect 7837 20961 7849 20964
rect 7883 20961 7895 20995
rect 7837 20955 7895 20961
rect 11054 20952 11060 21004
rect 11112 20992 11118 21004
rect 11241 20995 11299 21001
rect 11241 20992 11253 20995
rect 11112 20964 11253 20992
rect 11112 20952 11118 20964
rect 11241 20961 11253 20964
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 7926 20924 7932 20936
rect 7887 20896 7932 20924
rect 7926 20884 7932 20896
rect 7984 20884 7990 20936
rect 9769 20927 9827 20933
rect 9769 20893 9781 20927
rect 9815 20924 9827 20927
rect 9950 20924 9956 20936
rect 9815 20896 9956 20924
rect 9815 20893 9827 20896
rect 9769 20887 9827 20893
rect 9950 20884 9956 20896
rect 10008 20884 10014 20936
rect 10413 20927 10471 20933
rect 10413 20893 10425 20927
rect 10459 20924 10471 20927
rect 10594 20924 10600 20936
rect 10459 20896 10600 20924
rect 10459 20893 10471 20896
rect 10413 20887 10471 20893
rect 10594 20884 10600 20896
rect 10652 20884 10658 20936
rect 5350 20788 5356 20800
rect 5311 20760 5356 20788
rect 5350 20748 5356 20760
rect 5408 20748 5414 20800
rect 6914 20788 6920 20800
rect 6875 20760 6920 20788
rect 6914 20748 6920 20760
rect 6972 20748 6978 20800
rect 10410 20748 10416 20800
rect 10468 20788 10474 20800
rect 10689 20791 10747 20797
rect 10689 20788 10701 20791
rect 10468 20760 10701 20788
rect 10468 20748 10474 20760
rect 10689 20757 10701 20760
rect 10735 20757 10747 20791
rect 10689 20751 10747 20757
rect 10778 20748 10784 20800
rect 10836 20788 10842 20800
rect 11425 20791 11483 20797
rect 11425 20788 11437 20791
rect 10836 20760 11437 20788
rect 10836 20748 10842 20760
rect 11425 20757 11437 20760
rect 11471 20757 11483 20791
rect 11425 20751 11483 20757
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 2866 20584 2872 20596
rect 2827 20556 2872 20584
rect 2866 20544 2872 20556
rect 2924 20544 2930 20596
rect 4614 20544 4620 20596
rect 4672 20584 4678 20596
rect 4801 20587 4859 20593
rect 4801 20584 4813 20587
rect 4672 20556 4813 20584
rect 4672 20544 4678 20556
rect 4801 20553 4813 20556
rect 4847 20584 4859 20587
rect 5350 20584 5356 20596
rect 4847 20556 5356 20584
rect 4847 20553 4859 20556
rect 4801 20547 4859 20553
rect 5350 20544 5356 20556
rect 5408 20544 5414 20596
rect 5905 20587 5963 20593
rect 5905 20553 5917 20587
rect 5951 20584 5963 20587
rect 6638 20584 6644 20596
rect 5951 20556 6644 20584
rect 5951 20553 5963 20556
rect 5905 20547 5963 20553
rect 6638 20544 6644 20556
rect 6696 20584 6702 20596
rect 7466 20584 7472 20596
rect 6696 20556 7472 20584
rect 6696 20544 6702 20556
rect 7466 20544 7472 20556
rect 7524 20544 7530 20596
rect 9033 20587 9091 20593
rect 9033 20553 9045 20587
rect 9079 20584 9091 20587
rect 9769 20587 9827 20593
rect 9769 20584 9781 20587
rect 9079 20556 9781 20584
rect 9079 20553 9091 20556
rect 9033 20547 9091 20553
rect 9769 20553 9781 20556
rect 9815 20584 9827 20587
rect 9858 20584 9864 20596
rect 9815 20556 9864 20584
rect 9815 20553 9827 20556
rect 9769 20547 9827 20553
rect 9858 20544 9864 20556
rect 9916 20544 9922 20596
rect 4154 20516 4160 20528
rect 4126 20476 4160 20516
rect 4212 20476 4218 20528
rect 6549 20519 6607 20525
rect 6549 20485 6561 20519
rect 6595 20516 6607 20519
rect 6914 20516 6920 20528
rect 6595 20488 6920 20516
rect 6595 20485 6607 20488
rect 6549 20479 6607 20485
rect 6914 20476 6920 20488
rect 6972 20516 6978 20528
rect 12986 20516 12992 20528
rect 6972 20488 12992 20516
rect 6972 20476 6978 20488
rect 12986 20476 12992 20488
rect 13044 20476 13050 20528
rect 1762 20448 1768 20460
rect 1675 20420 1768 20448
rect 1762 20408 1768 20420
rect 1820 20448 1826 20460
rect 3789 20451 3847 20457
rect 1820 20420 2452 20448
rect 1820 20408 1826 20420
rect 1854 20380 1860 20392
rect 1815 20352 1860 20380
rect 1854 20340 1860 20352
rect 1912 20340 1918 20392
rect 2424 20389 2452 20420
rect 3789 20417 3801 20451
rect 3835 20448 3847 20451
rect 4126 20448 4154 20476
rect 4246 20448 4252 20460
rect 3835 20420 4154 20448
rect 4207 20420 4252 20448
rect 3835 20417 3847 20420
rect 3789 20411 3847 20417
rect 4246 20408 4252 20420
rect 4304 20408 4310 20460
rect 9953 20451 10011 20457
rect 9953 20417 9965 20451
rect 9999 20448 10011 20451
rect 10410 20448 10416 20460
rect 9999 20420 10416 20448
rect 9999 20417 10011 20420
rect 9953 20411 10011 20417
rect 10410 20408 10416 20420
rect 10468 20408 10474 20460
rect 2409 20383 2467 20389
rect 2409 20349 2421 20383
rect 2455 20380 2467 20383
rect 2958 20380 2964 20392
rect 2455 20352 2964 20380
rect 2455 20349 2467 20352
rect 2409 20343 2467 20349
rect 2958 20340 2964 20352
rect 3016 20340 3022 20392
rect 5629 20383 5687 20389
rect 5629 20349 5641 20383
rect 5675 20380 5687 20383
rect 5721 20383 5779 20389
rect 5721 20380 5733 20383
rect 5675 20352 5733 20380
rect 5675 20349 5687 20352
rect 5629 20343 5687 20349
rect 5721 20349 5733 20352
rect 5767 20380 5779 20383
rect 5902 20380 5908 20392
rect 5767 20352 5908 20380
rect 5767 20349 5779 20352
rect 5721 20343 5779 20349
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 7136 20383 7194 20389
rect 7136 20380 7148 20383
rect 6840 20352 7148 20380
rect 2590 20312 2596 20324
rect 2551 20284 2596 20312
rect 2590 20272 2596 20284
rect 2648 20272 2654 20324
rect 3605 20315 3663 20321
rect 3605 20281 3617 20315
rect 3651 20312 3663 20315
rect 3881 20315 3939 20321
rect 3881 20312 3893 20315
rect 3651 20284 3893 20312
rect 3651 20281 3663 20284
rect 3605 20275 3663 20281
rect 3881 20281 3893 20284
rect 3927 20312 3939 20315
rect 3970 20312 3976 20324
rect 3927 20284 3976 20312
rect 3927 20281 3939 20284
rect 3881 20275 3939 20281
rect 3970 20272 3976 20284
rect 4028 20272 4034 20324
rect 4154 20272 4160 20324
rect 4212 20312 4218 20324
rect 5810 20312 5816 20324
rect 4212 20284 5816 20312
rect 4212 20272 4218 20284
rect 5810 20272 5816 20284
rect 5868 20312 5874 20324
rect 6181 20315 6239 20321
rect 6181 20312 6193 20315
rect 5868 20284 6193 20312
rect 5868 20272 5874 20284
rect 6181 20281 6193 20284
rect 6227 20281 6239 20315
rect 6181 20275 6239 20281
rect 5534 20204 5540 20256
rect 5592 20244 5598 20256
rect 6840 20244 6868 20352
rect 7136 20349 7148 20352
rect 7182 20380 7194 20383
rect 7561 20383 7619 20389
rect 7561 20380 7573 20383
rect 7182 20352 7573 20380
rect 7182 20349 7194 20352
rect 7136 20343 7194 20349
rect 7561 20349 7573 20352
rect 7607 20380 7619 20383
rect 8018 20380 8024 20392
rect 7607 20352 8024 20380
rect 7607 20349 7619 20352
rect 7561 20343 7619 20349
rect 8018 20340 8024 20352
rect 8076 20340 8082 20392
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20380 8171 20383
rect 9309 20383 9367 20389
rect 9309 20380 9321 20383
rect 8159 20352 9321 20380
rect 8159 20349 8171 20352
rect 8113 20343 8171 20349
rect 9309 20349 9321 20352
rect 9355 20380 9367 20383
rect 9766 20380 9772 20392
rect 9355 20352 9772 20380
rect 9355 20349 9367 20352
rect 9309 20343 9367 20349
rect 9766 20340 9772 20352
rect 9824 20340 9830 20392
rect 7239 20315 7297 20321
rect 7239 20281 7251 20315
rect 7285 20312 7297 20315
rect 8294 20312 8300 20324
rect 7285 20284 8300 20312
rect 7285 20281 7297 20284
rect 7239 20275 7297 20281
rect 8294 20272 8300 20284
rect 8352 20272 8358 20324
rect 8434 20315 8492 20321
rect 8434 20281 8446 20315
rect 8480 20281 8492 20315
rect 8434 20275 8492 20281
rect 10045 20315 10103 20321
rect 10045 20281 10057 20315
rect 10091 20281 10103 20315
rect 10594 20312 10600 20324
rect 10555 20284 10600 20312
rect 10045 20275 10103 20281
rect 5592 20216 6868 20244
rect 8021 20247 8079 20253
rect 5592 20204 5598 20216
rect 8021 20213 8033 20247
rect 8067 20244 8079 20247
rect 8110 20244 8116 20256
rect 8067 20216 8116 20244
rect 8067 20213 8079 20216
rect 8021 20207 8079 20213
rect 8110 20204 8116 20216
rect 8168 20244 8174 20256
rect 8449 20244 8477 20275
rect 8168 20216 8477 20244
rect 8168 20204 8174 20216
rect 8754 20204 8760 20256
rect 8812 20244 8818 20256
rect 10060 20244 10088 20275
rect 10594 20272 10600 20284
rect 10652 20272 10658 20324
rect 10873 20247 10931 20253
rect 10873 20244 10885 20247
rect 8812 20216 10885 20244
rect 8812 20204 8818 20216
rect 10873 20213 10885 20216
rect 10919 20213 10931 20247
rect 10873 20207 10931 20213
rect 11054 20204 11060 20256
rect 11112 20244 11118 20256
rect 11241 20247 11299 20253
rect 11241 20244 11253 20247
rect 11112 20216 11253 20244
rect 11112 20204 11118 20216
rect 11241 20213 11253 20216
rect 11287 20213 11299 20247
rect 11241 20207 11299 20213
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 1578 20040 1584 20052
rect 1539 20012 1584 20040
rect 1578 20000 1584 20012
rect 1636 20000 1642 20052
rect 2590 20000 2596 20052
rect 2648 20040 2654 20052
rect 3421 20043 3479 20049
rect 3421 20040 3433 20043
rect 2648 20012 3433 20040
rect 2648 20000 2654 20012
rect 3421 20009 3433 20012
rect 3467 20009 3479 20043
rect 4890 20040 4896 20052
rect 3421 20003 3479 20009
rect 4632 20012 4896 20040
rect 3145 19975 3203 19981
rect 3145 19941 3157 19975
rect 3191 19972 3203 19975
rect 4062 19972 4068 19984
rect 3191 19944 4068 19972
rect 3191 19941 3203 19944
rect 3145 19935 3203 19941
rect 4062 19932 4068 19944
rect 4120 19972 4126 19984
rect 4632 19981 4660 20012
rect 4890 20000 4896 20012
rect 4948 20040 4954 20052
rect 5994 20040 6000 20052
rect 4948 20012 6000 20040
rect 4948 20000 4954 20012
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 8110 20000 8116 20052
rect 8168 20040 8174 20052
rect 8205 20043 8263 20049
rect 8205 20040 8217 20043
rect 8168 20012 8217 20040
rect 8168 20000 8174 20012
rect 8205 20009 8217 20012
rect 8251 20009 8263 20043
rect 8754 20040 8760 20052
rect 8715 20012 8760 20040
rect 8205 20003 8263 20009
rect 8754 20000 8760 20012
rect 8812 20000 8818 20052
rect 9766 20040 9772 20052
rect 9727 20012 9772 20040
rect 9766 20000 9772 20012
rect 9824 20000 9830 20052
rect 12986 20040 12992 20052
rect 12947 20012 12992 20040
rect 12986 20000 12992 20012
rect 13044 20000 13050 20052
rect 4249 19975 4307 19981
rect 4249 19972 4261 19975
rect 4120 19944 4261 19972
rect 4120 19932 4126 19944
rect 4249 19941 4261 19944
rect 4295 19941 4307 19975
rect 4249 19935 4307 19941
rect 4617 19975 4675 19981
rect 4617 19941 4629 19975
rect 4663 19941 4675 19975
rect 4617 19935 4675 19941
rect 4709 19975 4767 19981
rect 4709 19941 4721 19975
rect 4755 19972 4767 19975
rect 5258 19972 5264 19984
rect 4755 19944 5264 19972
rect 4755 19941 4767 19944
rect 4709 19935 4767 19941
rect 5258 19932 5264 19944
rect 5316 19932 5322 19984
rect 5350 19932 5356 19984
rect 5408 19972 5414 19984
rect 6362 19972 6368 19984
rect 5408 19944 6368 19972
rect 5408 19932 5414 19944
rect 6362 19932 6368 19944
rect 6420 19932 6426 19984
rect 8294 19932 8300 19984
rect 8352 19972 8358 19984
rect 10042 19972 10048 19984
rect 8352 19944 10048 19972
rect 8352 19932 8358 19944
rect 10042 19932 10048 19944
rect 10100 19972 10106 19984
rect 10689 19975 10747 19981
rect 10689 19972 10701 19975
rect 10100 19944 10701 19972
rect 10100 19932 10106 19944
rect 10689 19941 10701 19944
rect 10735 19941 10747 19975
rect 11422 19972 11428 19984
rect 11383 19944 11428 19972
rect 10689 19935 10747 19941
rect 11422 19932 11428 19944
rect 11480 19932 11486 19984
rect 1397 19907 1455 19913
rect 1397 19873 1409 19907
rect 1443 19904 1455 19907
rect 2685 19907 2743 19913
rect 1443 19876 2360 19904
rect 1443 19873 1455 19876
rect 1397 19867 1455 19873
rect 1854 19700 1860 19712
rect 1815 19672 1860 19700
rect 1854 19660 1860 19672
rect 1912 19660 1918 19712
rect 2332 19709 2360 19876
rect 2685 19873 2697 19907
rect 2731 19873 2743 19907
rect 2685 19867 2743 19873
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19904 2927 19907
rect 7837 19907 7895 19913
rect 2915 19876 3004 19904
rect 2915 19873 2927 19876
rect 2869 19867 2927 19873
rect 2406 19728 2412 19780
rect 2464 19768 2470 19780
rect 2700 19768 2728 19867
rect 2976 19848 3004 19876
rect 7837 19873 7849 19907
rect 7883 19904 7895 19907
rect 7926 19904 7932 19916
rect 7883 19876 7932 19904
rect 7883 19873 7895 19876
rect 7837 19867 7895 19873
rect 7926 19864 7932 19876
rect 7984 19864 7990 19916
rect 9306 19864 9312 19916
rect 9364 19904 9370 19916
rect 9674 19904 9680 19916
rect 9364 19876 9680 19904
rect 9364 19864 9370 19876
rect 9674 19864 9680 19876
rect 9732 19864 9738 19916
rect 9766 19864 9772 19916
rect 9824 19904 9830 19916
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9824 19876 10149 19904
rect 9824 19864 9830 19876
rect 10137 19873 10149 19876
rect 10183 19873 10195 19907
rect 10137 19867 10195 19873
rect 12618 19864 12624 19916
rect 12676 19904 12682 19916
rect 12805 19907 12863 19913
rect 12805 19904 12817 19907
rect 12676 19876 12817 19904
rect 12676 19864 12682 19876
rect 12805 19873 12817 19876
rect 12851 19873 12863 19907
rect 12805 19867 12863 19873
rect 2958 19796 2964 19848
rect 3016 19796 3022 19848
rect 3234 19796 3240 19848
rect 3292 19836 3298 19848
rect 4893 19839 4951 19845
rect 3292 19808 4568 19836
rect 3292 19796 3298 19808
rect 3970 19768 3976 19780
rect 2464 19740 3976 19768
rect 2464 19728 2470 19740
rect 3970 19728 3976 19740
rect 4028 19768 4034 19780
rect 4154 19768 4160 19780
rect 4028 19740 4160 19768
rect 4028 19728 4034 19740
rect 4154 19728 4160 19740
rect 4212 19728 4218 19780
rect 4540 19768 4568 19808
rect 4893 19805 4905 19839
rect 4939 19805 4951 19839
rect 4893 19799 4951 19805
rect 4908 19768 4936 19799
rect 5626 19796 5632 19848
rect 5684 19836 5690 19848
rect 6089 19839 6147 19845
rect 6089 19836 6101 19839
rect 5684 19808 6101 19836
rect 5684 19796 5690 19808
rect 6089 19805 6101 19808
rect 6135 19805 6147 19839
rect 6089 19799 6147 19805
rect 7469 19839 7527 19845
rect 7469 19805 7481 19839
rect 7515 19836 7527 19839
rect 7742 19836 7748 19848
rect 7515 19808 7748 19836
rect 7515 19805 7527 19808
rect 7469 19799 7527 19805
rect 7742 19796 7748 19808
rect 7800 19836 7806 19848
rect 9784 19836 9812 19864
rect 7800 19808 9812 19836
rect 11333 19839 11391 19845
rect 7800 19796 7806 19808
rect 11333 19805 11345 19839
rect 11379 19836 11391 19839
rect 11698 19836 11704 19848
rect 11379 19808 11704 19836
rect 11379 19805 11391 19808
rect 11333 19799 11391 19805
rect 11698 19796 11704 19808
rect 11756 19796 11762 19848
rect 10594 19768 10600 19780
rect 4540 19740 10600 19768
rect 10594 19728 10600 19740
rect 10652 19728 10658 19780
rect 11606 19728 11612 19780
rect 11664 19768 11670 19780
rect 11885 19771 11943 19777
rect 11885 19768 11897 19771
rect 11664 19740 11897 19768
rect 11664 19728 11670 19740
rect 11885 19737 11897 19740
rect 11931 19737 11943 19771
rect 11885 19731 11943 19737
rect 2317 19703 2375 19709
rect 2317 19669 2329 19703
rect 2363 19700 2375 19703
rect 4062 19700 4068 19712
rect 2363 19672 4068 19700
rect 2363 19669 2375 19672
rect 2317 19663 2375 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 5258 19660 5264 19712
rect 5316 19700 5322 19712
rect 7009 19703 7067 19709
rect 7009 19700 7021 19703
rect 5316 19672 7021 19700
rect 5316 19660 5322 19672
rect 7009 19669 7021 19672
rect 7055 19669 7067 19703
rect 7009 19663 7067 19669
rect 8018 19660 8024 19712
rect 8076 19700 8082 19712
rect 9033 19703 9091 19709
rect 9033 19700 9045 19703
rect 8076 19672 9045 19700
rect 8076 19660 8082 19672
rect 9033 19669 9045 19672
rect 9079 19669 9091 19703
rect 9033 19663 9091 19669
rect 9493 19703 9551 19709
rect 9493 19669 9505 19703
rect 9539 19700 9551 19703
rect 9950 19700 9956 19712
rect 9539 19672 9956 19700
rect 9539 19669 9551 19672
rect 9493 19663 9551 19669
rect 9950 19660 9956 19672
rect 10008 19700 10014 19712
rect 10778 19700 10784 19712
rect 10008 19672 10784 19700
rect 10008 19660 10014 19672
rect 10778 19660 10784 19672
rect 10836 19660 10842 19712
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 1762 19496 1768 19508
rect 1723 19468 1768 19496
rect 1762 19456 1768 19468
rect 1820 19456 1826 19508
rect 4890 19496 4896 19508
rect 4851 19468 4896 19496
rect 4890 19456 4896 19468
rect 4948 19456 4954 19508
rect 5258 19496 5264 19508
rect 5219 19468 5264 19496
rect 5258 19456 5264 19468
rect 5316 19456 5322 19508
rect 6638 19496 6644 19508
rect 6599 19468 6644 19496
rect 6638 19456 6644 19468
rect 6696 19456 6702 19508
rect 7101 19499 7159 19505
rect 7101 19465 7113 19499
rect 7147 19496 7159 19499
rect 7926 19496 7932 19508
rect 7147 19468 7932 19496
rect 7147 19465 7159 19468
rect 7101 19459 7159 19465
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 9950 19496 9956 19508
rect 9732 19468 9956 19496
rect 9732 19456 9738 19468
rect 9950 19456 9956 19468
rect 10008 19496 10014 19508
rect 10965 19499 11023 19505
rect 10965 19496 10977 19499
rect 10008 19468 10977 19496
rect 10008 19456 10014 19468
rect 10965 19465 10977 19468
rect 11011 19465 11023 19499
rect 11698 19496 11704 19508
rect 11659 19468 11704 19496
rect 10965 19459 11023 19465
rect 11698 19456 11704 19468
rect 11756 19496 11762 19508
rect 12575 19499 12633 19505
rect 12575 19496 12587 19499
rect 11756 19468 12587 19496
rect 11756 19456 11762 19468
rect 12575 19465 12587 19468
rect 12621 19465 12633 19499
rect 12575 19459 12633 19465
rect 1578 19388 1584 19440
rect 1636 19428 1642 19440
rect 7190 19428 7196 19440
rect 1636 19400 7196 19428
rect 1636 19388 1642 19400
rect 7190 19388 7196 19400
rect 7248 19388 7254 19440
rect 7466 19388 7472 19440
rect 7524 19428 7530 19440
rect 7524 19400 8156 19428
rect 7524 19388 7530 19400
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 3970 19360 3976 19372
rect 3375 19332 3976 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 3970 19320 3976 19332
rect 4028 19320 4034 19372
rect 6273 19363 6331 19369
rect 6273 19329 6285 19363
rect 6319 19360 6331 19363
rect 6362 19360 6368 19372
rect 6319 19332 6368 19360
rect 6319 19329 6331 19332
rect 6273 19323 6331 19329
rect 6362 19320 6368 19332
rect 6420 19360 6426 19372
rect 7484 19360 7512 19388
rect 8128 19372 8156 19400
rect 10594 19388 10600 19440
rect 10652 19428 10658 19440
rect 10652 19400 12515 19428
rect 10652 19388 10658 19400
rect 6420 19332 7512 19360
rect 7745 19363 7803 19369
rect 6420 19320 6426 19332
rect 7745 19329 7757 19363
rect 7791 19360 7803 19363
rect 7834 19360 7840 19372
rect 7791 19332 7840 19360
rect 7791 19329 7803 19332
rect 7745 19323 7803 19329
rect 2133 19295 2191 19301
rect 2133 19261 2145 19295
rect 2179 19292 2191 19295
rect 2501 19295 2559 19301
rect 2501 19292 2513 19295
rect 2179 19264 2513 19292
rect 2179 19261 2191 19264
rect 2133 19255 2191 19261
rect 2501 19261 2513 19264
rect 2547 19292 2559 19295
rect 2590 19292 2596 19304
rect 2547 19264 2596 19292
rect 2547 19261 2559 19264
rect 2501 19255 2559 19261
rect 2590 19252 2596 19264
rect 2648 19252 2654 19304
rect 2774 19292 2780 19304
rect 2735 19264 2780 19292
rect 2774 19252 2780 19264
rect 2832 19252 2838 19304
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 4798 19292 4804 19304
rect 4571 19264 4804 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 5721 19295 5779 19301
rect 5721 19261 5733 19295
rect 5767 19292 5779 19295
rect 6178 19292 6184 19304
rect 5767 19264 6184 19292
rect 5767 19261 5779 19264
rect 5721 19255 5779 19261
rect 6178 19252 6184 19264
rect 6236 19292 6242 19304
rect 6638 19292 6644 19304
rect 6236 19264 6644 19292
rect 6236 19252 6242 19264
rect 6638 19252 6644 19264
rect 6696 19252 6702 19304
rect 7260 19295 7318 19301
rect 7260 19261 7272 19295
rect 7306 19292 7318 19295
rect 7760 19292 7788 19323
rect 7834 19320 7840 19332
rect 7892 19320 7898 19372
rect 8110 19360 8116 19372
rect 8023 19332 8116 19360
rect 8110 19320 8116 19332
rect 8168 19360 8174 19372
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 8168 19332 9413 19360
rect 8168 19320 8174 19332
rect 7306 19264 7788 19292
rect 7306 19261 7318 19264
rect 7260 19255 7318 19261
rect 8018 19252 8024 19304
rect 8076 19292 8082 19304
rect 8205 19295 8263 19301
rect 8205 19292 8217 19295
rect 8076 19264 8217 19292
rect 8076 19252 8082 19264
rect 8205 19261 8217 19264
rect 8251 19261 8263 19295
rect 8205 19255 8263 19261
rect 2961 19227 3019 19233
rect 2961 19193 2973 19227
rect 3007 19224 3019 19227
rect 3418 19224 3424 19236
rect 3007 19196 3424 19224
rect 3007 19193 3019 19196
rect 2961 19187 3019 19193
rect 3418 19184 3424 19196
rect 3476 19184 3482 19236
rect 3878 19224 3884 19236
rect 3839 19196 3884 19224
rect 3878 19184 3884 19196
rect 3936 19184 3942 19236
rect 8541 19233 8569 19332
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 10042 19360 10048 19372
rect 10003 19332 10048 19360
rect 9401 19323 9459 19329
rect 10042 19320 10048 19332
rect 10100 19320 10106 19372
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19292 10747 19295
rect 10778 19292 10784 19304
rect 10735 19264 10784 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 10778 19252 10784 19264
rect 10836 19252 10842 19304
rect 11514 19252 11520 19304
rect 11572 19292 11578 19304
rect 12250 19292 12256 19304
rect 11572 19264 12256 19292
rect 11572 19252 11578 19264
rect 12250 19252 12256 19264
rect 12308 19252 12314 19304
rect 12487 19301 12515 19400
rect 12472 19295 12530 19301
rect 12472 19261 12484 19295
rect 12518 19292 12530 19295
rect 12897 19295 12955 19301
rect 12897 19292 12909 19295
rect 12518 19264 12909 19292
rect 12518 19261 12530 19264
rect 12472 19255 12530 19261
rect 12897 19261 12909 19264
rect 12943 19261 12955 19295
rect 12897 19255 12955 19261
rect 3982 19227 4040 19233
rect 3982 19193 3994 19227
rect 4028 19224 4040 19227
rect 8526 19227 8584 19233
rect 4028 19196 4108 19224
rect 4028 19193 4040 19196
rect 3982 19187 4040 19193
rect 3697 19159 3755 19165
rect 3697 19125 3709 19159
rect 3743 19156 3755 19159
rect 4080 19156 4108 19196
rect 8526 19193 8538 19227
rect 8572 19193 8584 19227
rect 8526 19187 8584 19193
rect 8754 19184 8760 19236
rect 8812 19224 8818 19236
rect 10137 19227 10195 19233
rect 10137 19224 10149 19227
rect 8812 19196 10149 19224
rect 8812 19184 8818 19196
rect 10137 19193 10149 19196
rect 10183 19224 10195 19227
rect 10502 19224 10508 19236
rect 10183 19196 10508 19224
rect 10183 19193 10195 19196
rect 10137 19187 10195 19193
rect 10502 19184 10508 19196
rect 10560 19184 10566 19236
rect 11333 19227 11391 19233
rect 11333 19224 11345 19227
rect 10796 19196 11345 19224
rect 4154 19156 4160 19168
rect 3743 19128 4160 19156
rect 3743 19125 3755 19128
rect 3697 19119 3755 19125
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 5626 19156 5632 19168
rect 5587 19128 5632 19156
rect 5626 19116 5632 19128
rect 5684 19116 5690 19168
rect 5718 19116 5724 19168
rect 5776 19156 5782 19168
rect 5905 19159 5963 19165
rect 5905 19156 5917 19159
rect 5776 19128 5917 19156
rect 5776 19116 5782 19128
rect 5905 19125 5917 19128
rect 5951 19125 5963 19159
rect 5905 19119 5963 19125
rect 7331 19159 7389 19165
rect 7331 19125 7343 19159
rect 7377 19156 7389 19159
rect 7558 19156 7564 19168
rect 7377 19128 7564 19156
rect 7377 19125 7389 19128
rect 7331 19119 7389 19125
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 9125 19159 9183 19165
rect 9125 19125 9137 19159
rect 9171 19156 9183 19159
rect 9306 19156 9312 19168
rect 9171 19128 9312 19156
rect 9171 19125 9183 19128
rect 9125 19119 9183 19125
rect 9306 19116 9312 19128
rect 9364 19116 9370 19168
rect 9766 19156 9772 19168
rect 9727 19128 9772 19156
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 10520 19156 10548 19184
rect 10796 19156 10824 19196
rect 11333 19193 11345 19196
rect 11379 19224 11391 19227
rect 11422 19224 11428 19236
rect 11379 19196 11428 19224
rect 11379 19193 11391 19196
rect 11333 19187 11391 19193
rect 11422 19184 11428 19196
rect 11480 19184 11486 19236
rect 12618 19184 12624 19236
rect 12676 19224 12682 19236
rect 13265 19227 13323 19233
rect 13265 19224 13277 19227
rect 12676 19196 13277 19224
rect 12676 19184 12682 19196
rect 13265 19193 13277 19196
rect 13311 19193 13323 19227
rect 13265 19187 13323 19193
rect 10520 19128 10824 19156
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 1670 18952 1676 18964
rect 1627 18924 1676 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 1670 18912 1676 18924
rect 1728 18912 1734 18964
rect 5626 18912 5632 18964
rect 5684 18952 5690 18964
rect 6273 18955 6331 18961
rect 6273 18952 6285 18955
rect 5684 18924 6285 18952
rect 5684 18912 5690 18924
rect 6273 18921 6285 18924
rect 6319 18921 6331 18955
rect 6273 18915 6331 18921
rect 8110 18912 8116 18964
rect 8168 18952 8174 18964
rect 8205 18955 8263 18961
rect 8205 18952 8217 18955
rect 8168 18924 8217 18952
rect 8168 18912 8174 18924
rect 8205 18921 8217 18924
rect 8251 18921 8263 18955
rect 9769 18955 9827 18961
rect 9769 18952 9781 18955
rect 8205 18915 8263 18921
rect 8680 18924 9781 18952
rect 2222 18844 2228 18896
rect 2280 18884 2286 18896
rect 3050 18884 3056 18896
rect 2280 18856 3056 18884
rect 2280 18844 2286 18856
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 2314 18816 2320 18828
rect 1443 18788 2320 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 2424 18825 2452 18856
rect 3050 18844 3056 18856
rect 3108 18844 3114 18896
rect 4522 18844 4528 18896
rect 4580 18884 4586 18896
rect 4617 18887 4675 18893
rect 4617 18884 4629 18887
rect 4580 18856 4629 18884
rect 4580 18844 4586 18856
rect 4617 18853 4629 18856
rect 4663 18853 4675 18887
rect 4617 18847 4675 18853
rect 2409 18819 2467 18825
rect 2409 18785 2421 18819
rect 2455 18785 2467 18819
rect 2774 18816 2780 18828
rect 2687 18788 2780 18816
rect 2409 18779 2467 18785
rect 1946 18748 1952 18760
rect 1907 18720 1952 18748
rect 1946 18708 1952 18720
rect 2004 18708 2010 18760
rect 2700 18748 2728 18788
rect 2774 18776 2780 18788
rect 2832 18816 2838 18828
rect 2869 18819 2927 18825
rect 2869 18816 2881 18819
rect 2832 18788 2881 18816
rect 2832 18776 2838 18788
rect 2869 18785 2881 18788
rect 2915 18785 2927 18819
rect 6178 18816 6184 18828
rect 6139 18788 6184 18816
rect 2869 18779 2927 18785
rect 6178 18776 6184 18788
rect 6236 18776 6242 18828
rect 6730 18816 6736 18828
rect 6691 18788 6736 18816
rect 6730 18776 6736 18788
rect 6788 18776 6794 18828
rect 7837 18819 7895 18825
rect 7837 18785 7849 18819
rect 7883 18816 7895 18819
rect 8478 18816 8484 18828
rect 7883 18788 8484 18816
rect 7883 18785 7895 18788
rect 7837 18779 7895 18785
rect 8478 18776 8484 18788
rect 8536 18816 8542 18828
rect 8680 18816 8708 18924
rect 9769 18921 9781 18924
rect 9815 18921 9827 18955
rect 9769 18915 9827 18921
rect 10502 18912 10508 18964
rect 10560 18952 10566 18964
rect 10689 18955 10747 18961
rect 10689 18952 10701 18955
rect 10560 18924 10701 18952
rect 10560 18912 10566 18924
rect 10689 18921 10701 18924
rect 10735 18921 10747 18955
rect 10689 18915 10747 18921
rect 10962 18884 10968 18896
rect 9692 18856 10968 18884
rect 8536 18788 8708 18816
rect 8536 18776 8542 18788
rect 8754 18776 8760 18828
rect 8812 18816 8818 18828
rect 8812 18788 8857 18816
rect 8812 18776 8818 18788
rect 9398 18776 9404 18828
rect 9456 18816 9462 18828
rect 9692 18825 9720 18856
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 11422 18884 11428 18896
rect 11383 18856 11428 18884
rect 11422 18844 11428 18856
rect 11480 18844 11486 18896
rect 9677 18819 9735 18825
rect 9677 18816 9689 18819
rect 9456 18788 9689 18816
rect 9456 18776 9462 18788
rect 9677 18785 9689 18788
rect 9723 18785 9735 18819
rect 9677 18779 9735 18785
rect 9766 18776 9772 18828
rect 9824 18816 9830 18828
rect 10137 18819 10195 18825
rect 10137 18816 10149 18819
rect 9824 18788 10149 18816
rect 9824 18776 9830 18788
rect 10137 18785 10149 18788
rect 10183 18785 10195 18819
rect 10137 18779 10195 18785
rect 12872 18819 12930 18825
rect 12872 18785 12884 18819
rect 12918 18816 12930 18819
rect 13262 18816 13268 18828
rect 12918 18788 13268 18816
rect 12918 18785 12930 18788
rect 12872 18779 12930 18785
rect 13262 18776 13268 18788
rect 13320 18776 13326 18828
rect 2958 18748 2964 18760
rect 2240 18720 2728 18748
rect 2919 18720 2964 18748
rect 2038 18572 2044 18624
rect 2096 18612 2102 18624
rect 2240 18621 2268 18720
rect 2958 18708 2964 18720
rect 3016 18708 3022 18760
rect 3881 18751 3939 18757
rect 3881 18717 3893 18751
rect 3927 18748 3939 18751
rect 3970 18748 3976 18760
rect 3927 18720 3976 18748
rect 3927 18717 3939 18720
rect 3881 18711 3939 18717
rect 3970 18708 3976 18720
rect 4028 18708 4034 18760
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18748 4583 18751
rect 4706 18748 4712 18760
rect 4571 18720 4712 18748
rect 4571 18717 4583 18720
rect 4525 18711 4583 18717
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 4798 18708 4804 18760
rect 4856 18748 4862 18760
rect 4856 18720 4901 18748
rect 4856 18708 4862 18720
rect 8754 18640 8760 18692
rect 8812 18680 8818 18692
rect 9416 18680 9444 18776
rect 10870 18708 10876 18760
rect 10928 18748 10934 18760
rect 11333 18751 11391 18757
rect 11333 18748 11345 18751
rect 10928 18720 11345 18748
rect 10928 18708 10934 18720
rect 11333 18717 11345 18720
rect 11379 18717 11391 18751
rect 11333 18711 11391 18717
rect 11609 18751 11667 18757
rect 11609 18717 11621 18751
rect 11655 18717 11667 18751
rect 11609 18711 11667 18717
rect 8812 18652 9444 18680
rect 8812 18640 8818 18652
rect 10410 18640 10416 18692
rect 10468 18680 10474 18692
rect 11514 18680 11520 18692
rect 10468 18652 11520 18680
rect 10468 18640 10474 18652
rect 11514 18640 11520 18652
rect 11572 18680 11578 18692
rect 11624 18680 11652 18711
rect 11572 18652 11652 18680
rect 11572 18640 11578 18652
rect 2225 18615 2283 18621
rect 2225 18612 2237 18615
rect 2096 18584 2237 18612
rect 2096 18572 2102 18584
rect 2225 18581 2237 18584
rect 2271 18581 2283 18615
rect 2225 18575 2283 18581
rect 8846 18572 8852 18624
rect 8904 18612 8910 18624
rect 9033 18615 9091 18621
rect 9033 18612 9045 18615
rect 8904 18584 9045 18612
rect 8904 18572 8910 18584
rect 9033 18581 9045 18584
rect 9079 18581 9091 18615
rect 9033 18575 9091 18581
rect 11330 18572 11336 18624
rect 11388 18612 11394 18624
rect 12943 18615 13001 18621
rect 12943 18612 12955 18615
rect 11388 18584 12955 18612
rect 11388 18572 11394 18584
rect 12943 18581 12955 18584
rect 12989 18581 13001 18615
rect 12943 18575 13001 18581
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 2041 18411 2099 18417
rect 2041 18377 2053 18411
rect 2087 18408 2099 18411
rect 2406 18408 2412 18420
rect 2087 18380 2412 18408
rect 2087 18377 2099 18380
rect 2041 18371 2099 18377
rect 2406 18368 2412 18380
rect 2464 18368 2470 18420
rect 3789 18411 3847 18417
rect 3789 18377 3801 18411
rect 3835 18408 3847 18411
rect 4154 18408 4160 18420
rect 3835 18380 4160 18408
rect 3835 18377 3847 18380
rect 3789 18371 3847 18377
rect 4154 18368 4160 18380
rect 4212 18408 4218 18420
rect 4798 18408 4804 18420
rect 4212 18380 4804 18408
rect 4212 18368 4218 18380
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 6178 18368 6184 18420
rect 6236 18408 6242 18420
rect 6549 18411 6607 18417
rect 6549 18408 6561 18411
rect 6236 18380 6561 18408
rect 6236 18368 6242 18380
rect 6549 18377 6561 18380
rect 6595 18377 6607 18411
rect 6549 18371 6607 18377
rect 7331 18411 7389 18417
rect 7331 18377 7343 18411
rect 7377 18408 7389 18411
rect 10870 18408 10876 18420
rect 7377 18380 10876 18408
rect 7377 18377 7389 18380
rect 7331 18371 7389 18377
rect 10870 18368 10876 18380
rect 10928 18408 10934 18420
rect 12069 18411 12127 18417
rect 12069 18408 12081 18411
rect 10928 18380 12081 18408
rect 10928 18368 10934 18380
rect 12069 18377 12081 18380
rect 12115 18377 12127 18411
rect 13262 18408 13268 18420
rect 13223 18380 13268 18408
rect 12069 18371 12127 18377
rect 13262 18368 13268 18380
rect 13320 18368 13326 18420
rect 1762 18300 1768 18352
rect 1820 18340 1826 18352
rect 5534 18340 5540 18352
rect 1820 18312 5540 18340
rect 1820 18300 1826 18312
rect 5534 18300 5540 18312
rect 5592 18300 5598 18352
rect 6273 18343 6331 18349
rect 6273 18309 6285 18343
rect 6319 18340 6331 18343
rect 6730 18340 6736 18352
rect 6319 18312 6736 18340
rect 6319 18309 6331 18312
rect 6273 18303 6331 18309
rect 6730 18300 6736 18312
rect 6788 18300 6794 18352
rect 7101 18343 7159 18349
rect 7101 18309 7113 18343
rect 7147 18340 7159 18343
rect 7466 18340 7472 18352
rect 7147 18312 7472 18340
rect 7147 18309 7159 18312
rect 7101 18303 7159 18309
rect 7466 18300 7472 18312
rect 7524 18340 7530 18352
rect 8021 18343 8079 18349
rect 8021 18340 8033 18343
rect 7524 18312 8033 18340
rect 7524 18300 7530 18312
rect 8021 18309 8033 18312
rect 8067 18340 8079 18343
rect 8386 18340 8392 18352
rect 8067 18312 8392 18340
rect 8067 18309 8079 18312
rect 8021 18303 8079 18309
rect 8386 18300 8392 18312
rect 8444 18300 8450 18352
rect 9125 18343 9183 18349
rect 9125 18309 9137 18343
rect 9171 18340 9183 18343
rect 11333 18343 11391 18349
rect 11333 18340 11345 18343
rect 9171 18312 11345 18340
rect 9171 18309 9183 18312
rect 9125 18303 9183 18309
rect 11333 18309 11345 18312
rect 11379 18340 11391 18343
rect 11422 18340 11428 18352
rect 11379 18312 11428 18340
rect 11379 18309 11391 18312
rect 11333 18303 11391 18309
rect 11422 18300 11428 18312
rect 11480 18300 11486 18352
rect 2869 18275 2927 18281
rect 2869 18241 2881 18275
rect 2915 18272 2927 18275
rect 2958 18272 2964 18284
rect 2915 18244 2964 18272
rect 2915 18241 2927 18244
rect 2869 18235 2927 18241
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 4706 18232 4712 18284
rect 4764 18272 4770 18284
rect 5721 18275 5779 18281
rect 5721 18272 5733 18275
rect 4764 18244 5733 18272
rect 4764 18232 4770 18244
rect 5721 18241 5733 18244
rect 5767 18272 5779 18275
rect 5767 18244 7788 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 1857 18207 1915 18213
rect 1857 18173 1869 18207
rect 1903 18204 1915 18207
rect 1946 18204 1952 18216
rect 1903 18176 1952 18204
rect 1903 18173 1915 18176
rect 1857 18167 1915 18173
rect 1946 18164 1952 18176
rect 2004 18164 2010 18216
rect 5353 18207 5411 18213
rect 5353 18173 5365 18207
rect 5399 18204 5411 18207
rect 6178 18204 6184 18216
rect 5399 18176 6184 18204
rect 5399 18173 5411 18176
rect 5353 18167 5411 18173
rect 6178 18164 6184 18176
rect 6236 18164 6242 18216
rect 7260 18207 7318 18213
rect 7260 18173 7272 18207
rect 7306 18173 7318 18207
rect 7760 18204 7788 18244
rect 8110 18232 8116 18284
rect 8168 18272 8174 18284
rect 8205 18275 8263 18281
rect 8205 18272 8217 18275
rect 8168 18244 8217 18272
rect 8168 18232 8174 18244
rect 8205 18241 8217 18244
rect 8251 18272 8263 18275
rect 8846 18272 8852 18284
rect 8251 18244 8852 18272
rect 8251 18241 8263 18244
rect 8205 18235 8263 18241
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18272 10103 18275
rect 10686 18272 10692 18284
rect 10091 18244 10692 18272
rect 10091 18241 10103 18244
rect 10045 18235 10103 18241
rect 10686 18232 10692 18244
rect 10744 18272 10750 18284
rect 11701 18275 11759 18281
rect 11701 18272 11713 18275
rect 10744 18244 11713 18272
rect 10744 18232 10750 18244
rect 11701 18241 11713 18244
rect 11747 18241 11759 18275
rect 11701 18235 11759 18241
rect 12066 18232 12072 18284
rect 12124 18272 12130 18284
rect 13906 18272 13912 18284
rect 12124 18244 13912 18272
rect 12124 18232 12130 18244
rect 9766 18204 9772 18216
rect 7760 18176 9772 18204
rect 7260 18167 7318 18173
rect 3190 18139 3248 18145
rect 3190 18136 3202 18139
rect 2792 18108 3202 18136
rect 2792 18080 2820 18108
rect 3190 18105 3202 18108
rect 3236 18105 3248 18139
rect 4706 18136 4712 18148
rect 4667 18108 4712 18136
rect 3190 18099 3248 18105
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 4798 18096 4804 18148
rect 4856 18136 4862 18148
rect 7275 18136 7303 18167
rect 9766 18164 9772 18176
rect 9824 18164 9830 18216
rect 10870 18204 10876 18216
rect 10704 18176 10876 18204
rect 7745 18139 7803 18145
rect 7745 18136 7757 18139
rect 4856 18108 4901 18136
rect 7275 18108 7757 18136
rect 4856 18096 4862 18108
rect 7745 18105 7757 18108
rect 7791 18136 7803 18139
rect 7791 18108 8156 18136
rect 7791 18105 7803 18108
rect 7745 18099 7803 18105
rect 1765 18071 1823 18077
rect 1765 18037 1777 18071
rect 1811 18068 1823 18071
rect 1946 18068 1952 18080
rect 1811 18040 1952 18068
rect 1811 18037 1823 18040
rect 1765 18031 1823 18037
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 2222 18028 2228 18080
rect 2280 18068 2286 18080
rect 2317 18071 2375 18077
rect 2317 18068 2329 18071
rect 2280 18040 2329 18068
rect 2280 18028 2286 18040
rect 2317 18037 2329 18040
rect 2363 18037 2375 18071
rect 2774 18068 2780 18080
rect 2735 18040 2780 18068
rect 2317 18031 2375 18037
rect 2774 18028 2780 18040
rect 2832 18028 2838 18080
rect 4522 18068 4528 18080
rect 4483 18040 4528 18068
rect 4522 18028 4528 18040
rect 4580 18028 4586 18080
rect 8128 18068 8156 18108
rect 8386 18096 8392 18148
rect 8444 18136 8450 18148
rect 8526 18139 8584 18145
rect 8526 18136 8538 18139
rect 8444 18108 8538 18136
rect 8444 18096 8450 18108
rect 8526 18105 8538 18108
rect 8572 18105 8584 18139
rect 8526 18099 8584 18105
rect 9306 18096 9312 18148
rect 9364 18136 9370 18148
rect 9858 18136 9864 18148
rect 9364 18108 9864 18136
rect 9364 18096 9370 18108
rect 9858 18096 9864 18108
rect 9916 18136 9922 18148
rect 10704 18145 10732 18176
rect 10870 18164 10876 18176
rect 10928 18164 10934 18216
rect 10962 18164 10968 18216
rect 11020 18204 11026 18216
rect 12342 18204 12348 18216
rect 11020 18176 11065 18204
rect 12084 18176 12348 18204
rect 11020 18164 11026 18176
rect 12084 18148 12112 18176
rect 12342 18164 12348 18176
rect 12400 18204 12406 18216
rect 13531 18213 13559 18244
rect 13906 18232 13912 18244
rect 13964 18232 13970 18284
rect 12472 18207 12530 18213
rect 12472 18204 12484 18207
rect 12400 18176 12484 18204
rect 12400 18164 12406 18176
rect 12472 18173 12484 18176
rect 12518 18204 12530 18207
rect 12897 18207 12955 18213
rect 12897 18204 12909 18207
rect 12518 18176 12909 18204
rect 12518 18173 12530 18176
rect 12472 18167 12530 18173
rect 12897 18173 12909 18176
rect 12943 18173 12955 18207
rect 13516 18207 13574 18213
rect 13516 18204 13528 18207
rect 13494 18176 13528 18204
rect 12897 18167 12955 18173
rect 13516 18173 13528 18176
rect 13562 18173 13574 18207
rect 13516 18167 13574 18173
rect 10137 18139 10195 18145
rect 10137 18136 10149 18139
rect 9916 18108 10149 18136
rect 9916 18096 9922 18108
rect 10137 18105 10149 18108
rect 10183 18105 10195 18139
rect 10137 18099 10195 18105
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18105 10747 18139
rect 10689 18099 10747 18105
rect 10796 18108 11468 18136
rect 8202 18068 8208 18080
rect 8128 18040 8208 18068
rect 8202 18028 8208 18040
rect 8260 18068 8266 18080
rect 9398 18068 9404 18080
rect 8260 18040 9404 18068
rect 8260 18028 8266 18040
rect 9398 18028 9404 18040
rect 9456 18028 9462 18080
rect 9674 18068 9680 18080
rect 9635 18040 9680 18068
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10796 18068 10824 18108
rect 9824 18040 10824 18068
rect 11440 18068 11468 18108
rect 12066 18096 12072 18148
rect 12124 18096 12130 18148
rect 12575 18071 12633 18077
rect 12575 18068 12587 18071
rect 11440 18040 12587 18068
rect 9824 18028 9830 18040
rect 12575 18037 12587 18040
rect 12621 18037 12633 18071
rect 12575 18031 12633 18037
rect 13354 18028 13360 18080
rect 13412 18068 13418 18080
rect 13587 18071 13645 18077
rect 13587 18068 13599 18071
rect 13412 18040 13599 18068
rect 13412 18028 13418 18040
rect 13587 18037 13599 18040
rect 13633 18037 13645 18071
rect 13906 18068 13912 18080
rect 13867 18040 13912 18068
rect 13587 18031 13645 18037
rect 13906 18028 13912 18040
rect 13964 18028 13970 18080
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 2958 17824 2964 17876
rect 3016 17864 3022 17876
rect 3329 17867 3387 17873
rect 3329 17864 3341 17867
rect 3016 17836 3341 17864
rect 3016 17824 3022 17836
rect 3329 17833 3341 17836
rect 3375 17833 3387 17867
rect 3329 17827 3387 17833
rect 4338 17824 4344 17876
rect 4396 17864 4402 17876
rect 4433 17867 4491 17873
rect 4433 17864 4445 17867
rect 4396 17836 4445 17864
rect 4396 17824 4402 17836
rect 4433 17833 4445 17836
rect 4479 17833 4491 17867
rect 4433 17827 4491 17833
rect 2133 17799 2191 17805
rect 2133 17765 2145 17799
rect 2179 17796 2191 17799
rect 2682 17796 2688 17808
rect 2179 17768 2688 17796
rect 2179 17765 2191 17768
rect 2133 17759 2191 17765
rect 2682 17756 2688 17768
rect 2740 17796 2746 17808
rect 3697 17799 3755 17805
rect 3697 17796 3709 17799
rect 2740 17768 3709 17796
rect 2740 17756 2746 17768
rect 3697 17765 3709 17768
rect 3743 17765 3755 17799
rect 4448 17796 4476 17827
rect 4522 17824 4528 17876
rect 4580 17864 4586 17876
rect 4985 17867 5043 17873
rect 4985 17864 4997 17867
rect 4580 17836 4997 17864
rect 4580 17824 4586 17836
rect 4985 17833 4997 17836
rect 5031 17833 5043 17867
rect 8478 17864 8484 17876
rect 8439 17836 8484 17864
rect 4985 17827 5043 17833
rect 4614 17796 4620 17808
rect 4448 17768 4620 17796
rect 3697 17759 3755 17765
rect 4614 17756 4620 17768
rect 4672 17756 4678 17808
rect 5000 17796 5028 17827
rect 8478 17824 8484 17836
rect 8536 17824 8542 17876
rect 9582 17824 9588 17876
rect 9640 17864 9646 17876
rect 9640 17836 12915 17864
rect 9640 17824 9646 17836
rect 5994 17796 6000 17808
rect 5000 17768 6000 17796
rect 5994 17756 6000 17768
rect 6052 17756 6058 17808
rect 8110 17796 8116 17808
rect 8071 17768 8116 17796
rect 8110 17756 8116 17768
rect 8168 17756 8174 17808
rect 8386 17756 8392 17808
rect 8444 17796 8450 17808
rect 9490 17796 9496 17808
rect 8444 17768 9496 17796
rect 8444 17756 8450 17768
rect 9490 17756 9496 17768
rect 9548 17756 9554 17808
rect 9858 17796 9864 17808
rect 9819 17768 9864 17796
rect 9858 17756 9864 17768
rect 9916 17796 9922 17808
rect 10689 17799 10747 17805
rect 10689 17796 10701 17799
rect 9916 17768 10701 17796
rect 9916 17756 9922 17768
rect 10689 17765 10701 17768
rect 10735 17765 10747 17799
rect 11330 17796 11336 17808
rect 11291 17768 11336 17796
rect 10689 17759 10747 17765
rect 11330 17756 11336 17768
rect 11388 17756 11394 17808
rect 11422 17756 11428 17808
rect 11480 17796 11486 17808
rect 11480 17768 11525 17796
rect 11480 17756 11486 17768
rect 3418 17688 3424 17740
rect 3476 17728 3482 17740
rect 4065 17731 4123 17737
rect 4065 17728 4077 17731
rect 3476 17700 4077 17728
rect 3476 17688 3482 17700
rect 4065 17697 4077 17700
rect 4111 17697 4123 17731
rect 7374 17728 7380 17740
rect 7335 17700 7380 17728
rect 4065 17691 4123 17697
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 7834 17688 7840 17740
rect 7892 17728 7898 17740
rect 7929 17731 7987 17737
rect 7929 17728 7941 17731
rect 7892 17700 7941 17728
rect 7892 17688 7898 17700
rect 7929 17697 7941 17700
rect 7975 17728 7987 17731
rect 9582 17728 9588 17740
rect 7975 17700 9588 17728
rect 7975 17697 7987 17700
rect 7929 17691 7987 17697
rect 9582 17688 9588 17700
rect 9640 17688 9646 17740
rect 10410 17688 10416 17740
rect 10468 17728 10474 17740
rect 12887 17737 12915 17836
rect 12872 17731 12930 17737
rect 10468 17700 10513 17728
rect 10468 17688 10474 17700
rect 12872 17697 12884 17731
rect 12918 17728 12930 17731
rect 13262 17728 13268 17740
rect 12918 17700 13268 17728
rect 12918 17697 12930 17700
rect 12872 17691 12930 17697
rect 13262 17688 13268 17700
rect 13320 17688 13326 17740
rect 2038 17660 2044 17672
rect 1999 17632 2044 17660
rect 2038 17620 2044 17632
rect 2096 17620 2102 17672
rect 2314 17620 2320 17672
rect 2372 17660 2378 17672
rect 2961 17663 3019 17669
rect 2961 17660 2973 17663
rect 2372 17632 2973 17660
rect 2372 17620 2378 17632
rect 2961 17629 2973 17632
rect 3007 17660 3019 17663
rect 5626 17660 5632 17672
rect 3007 17632 5632 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 5626 17620 5632 17632
rect 5684 17620 5690 17672
rect 5721 17663 5779 17669
rect 5721 17629 5733 17663
rect 5767 17660 5779 17663
rect 5905 17663 5963 17669
rect 5905 17660 5917 17663
rect 5767 17632 5917 17660
rect 5767 17629 5779 17632
rect 5721 17623 5779 17629
rect 5905 17629 5917 17632
rect 5951 17629 5963 17663
rect 6178 17660 6184 17672
rect 6139 17632 6184 17660
rect 5905 17623 5963 17629
rect 2593 17595 2651 17601
rect 2593 17561 2605 17595
rect 2639 17561 2651 17595
rect 5920 17592 5948 17623
rect 6178 17620 6184 17632
rect 6236 17620 6242 17672
rect 7558 17620 7564 17672
rect 7616 17660 7622 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 7616 17632 9781 17660
rect 7616 17620 7622 17632
rect 9769 17629 9781 17632
rect 9815 17660 9827 17663
rect 10042 17660 10048 17672
rect 9815 17632 10048 17660
rect 9815 17629 9827 17632
rect 9769 17623 9827 17629
rect 10042 17620 10048 17632
rect 10100 17620 10106 17672
rect 13354 17660 13360 17672
rect 10152 17632 13360 17660
rect 10152 17592 10180 17632
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 5920 17564 10180 17592
rect 2593 17555 2651 17561
rect 1673 17527 1731 17533
rect 1673 17493 1685 17527
rect 1719 17524 1731 17527
rect 1946 17524 1952 17536
rect 1719 17496 1952 17524
rect 1719 17493 1731 17496
rect 1673 17487 1731 17493
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 2314 17484 2320 17536
rect 2372 17524 2378 17536
rect 2608 17524 2636 17555
rect 10870 17552 10876 17604
rect 10928 17592 10934 17604
rect 11885 17595 11943 17601
rect 11885 17592 11897 17595
rect 10928 17564 11897 17592
rect 10928 17552 10934 17564
rect 11885 17561 11897 17564
rect 11931 17561 11943 17595
rect 11885 17555 11943 17561
rect 2372 17496 2636 17524
rect 2372 17484 2378 17496
rect 4706 17484 4712 17536
rect 4764 17524 4770 17536
rect 5353 17527 5411 17533
rect 5353 17524 5365 17527
rect 4764 17496 5365 17524
rect 4764 17484 4770 17496
rect 5353 17493 5365 17496
rect 5399 17524 5411 17527
rect 7374 17524 7380 17536
rect 5399 17496 7380 17524
rect 5399 17493 5411 17496
rect 5353 17487 5411 17493
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 8941 17527 8999 17533
rect 8941 17493 8953 17527
rect 8987 17524 8999 17527
rect 9306 17524 9312 17536
rect 8987 17496 9312 17524
rect 8987 17493 8999 17496
rect 8941 17487 8999 17493
rect 9306 17484 9312 17496
rect 9364 17484 9370 17536
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 12943 17527 13001 17533
rect 12943 17524 12955 17527
rect 10836 17496 12955 17524
rect 10836 17484 10842 17496
rect 12943 17493 12955 17496
rect 12989 17493 13001 17527
rect 12943 17487 13001 17493
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 2593 17323 2651 17329
rect 2593 17289 2605 17323
rect 2639 17320 2651 17323
rect 5718 17320 5724 17332
rect 2639 17292 5724 17320
rect 2639 17289 2651 17292
rect 2593 17283 2651 17289
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 5994 17320 6000 17332
rect 5955 17292 6000 17320
rect 5994 17280 6000 17292
rect 6052 17280 6058 17332
rect 9858 17320 9864 17332
rect 9819 17292 9864 17320
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 10042 17280 10048 17332
rect 10100 17320 10106 17332
rect 10229 17323 10287 17329
rect 10229 17320 10241 17323
rect 10100 17292 10241 17320
rect 10100 17280 10106 17292
rect 10229 17289 10241 17292
rect 10275 17289 10287 17323
rect 10229 17283 10287 17289
rect 11330 17280 11336 17332
rect 11388 17320 11394 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11388 17292 11621 17320
rect 11388 17280 11394 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 13262 17320 13268 17332
rect 13223 17292 13268 17320
rect 11609 17283 11667 17289
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 6638 17212 6644 17264
rect 6696 17252 6702 17264
rect 13587 17255 13645 17261
rect 13587 17252 13599 17255
rect 6696 17224 13599 17252
rect 6696 17212 6702 17224
rect 13587 17221 13599 17224
rect 13633 17221 13645 17255
rect 13587 17215 13645 17221
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17184 6607 17187
rect 6730 17184 6736 17196
rect 6595 17156 6736 17184
rect 6595 17153 6607 17156
rect 6549 17147 6607 17153
rect 6730 17144 6736 17156
rect 6788 17184 6794 17196
rect 7193 17187 7251 17193
rect 7193 17184 7205 17187
rect 6788 17156 7205 17184
rect 6788 17144 6794 17156
rect 7193 17153 7205 17156
rect 7239 17184 7251 17187
rect 8018 17184 8024 17196
rect 7239 17156 7880 17184
rect 7979 17156 8024 17184
rect 7239 17153 7251 17156
rect 7193 17147 7251 17153
rect 7852 17128 7880 17156
rect 8018 17144 8024 17156
rect 8076 17144 8082 17196
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17184 8815 17187
rect 8941 17187 8999 17193
rect 8941 17184 8953 17187
rect 8803 17156 8953 17184
rect 8803 17153 8815 17156
rect 8757 17147 8815 17153
rect 8941 17153 8953 17156
rect 8987 17184 8999 17187
rect 9214 17184 9220 17196
rect 8987 17156 9220 17184
rect 8987 17153 8999 17156
rect 8941 17147 8999 17153
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 10551 17187 10609 17193
rect 10551 17153 10563 17187
rect 10597 17184 10609 17187
rect 10686 17184 10692 17196
rect 10597 17156 10692 17184
rect 10597 17153 10609 17156
rect 10551 17147 10609 17153
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 11333 17187 11391 17193
rect 11333 17153 11345 17187
rect 11379 17184 11391 17187
rect 11422 17184 11428 17196
rect 11379 17156 11428 17184
rect 11379 17153 11391 17156
rect 11333 17147 11391 17153
rect 11422 17144 11428 17156
rect 11480 17144 11486 17196
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17085 1731 17119
rect 1946 17116 1952 17128
rect 1907 17088 1952 17116
rect 1673 17079 1731 17085
rect 1688 17048 1716 17079
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 2961 17119 3019 17125
rect 2961 17085 2973 17119
rect 3007 17116 3019 17119
rect 3142 17116 3148 17128
rect 3007 17088 3148 17116
rect 3007 17085 3019 17088
rect 2961 17079 3019 17085
rect 3142 17076 3148 17088
rect 3200 17076 3206 17128
rect 4798 17116 4804 17128
rect 4759 17088 4804 17116
rect 4798 17076 4804 17088
rect 4856 17076 4862 17128
rect 5810 17076 5816 17128
rect 5868 17116 5874 17128
rect 6822 17116 6828 17128
rect 5868 17088 6828 17116
rect 5868 17076 5874 17088
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 7558 17116 7564 17128
rect 7519 17088 7564 17116
rect 7558 17076 7564 17088
rect 7616 17076 7622 17128
rect 7834 17116 7840 17128
rect 7795 17088 7840 17116
rect 7834 17076 7840 17088
rect 7892 17076 7898 17128
rect 8662 17076 8668 17128
rect 8720 17116 8726 17128
rect 8849 17119 8907 17125
rect 8849 17116 8861 17119
rect 8720 17088 8861 17116
rect 8720 17076 8726 17088
rect 8849 17085 8861 17088
rect 8895 17085 8907 17119
rect 8849 17079 8907 17085
rect 9125 17119 9183 17125
rect 9125 17085 9137 17119
rect 9171 17116 9183 17119
rect 9306 17116 9312 17128
rect 9171 17088 9312 17116
rect 9171 17085 9183 17088
rect 9125 17079 9183 17085
rect 9306 17076 9312 17088
rect 9364 17116 9370 17128
rect 9950 17116 9956 17128
rect 9364 17088 9956 17116
rect 9364 17076 9370 17088
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 10464 17119 10522 17125
rect 10464 17085 10476 17119
rect 10510 17116 10522 17119
rect 10870 17116 10876 17128
rect 10510 17088 10876 17116
rect 10510 17085 10522 17088
rect 10464 17079 10522 17085
rect 10870 17076 10876 17088
rect 10928 17076 10934 17128
rect 12158 17076 12164 17128
rect 12216 17116 12222 17128
rect 12472 17119 12530 17125
rect 12472 17116 12484 17119
rect 12216 17088 12484 17116
rect 12216 17076 12222 17088
rect 12472 17085 12484 17088
rect 12518 17116 12530 17119
rect 12894 17116 12900 17128
rect 12518 17088 12900 17116
rect 12518 17085 12530 17088
rect 12472 17079 12530 17085
rect 12894 17076 12900 17088
rect 12952 17076 12958 17128
rect 13516 17119 13574 17125
rect 13516 17085 13528 17119
rect 13562 17116 13574 17119
rect 13722 17116 13728 17128
rect 13562 17088 13728 17116
rect 13562 17085 13574 17088
rect 13516 17079 13574 17085
rect 13722 17076 13728 17088
rect 13780 17116 13786 17128
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13780 17088 13921 17116
rect 13780 17076 13786 17088
rect 13909 17085 13921 17088
rect 13955 17085 13967 17119
rect 13909 17079 13967 17085
rect 1688 17020 1900 17048
rect 1872 16992 1900 17020
rect 2130 17008 2136 17060
rect 2188 17048 2194 17060
rect 2774 17048 2780 17060
rect 2188 17020 2780 17048
rect 2188 17008 2194 17020
rect 2774 17008 2780 17020
rect 2832 17048 2838 17060
rect 3282 17051 3340 17057
rect 3282 17048 3294 17051
rect 2832 17020 3294 17048
rect 2832 17008 2838 17020
rect 3282 17017 3294 17020
rect 3328 17048 3340 17051
rect 4157 17051 4215 17057
rect 4157 17048 4169 17051
rect 3328 17020 4169 17048
rect 3328 17017 3340 17020
rect 3282 17011 3340 17017
rect 4157 17017 4169 17020
rect 4203 17048 4215 17051
rect 4338 17048 4344 17060
rect 4203 17020 4344 17048
rect 4203 17017 4215 17020
rect 4157 17011 4215 17017
rect 4338 17008 4344 17020
rect 4396 17048 4402 17060
rect 4617 17051 4675 17057
rect 4617 17048 4629 17051
rect 4396 17020 4629 17048
rect 4396 17008 4402 17020
rect 4617 17017 4629 17020
rect 4663 17048 4675 17051
rect 5122 17051 5180 17057
rect 5122 17048 5134 17051
rect 4663 17020 5134 17048
rect 4663 17017 4675 17020
rect 4617 17011 4675 17017
rect 5122 17017 5134 17020
rect 5168 17017 5180 17051
rect 5122 17011 5180 17017
rect 5534 17008 5540 17060
rect 5592 17048 5598 17060
rect 12575 17051 12633 17057
rect 12575 17048 12587 17051
rect 5592 17020 12587 17048
rect 5592 17008 5598 17020
rect 12575 17017 12587 17020
rect 12621 17017 12633 17051
rect 12575 17011 12633 17017
rect 1670 16980 1676 16992
rect 1631 16952 1676 16980
rect 1670 16940 1676 16952
rect 1728 16940 1734 16992
rect 1854 16940 1860 16992
rect 1912 16980 1918 16992
rect 2409 16983 2467 16989
rect 2409 16980 2421 16983
rect 1912 16952 2421 16980
rect 1912 16940 1918 16952
rect 2409 16949 2421 16952
rect 2455 16980 2467 16983
rect 2593 16983 2651 16989
rect 2593 16980 2605 16983
rect 2455 16952 2605 16980
rect 2455 16949 2467 16952
rect 2409 16943 2467 16949
rect 2593 16949 2605 16952
rect 2639 16949 2651 16983
rect 3878 16980 3884 16992
rect 3839 16952 3884 16980
rect 2593 16943 2651 16949
rect 3878 16940 3884 16952
rect 3936 16940 3942 16992
rect 5718 16980 5724 16992
rect 5679 16952 5724 16980
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 7558 16940 7564 16992
rect 7616 16980 7622 16992
rect 8386 16980 8392 16992
rect 7616 16952 8392 16980
rect 7616 16940 7622 16952
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 8846 16940 8852 16992
rect 8904 16980 8910 16992
rect 9309 16983 9367 16989
rect 9309 16980 9321 16983
rect 8904 16952 9321 16980
rect 8904 16940 8910 16952
rect 9309 16949 9321 16952
rect 9355 16949 9367 16983
rect 9309 16943 9367 16949
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 2593 16779 2651 16785
rect 2593 16745 2605 16779
rect 2639 16776 2651 16779
rect 2682 16776 2688 16788
rect 2639 16748 2688 16776
rect 2639 16745 2651 16748
rect 2593 16739 2651 16745
rect 2682 16736 2688 16748
rect 2740 16736 2746 16788
rect 3418 16736 3424 16788
rect 3476 16776 3482 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 3476 16748 3801 16776
rect 3476 16736 3482 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 3789 16739 3847 16745
rect 4798 16736 4804 16788
rect 4856 16776 4862 16788
rect 5169 16779 5227 16785
rect 5169 16776 5181 16779
rect 4856 16748 5181 16776
rect 4856 16736 4862 16748
rect 5169 16745 5181 16748
rect 5215 16776 5227 16779
rect 7285 16779 7343 16785
rect 7285 16776 7297 16779
rect 5215 16748 7297 16776
rect 5215 16745 5227 16748
rect 5169 16739 5227 16745
rect 7285 16745 7297 16748
rect 7331 16745 7343 16779
rect 7285 16739 7343 16745
rect 7374 16736 7380 16788
rect 7432 16776 7438 16788
rect 12391 16779 12449 16785
rect 12391 16776 12403 16779
rect 7432 16748 12403 16776
rect 7432 16736 7438 16748
rect 12391 16745 12403 16748
rect 12437 16745 12449 16779
rect 12391 16739 12449 16745
rect 2035 16711 2093 16717
rect 2035 16677 2047 16711
rect 2081 16708 2093 16711
rect 2130 16708 2136 16720
rect 2081 16680 2136 16708
rect 2081 16677 2093 16680
rect 2035 16671 2093 16677
rect 2130 16668 2136 16680
rect 2188 16668 2194 16720
rect 3878 16668 3884 16720
rect 3936 16708 3942 16720
rect 4246 16708 4252 16720
rect 3936 16680 4252 16708
rect 3936 16668 3942 16680
rect 4246 16668 4252 16680
rect 4304 16668 4310 16720
rect 5534 16708 5540 16720
rect 5495 16680 5540 16708
rect 5534 16668 5540 16680
rect 5592 16668 5598 16720
rect 5718 16668 5724 16720
rect 5776 16708 5782 16720
rect 5813 16711 5871 16717
rect 5813 16708 5825 16711
rect 5776 16680 5825 16708
rect 5776 16668 5782 16680
rect 5813 16677 5825 16680
rect 5859 16677 5871 16711
rect 5813 16671 5871 16677
rect 7466 16668 7472 16720
rect 7524 16708 7530 16720
rect 8297 16711 8355 16717
rect 8297 16708 8309 16711
rect 7524 16680 8309 16708
rect 7524 16668 7530 16680
rect 8297 16677 8309 16680
rect 8343 16708 8355 16711
rect 10962 16708 10968 16720
rect 8343 16680 10968 16708
rect 8343 16677 8355 16680
rect 8297 16671 8355 16677
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 11514 16668 11520 16720
rect 11572 16708 11578 16720
rect 11572 16680 12363 16708
rect 11572 16668 11578 16680
rect 1670 16640 1676 16652
rect 1631 16612 1676 16640
rect 1670 16600 1676 16612
rect 1728 16600 1734 16652
rect 7190 16640 7196 16652
rect 7151 16612 7196 16640
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 7745 16643 7803 16649
rect 7745 16609 7757 16643
rect 7791 16640 7803 16643
rect 8202 16640 8208 16652
rect 7791 16612 8208 16640
rect 7791 16609 7803 16612
rect 7745 16603 7803 16609
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 9674 16640 9680 16652
rect 9635 16612 9680 16640
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 9950 16640 9956 16652
rect 9911 16612 9956 16640
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 11238 16640 11244 16652
rect 11199 16612 11244 16640
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 12335 16649 12363 16680
rect 12320 16643 12378 16649
rect 12320 16609 12332 16643
rect 12366 16640 12378 16643
rect 12618 16640 12624 16652
rect 12366 16612 12624 16640
rect 12366 16609 12378 16612
rect 12320 16603 12378 16609
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 3970 16532 3976 16584
rect 4028 16572 4034 16584
rect 4157 16575 4215 16581
rect 4157 16572 4169 16575
rect 4028 16544 4169 16572
rect 4028 16532 4034 16544
rect 4157 16541 4169 16544
rect 4203 16541 4215 16575
rect 4798 16572 4804 16584
rect 4759 16544 4804 16572
rect 4157 16535 4215 16541
rect 4172 16504 4200 16535
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 5721 16575 5779 16581
rect 5721 16541 5733 16575
rect 5767 16572 5779 16575
rect 5994 16572 6000 16584
rect 5767 16544 6000 16572
rect 5767 16541 5779 16544
rect 5721 16535 5779 16541
rect 5994 16532 6000 16544
rect 6052 16532 6058 16584
rect 6178 16572 6184 16584
rect 6139 16544 6184 16572
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 6730 16532 6736 16584
rect 6788 16572 6794 16584
rect 10137 16575 10195 16581
rect 10137 16572 10149 16575
rect 6788 16544 10149 16572
rect 6788 16532 6794 16544
rect 10137 16541 10149 16544
rect 10183 16541 10195 16575
rect 10137 16535 10195 16541
rect 10870 16532 10876 16584
rect 10928 16572 10934 16584
rect 13170 16572 13176 16584
rect 10928 16544 13176 16572
rect 10928 16532 10934 16544
rect 13170 16532 13176 16544
rect 13228 16532 13234 16584
rect 6196 16504 6224 16532
rect 8662 16504 8668 16516
rect 4172 16476 6224 16504
rect 6840 16476 8668 16504
rect 6840 16448 6868 16476
rect 8662 16464 8668 16476
rect 8720 16504 8726 16516
rect 8849 16507 8907 16513
rect 8849 16504 8861 16507
rect 8720 16476 8861 16504
rect 8720 16464 8726 16476
rect 8849 16473 8861 16476
rect 8895 16473 8907 16507
rect 8849 16467 8907 16473
rect 9306 16464 9312 16516
rect 9364 16504 9370 16516
rect 9769 16507 9827 16513
rect 9769 16504 9781 16507
rect 9364 16476 9781 16504
rect 9364 16464 9370 16476
rect 9769 16473 9781 16476
rect 9815 16473 9827 16507
rect 9769 16467 9827 16473
rect 9858 16464 9864 16516
rect 9916 16504 9922 16516
rect 11425 16507 11483 16513
rect 11425 16504 11437 16507
rect 9916 16476 11437 16504
rect 9916 16464 9922 16476
rect 11425 16473 11437 16476
rect 11471 16473 11483 16507
rect 11425 16467 11483 16473
rect 3050 16436 3056 16448
rect 3011 16408 3056 16436
rect 3050 16396 3056 16408
rect 3108 16396 3114 16448
rect 3142 16396 3148 16448
rect 3200 16436 3206 16448
rect 3329 16439 3387 16445
rect 3329 16436 3341 16439
rect 3200 16408 3341 16436
rect 3200 16396 3206 16408
rect 3329 16405 3341 16408
rect 3375 16405 3387 16439
rect 6822 16436 6828 16448
rect 6783 16408 6828 16436
rect 3329 16399 3387 16405
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 9401 16439 9459 16445
rect 9401 16405 9413 16439
rect 9447 16436 9459 16439
rect 9582 16436 9588 16448
rect 9447 16408 9588 16436
rect 9447 16405 9459 16408
rect 9401 16399 9459 16405
rect 9582 16396 9588 16408
rect 9640 16396 9646 16448
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 2038 16192 2044 16244
rect 2096 16232 2102 16244
rect 2225 16235 2283 16241
rect 2225 16232 2237 16235
rect 2096 16204 2237 16232
rect 2096 16192 2102 16204
rect 2225 16201 2237 16204
rect 2271 16201 2283 16235
rect 4246 16232 4252 16244
rect 4207 16204 4252 16232
rect 2225 16195 2283 16201
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 4709 16235 4767 16241
rect 4709 16201 4721 16235
rect 4755 16232 4767 16235
rect 4982 16232 4988 16244
rect 4755 16204 4988 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 4982 16192 4988 16204
rect 5040 16232 5046 16244
rect 5718 16232 5724 16244
rect 5040 16204 5724 16232
rect 5040 16192 5046 16204
rect 5718 16192 5724 16204
rect 5776 16232 5782 16244
rect 5813 16235 5871 16241
rect 5813 16232 5825 16235
rect 5776 16204 5825 16232
rect 5776 16192 5782 16204
rect 5813 16201 5825 16204
rect 5859 16201 5871 16235
rect 5813 16195 5871 16201
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6273 16235 6331 16241
rect 6273 16232 6285 16235
rect 6052 16204 6285 16232
rect 6052 16192 6058 16204
rect 6273 16201 6285 16204
rect 6319 16232 6331 16235
rect 6638 16232 6644 16244
rect 6319 16204 6644 16232
rect 6319 16201 6331 16204
rect 6273 16195 6331 16201
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 7190 16192 7196 16244
rect 7248 16232 7254 16244
rect 7650 16232 7656 16244
rect 7248 16204 7656 16232
rect 7248 16192 7254 16204
rect 7650 16192 7656 16204
rect 7708 16232 7714 16244
rect 7837 16235 7895 16241
rect 7837 16232 7849 16235
rect 7708 16204 7849 16232
rect 7708 16192 7714 16204
rect 7837 16201 7849 16204
rect 7883 16201 7895 16235
rect 7837 16195 7895 16201
rect 8849 16235 8907 16241
rect 8849 16201 8861 16235
rect 8895 16232 8907 16235
rect 9950 16232 9956 16244
rect 8895 16204 9956 16232
rect 8895 16201 8907 16204
rect 8849 16195 8907 16201
rect 9950 16192 9956 16204
rect 10008 16192 10014 16244
rect 10962 16192 10968 16244
rect 11020 16232 11026 16244
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 11020 16204 11069 16232
rect 11020 16192 11026 16204
rect 11057 16201 11069 16204
rect 11103 16201 11115 16235
rect 12618 16232 12624 16244
rect 12579 16204 12624 16232
rect 11057 16195 11115 16201
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 3234 16124 3240 16176
rect 3292 16164 3298 16176
rect 3292 16136 10916 16164
rect 3292 16124 3298 16136
rect 1302 16056 1308 16108
rect 1360 16096 1366 16108
rect 1535 16099 1593 16105
rect 1535 16096 1547 16099
rect 1360 16068 1547 16096
rect 1360 16056 1366 16068
rect 1535 16065 1547 16068
rect 1581 16065 1593 16099
rect 1535 16059 1593 16065
rect 4890 16056 4896 16108
rect 4948 16096 4954 16108
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 4948 16068 5181 16096
rect 4948 16056 4954 16068
rect 5169 16065 5181 16068
rect 5215 16065 5227 16099
rect 5169 16059 5227 16065
rect 5902 16056 5908 16108
rect 5960 16096 5966 16108
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 5960 16068 7297 16096
rect 5960 16056 5966 16068
rect 7285 16065 7297 16068
rect 7331 16065 7343 16099
rect 9214 16096 9220 16108
rect 9175 16068 9220 16096
rect 7285 16059 7343 16065
rect 9214 16056 9220 16068
rect 9272 16056 9278 16108
rect 9401 16099 9459 16105
rect 9401 16065 9413 16099
rect 9447 16096 9459 16099
rect 9582 16096 9588 16108
rect 9447 16068 9588 16096
rect 9447 16065 9459 16068
rect 9401 16059 9459 16065
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 9674 16056 9680 16108
rect 9732 16096 9738 16108
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 9732 16068 10333 16096
rect 9732 16056 9738 16068
rect 10321 16065 10333 16068
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 1448 16031 1506 16037
rect 1448 15997 1460 16031
rect 1494 16028 1506 16031
rect 2314 16028 2320 16040
rect 1494 16000 2320 16028
rect 1494 15997 1506 16000
rect 1448 15991 1506 15997
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 2961 16031 3019 16037
rect 2961 15997 2973 16031
rect 3007 16028 3019 16031
rect 3050 16028 3056 16040
rect 3007 16000 3056 16028
rect 3007 15997 3019 16000
rect 2961 15991 3019 15997
rect 3050 15988 3056 16000
rect 3108 15988 3114 16040
rect 6822 16028 6828 16040
rect 6783 16000 6828 16028
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 6914 15988 6920 16040
rect 6972 16028 6978 16040
rect 7101 16031 7159 16037
rect 6972 16000 7017 16028
rect 6972 15988 6978 16000
rect 7101 15997 7113 16031
rect 7147 16028 7159 16031
rect 7558 16028 7564 16040
rect 7147 16000 7564 16028
rect 7147 15997 7159 16000
rect 7101 15991 7159 15997
rect 1949 15963 2007 15969
rect 1949 15929 1961 15963
rect 1995 15960 2007 15963
rect 2130 15960 2136 15972
rect 1995 15932 2136 15960
rect 1995 15929 2007 15932
rect 1949 15923 2007 15929
rect 2130 15920 2136 15932
rect 2188 15960 2194 15972
rect 2869 15963 2927 15969
rect 2869 15960 2881 15963
rect 2188 15932 2881 15960
rect 2188 15920 2194 15932
rect 2869 15929 2881 15932
rect 2915 15960 2927 15963
rect 3323 15963 3381 15969
rect 3323 15960 3335 15963
rect 2915 15932 3335 15960
rect 2915 15929 2927 15932
rect 2869 15923 2927 15929
rect 3323 15929 3335 15932
rect 3369 15960 3381 15963
rect 4246 15960 4252 15972
rect 3369 15932 4252 15960
rect 3369 15929 3381 15932
rect 3323 15923 3381 15929
rect 4246 15920 4252 15932
rect 4304 15920 4310 15972
rect 4893 15963 4951 15969
rect 4893 15929 4905 15963
rect 4939 15929 4951 15963
rect 4893 15923 4951 15929
rect 3878 15892 3884 15904
rect 3839 15864 3884 15892
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 4908 15892 4936 15923
rect 4982 15920 4988 15972
rect 5040 15960 5046 15972
rect 6641 15963 6699 15969
rect 5040 15932 5085 15960
rect 5040 15920 5046 15932
rect 6641 15929 6653 15963
rect 6687 15960 6699 15963
rect 7116 15960 7144 15991
rect 7558 15988 7564 16000
rect 7616 15988 7622 16040
rect 10888 16037 10916 16136
rect 10873 16031 10931 16037
rect 10873 15997 10885 16031
rect 10919 16028 10931 16031
rect 11701 16031 11759 16037
rect 11701 16028 11713 16031
rect 10919 16000 11713 16028
rect 10919 15997 10931 16000
rect 10873 15991 10931 15997
rect 11701 15997 11713 16000
rect 11747 15997 11759 16031
rect 11701 15991 11759 15997
rect 6687 15932 7144 15960
rect 6687 15929 6699 15932
rect 6641 15923 6699 15929
rect 9490 15920 9496 15972
rect 9548 15960 9554 15972
rect 10045 15963 10103 15969
rect 9548 15932 9593 15960
rect 9548 15920 9554 15932
rect 10045 15929 10057 15963
rect 10091 15960 10103 15963
rect 10226 15960 10232 15972
rect 10091 15932 10232 15960
rect 10091 15929 10103 15932
rect 10045 15923 10103 15929
rect 10226 15920 10232 15932
rect 10284 15920 10290 15972
rect 10686 15920 10692 15972
rect 10744 15960 10750 15972
rect 11238 15960 11244 15972
rect 10744 15932 11244 15960
rect 10744 15920 10750 15932
rect 11238 15920 11244 15932
rect 11296 15960 11302 15972
rect 11333 15963 11391 15969
rect 11333 15960 11345 15963
rect 11296 15932 11345 15960
rect 11296 15920 11302 15932
rect 11333 15929 11345 15932
rect 11379 15929 11391 15963
rect 11333 15923 11391 15929
rect 5534 15892 5540 15904
rect 4908 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 8202 15892 8208 15904
rect 8163 15864 8208 15892
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 1857 15691 1915 15697
rect 1857 15688 1869 15691
rect 1728 15660 1869 15688
rect 1728 15648 1734 15660
rect 1857 15657 1869 15660
rect 1903 15657 1915 15691
rect 1857 15651 1915 15657
rect 3513 15691 3571 15697
rect 3513 15657 3525 15691
rect 3559 15688 3571 15691
rect 3970 15688 3976 15700
rect 3559 15660 3976 15688
rect 3559 15657 3571 15660
rect 3513 15651 3571 15657
rect 3970 15648 3976 15660
rect 4028 15648 4034 15700
rect 4062 15648 4068 15700
rect 4120 15688 4126 15700
rect 5258 15688 5264 15700
rect 4120 15660 4844 15688
rect 5219 15660 5264 15688
rect 4120 15648 4126 15660
rect 4816 15632 4844 15660
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 9582 15648 9588 15700
rect 9640 15688 9646 15700
rect 12943 15691 13001 15697
rect 12943 15688 12955 15691
rect 9640 15660 12955 15688
rect 9640 15648 9646 15660
rect 12943 15657 12955 15660
rect 12989 15657 13001 15691
rect 12943 15651 13001 15657
rect 1397 15623 1455 15629
rect 1397 15589 1409 15623
rect 1443 15620 1455 15623
rect 2038 15620 2044 15632
rect 1443 15592 2044 15620
rect 1443 15589 1455 15592
rect 1397 15583 1455 15589
rect 2038 15580 2044 15592
rect 2096 15580 2102 15632
rect 3142 15620 3148 15632
rect 3103 15592 3148 15620
rect 3142 15580 3148 15592
rect 3200 15580 3206 15632
rect 3878 15580 3884 15632
rect 3936 15620 3942 15632
rect 4249 15623 4307 15629
rect 4249 15620 4261 15623
rect 3936 15592 4261 15620
rect 3936 15580 3942 15592
rect 4249 15589 4261 15592
rect 4295 15620 4307 15623
rect 4614 15620 4620 15632
rect 4295 15592 4620 15620
rect 4295 15589 4307 15592
rect 4249 15583 4307 15589
rect 4614 15580 4620 15592
rect 4672 15580 4678 15632
rect 4798 15620 4804 15632
rect 4759 15592 4804 15620
rect 4798 15580 4804 15592
rect 4856 15580 4862 15632
rect 9214 15620 9220 15632
rect 6380 15592 9220 15620
rect 2406 15552 2412 15564
rect 2367 15524 2412 15552
rect 2406 15512 2412 15524
rect 2464 15512 2470 15564
rect 2958 15552 2964 15564
rect 2919 15524 2964 15552
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 6270 15512 6276 15564
rect 6328 15552 6334 15564
rect 6380 15561 6408 15592
rect 9214 15580 9220 15592
rect 9272 15580 9278 15632
rect 9401 15623 9459 15629
rect 9401 15589 9413 15623
rect 9447 15620 9459 15623
rect 9490 15620 9496 15632
rect 9447 15592 9496 15620
rect 9447 15589 9459 15592
rect 9401 15583 9459 15589
rect 9490 15580 9496 15592
rect 9548 15620 9554 15632
rect 9858 15620 9864 15632
rect 9548 15592 9864 15620
rect 9548 15580 9554 15592
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 11241 15623 11299 15629
rect 11241 15620 11253 15623
rect 10008 15592 11253 15620
rect 10008 15580 10014 15592
rect 11241 15589 11253 15592
rect 11287 15589 11299 15623
rect 11241 15583 11299 15589
rect 6365 15555 6423 15561
rect 6365 15552 6377 15555
rect 6328 15524 6377 15552
rect 6328 15512 6334 15524
rect 6365 15521 6377 15524
rect 6411 15521 6423 15555
rect 6365 15515 6423 15521
rect 7285 15555 7343 15561
rect 7285 15521 7297 15555
rect 7331 15552 7343 15555
rect 7331 15524 7512 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 3881 15487 3939 15493
rect 3881 15453 3893 15487
rect 3927 15484 3939 15487
rect 4157 15487 4215 15493
rect 4157 15484 4169 15487
rect 3927 15456 4169 15484
rect 3927 15453 3939 15456
rect 3881 15447 3939 15453
rect 4157 15453 4169 15456
rect 4203 15484 4215 15487
rect 4890 15484 4896 15496
rect 4203 15456 4896 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15453 6515 15487
rect 6457 15447 6515 15453
rect 2314 15416 2320 15428
rect 2227 15388 2320 15416
rect 2314 15376 2320 15388
rect 2372 15416 2378 15428
rect 4062 15416 4068 15428
rect 2372 15388 4068 15416
rect 2372 15376 2378 15388
rect 4062 15376 4068 15388
rect 4120 15376 4126 15428
rect 6472 15416 6500 15447
rect 7484 15428 7512 15524
rect 7558 15512 7564 15564
rect 7616 15552 7622 15564
rect 11422 15552 11428 15564
rect 7616 15524 7661 15552
rect 11383 15524 11428 15552
rect 7616 15512 7622 15524
rect 11422 15512 11428 15524
rect 11480 15512 11486 15564
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 12872 15555 12930 15561
rect 12872 15552 12884 15555
rect 12492 15524 12884 15552
rect 12492 15512 12498 15524
rect 12872 15521 12884 15524
rect 12918 15552 12930 15555
rect 13446 15552 13452 15564
rect 12918 15524 13452 15552
rect 12918 15521 12930 15524
rect 12872 15515 12930 15521
rect 13446 15512 13452 15524
rect 13504 15512 13510 15564
rect 7742 15484 7748 15496
rect 7703 15456 7748 15484
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 9769 15487 9827 15493
rect 9769 15453 9781 15487
rect 9815 15484 9827 15487
rect 9950 15484 9956 15496
rect 9815 15456 9956 15484
rect 9815 15453 9827 15456
rect 9769 15447 9827 15453
rect 9950 15444 9956 15456
rect 10008 15444 10014 15496
rect 10410 15484 10416 15496
rect 10371 15456 10416 15484
rect 10410 15444 10416 15456
rect 10468 15444 10474 15496
rect 6914 15416 6920 15428
rect 6472 15388 6920 15416
rect 6914 15376 6920 15388
rect 6972 15416 6978 15428
rect 7374 15416 7380 15428
rect 6972 15388 7380 15416
rect 6972 15376 6978 15388
rect 7374 15376 7380 15388
rect 7432 15376 7438 15428
rect 7466 15376 7472 15428
rect 7524 15416 7530 15428
rect 8110 15416 8116 15428
rect 7524 15388 8116 15416
rect 7524 15376 7530 15388
rect 8110 15376 8116 15388
rect 8168 15416 8174 15428
rect 9674 15416 9680 15428
rect 8168 15388 9680 15416
rect 8168 15376 8174 15388
rect 9674 15376 9680 15388
rect 9732 15376 9738 15428
rect 8294 15348 8300 15360
rect 8255 15320 8300 15348
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 8754 15348 8760 15360
rect 8667 15320 8760 15348
rect 8754 15308 8760 15320
rect 8812 15348 8818 15360
rect 11330 15348 11336 15360
rect 8812 15320 11336 15348
rect 8812 15308 8818 15320
rect 11330 15308 11336 15320
rect 11388 15308 11394 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 1673 15147 1731 15153
rect 1673 15113 1685 15147
rect 1719 15144 1731 15147
rect 1946 15144 1952 15156
rect 1719 15116 1952 15144
rect 1719 15113 1731 15116
rect 1673 15107 1731 15113
rect 1946 15104 1952 15116
rect 2004 15144 2010 15156
rect 2958 15144 2964 15156
rect 2004 15116 2964 15144
rect 2004 15104 2010 15116
rect 2958 15104 2964 15116
rect 3016 15104 3022 15156
rect 4433 15147 4491 15153
rect 4433 15113 4445 15147
rect 4479 15144 4491 15147
rect 4709 15147 4767 15153
rect 4709 15144 4721 15147
rect 4479 15116 4721 15144
rect 4479 15113 4491 15116
rect 4433 15107 4491 15113
rect 4709 15113 4721 15116
rect 4755 15144 4767 15147
rect 6730 15144 6736 15156
rect 4755 15116 6736 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 7377 15147 7435 15153
rect 7377 15113 7389 15147
rect 7423 15144 7435 15147
rect 7466 15144 7472 15156
rect 7423 15116 7472 15144
rect 7423 15113 7435 15116
rect 7377 15107 7435 15113
rect 7466 15104 7472 15116
rect 7524 15104 7530 15156
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 7745 15147 7803 15153
rect 7745 15144 7757 15147
rect 7616 15116 7757 15144
rect 7616 15104 7622 15116
rect 7745 15113 7757 15116
rect 7791 15144 7803 15147
rect 9309 15147 9367 15153
rect 7791 15116 8340 15144
rect 7791 15113 7803 15116
rect 7745 15107 7803 15113
rect 1578 15036 1584 15088
rect 1636 15076 1642 15088
rect 2041 15079 2099 15085
rect 2041 15076 2053 15079
rect 1636 15048 2053 15076
rect 1636 15036 1642 15048
rect 2041 15045 2053 15048
rect 2087 15045 2099 15079
rect 2406 15076 2412 15088
rect 2367 15048 2412 15076
rect 2041 15039 2099 15045
rect 1489 14943 1547 14949
rect 1489 14909 1501 14943
rect 1535 14940 1547 14943
rect 1578 14940 1584 14952
rect 1535 14912 1584 14940
rect 1535 14909 1547 14912
rect 1489 14903 1547 14909
rect 1578 14900 1584 14912
rect 1636 14900 1642 14952
rect 2056 14940 2084 15039
rect 2406 15036 2412 15048
rect 2464 15036 2470 15088
rect 3605 15079 3663 15085
rect 3605 15045 3617 15079
rect 3651 15076 3663 15079
rect 3973 15079 4031 15085
rect 3973 15076 3985 15079
rect 3651 15048 3985 15076
rect 3651 15045 3663 15048
rect 3605 15039 3663 15045
rect 3973 15045 3985 15048
rect 4019 15076 4031 15079
rect 8202 15076 8208 15088
rect 4019 15048 8208 15076
rect 4019 15045 4031 15048
rect 3973 15039 4031 15045
rect 3050 15008 3056 15020
rect 3011 14980 3056 15008
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 2501 14943 2559 14949
rect 2501 14940 2513 14943
rect 2056 14912 2513 14940
rect 2501 14909 2513 14912
rect 2547 14940 2559 14943
rect 2774 14940 2780 14952
rect 2547 14912 2780 14940
rect 2547 14909 2559 14912
rect 2501 14903 2559 14909
rect 2774 14900 2780 14912
rect 2832 14900 2838 14952
rect 2958 14940 2964 14952
rect 2871 14912 2964 14940
rect 2958 14900 2964 14912
rect 3016 14940 3022 14952
rect 3620 14940 3648 15039
rect 8202 15036 8208 15048
rect 8260 15036 8266 15088
rect 8312 15076 8340 15116
rect 9309 15113 9321 15147
rect 9355 15144 9367 15147
rect 9858 15144 9864 15156
rect 9355 15116 9864 15144
rect 9355 15113 9367 15116
rect 9309 15107 9367 15113
rect 9858 15104 9864 15116
rect 9916 15144 9922 15156
rect 10689 15147 10747 15153
rect 10689 15144 10701 15147
rect 9916 15116 10701 15144
rect 9916 15104 9922 15116
rect 10689 15113 10701 15116
rect 10735 15113 10747 15147
rect 10689 15107 10747 15113
rect 11333 15147 11391 15153
rect 11333 15113 11345 15147
rect 11379 15144 11391 15147
rect 11422 15144 11428 15156
rect 11379 15116 11428 15144
rect 11379 15113 11391 15116
rect 11333 15107 11391 15113
rect 11348 15076 11376 15107
rect 11422 15104 11428 15116
rect 11480 15104 11486 15156
rect 8312 15048 11376 15076
rect 6270 15008 6276 15020
rect 6231 14980 6276 15008
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 15008 8079 15011
rect 8754 15008 8760 15020
rect 8067 14980 8760 15008
rect 8067 14977 8079 14980
rect 8021 14971 8079 14977
rect 8754 14968 8760 14980
rect 8812 14968 8818 15020
rect 3016 14912 3648 14940
rect 4157 14943 4215 14949
rect 3016 14900 3022 14912
rect 4157 14909 4169 14943
rect 4203 14940 4215 14943
rect 4433 14943 4491 14949
rect 4433 14940 4445 14943
rect 4203 14912 4445 14940
rect 4203 14909 4215 14912
rect 4157 14903 4215 14909
rect 4433 14909 4445 14912
rect 4479 14909 4491 14943
rect 4433 14903 4491 14909
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14940 5135 14943
rect 5169 14943 5227 14949
rect 5169 14940 5181 14943
rect 5123 14912 5181 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 5169 14909 5181 14912
rect 5215 14909 5227 14943
rect 5169 14903 5227 14909
rect 5184 14872 5212 14903
rect 5258 14900 5264 14952
rect 5316 14940 5322 14952
rect 5718 14940 5724 14952
rect 5316 14912 5724 14940
rect 5316 14900 5322 14912
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 5902 14940 5908 14952
rect 5863 14912 5908 14940
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14940 6699 14943
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6687 14912 6837 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 6825 14909 6837 14912
rect 6871 14940 6883 14943
rect 7742 14940 7748 14952
rect 6871 14912 7748 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 7742 14900 7748 14912
rect 7800 14900 7806 14952
rect 9766 14940 9772 14952
rect 9727 14912 9772 14940
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 11514 14900 11520 14952
rect 11572 14940 11578 14952
rect 12253 14943 12311 14949
rect 12253 14940 12265 14943
rect 11572 14912 12265 14940
rect 11572 14900 11578 14912
rect 12253 14909 12265 14912
rect 12299 14940 12311 14943
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12299 14912 12449 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 12710 14900 12716 14952
rect 12768 14940 12774 14952
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12768 14912 12909 14940
rect 12768 14900 12774 14912
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 7926 14872 7932 14884
rect 5184 14844 7932 14872
rect 7926 14832 7932 14844
rect 7984 14832 7990 14884
rect 9585 14875 9643 14881
rect 9585 14872 9597 14875
rect 8404 14844 9597 14872
rect 4341 14807 4399 14813
rect 4341 14773 4353 14807
rect 4387 14804 4399 14807
rect 4430 14804 4436 14816
rect 4387 14776 4436 14804
rect 4387 14773 4399 14776
rect 4341 14767 4399 14773
rect 4430 14764 4436 14776
rect 4488 14764 4494 14816
rect 5718 14764 5724 14816
rect 5776 14804 5782 14816
rect 7009 14807 7067 14813
rect 7009 14804 7021 14807
rect 5776 14776 7021 14804
rect 5776 14764 5782 14776
rect 7009 14773 7021 14776
rect 7055 14773 7067 14807
rect 7009 14767 7067 14773
rect 8294 14764 8300 14816
rect 8352 14804 8358 14816
rect 8404 14813 8432 14844
rect 9585 14841 9597 14844
rect 9631 14872 9643 14875
rect 10090 14875 10148 14881
rect 10090 14872 10102 14875
rect 9631 14844 10102 14872
rect 9631 14841 9643 14844
rect 9585 14835 9643 14841
rect 10090 14841 10102 14844
rect 10136 14841 10148 14875
rect 10090 14835 10148 14841
rect 8389 14807 8447 14813
rect 8389 14804 8401 14807
rect 8352 14776 8401 14804
rect 8352 14764 8358 14776
rect 8389 14773 8401 14776
rect 8435 14773 8447 14807
rect 8938 14804 8944 14816
rect 8899 14776 8944 14804
rect 8389 14767 8447 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 11330 14764 11336 14816
rect 11388 14804 11394 14816
rect 12529 14807 12587 14813
rect 12529 14804 12541 14807
rect 11388 14776 12541 14804
rect 11388 14764 11394 14776
rect 12529 14773 12541 14776
rect 12575 14773 12587 14807
rect 13446 14804 13452 14816
rect 13407 14776 13452 14804
rect 12529 14767 12587 14773
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 4614 14600 4620 14612
rect 4575 14572 4620 14600
rect 4614 14560 4620 14572
rect 4672 14560 4678 14612
rect 7374 14600 7380 14612
rect 7335 14572 7380 14600
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 9493 14603 9551 14609
rect 9493 14569 9505 14603
rect 9539 14600 9551 14603
rect 9766 14600 9772 14612
rect 9539 14572 9772 14600
rect 9539 14569 9551 14572
rect 9493 14563 9551 14569
rect 9766 14560 9772 14572
rect 9824 14600 9830 14612
rect 11333 14603 11391 14609
rect 11333 14600 11345 14603
rect 9824 14572 11345 14600
rect 9824 14560 9830 14572
rect 11333 14569 11345 14572
rect 11379 14569 11391 14603
rect 11333 14563 11391 14569
rect 1535 14535 1593 14541
rect 1535 14501 1547 14535
rect 1581 14532 1593 14535
rect 3789 14535 3847 14541
rect 3789 14532 3801 14535
rect 1581 14504 3801 14532
rect 1581 14501 1593 14504
rect 1535 14495 1593 14501
rect 3789 14501 3801 14504
rect 3835 14532 3847 14535
rect 4338 14532 4344 14544
rect 3835 14504 4344 14532
rect 3835 14501 3847 14504
rect 3789 14495 3847 14501
rect 4338 14492 4344 14504
rect 4396 14492 4402 14544
rect 4982 14532 4988 14544
rect 4943 14504 4988 14532
rect 4982 14492 4988 14504
rect 5040 14492 5046 14544
rect 6178 14492 6184 14544
rect 6236 14532 6242 14544
rect 7006 14532 7012 14544
rect 6236 14504 7012 14532
rect 6236 14492 6242 14504
rect 1448 14467 1506 14473
rect 1448 14433 1460 14467
rect 1494 14464 1506 14467
rect 1762 14464 1768 14476
rect 1494 14436 1768 14464
rect 1494 14433 1506 14436
rect 1448 14427 1506 14433
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 2406 14464 2412 14476
rect 2367 14436 2412 14464
rect 2406 14424 2412 14436
rect 2464 14424 2470 14476
rect 2682 14464 2688 14476
rect 2643 14436 2688 14464
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14464 3203 14467
rect 3234 14464 3240 14476
rect 3191 14436 3240 14464
rect 3191 14433 3203 14436
rect 3145 14427 3203 14433
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 6362 14464 6368 14476
rect 6323 14436 6368 14464
rect 6362 14424 6368 14436
rect 6420 14424 6426 14476
rect 6472 14473 6500 14504
rect 7006 14492 7012 14504
rect 7064 14492 7070 14544
rect 8662 14532 8668 14544
rect 8496 14504 8668 14532
rect 6457 14467 6515 14473
rect 6457 14433 6469 14467
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 6546 14424 6552 14476
rect 6604 14464 6610 14476
rect 6641 14467 6699 14473
rect 6641 14464 6653 14467
rect 6604 14436 6653 14464
rect 6604 14424 6610 14436
rect 6641 14433 6653 14436
rect 6687 14464 6699 14467
rect 7558 14464 7564 14476
rect 6687 14436 7564 14464
rect 6687 14433 6699 14436
rect 6641 14427 6699 14433
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 7926 14464 7932 14476
rect 7887 14436 7932 14464
rect 7926 14424 7932 14436
rect 7984 14424 7990 14476
rect 8496 14473 8524 14504
rect 8662 14492 8668 14504
rect 8720 14492 8726 14544
rect 8938 14492 8944 14544
rect 8996 14532 9002 14544
rect 9582 14532 9588 14544
rect 8996 14504 9588 14532
rect 8996 14492 9002 14504
rect 9582 14492 9588 14504
rect 9640 14532 9646 14544
rect 9861 14535 9919 14541
rect 9861 14532 9873 14535
rect 9640 14504 9873 14532
rect 9640 14492 9646 14504
rect 9861 14501 9873 14504
rect 9907 14501 9919 14535
rect 10410 14532 10416 14544
rect 10371 14504 10416 14532
rect 9861 14495 9919 14501
rect 10410 14492 10416 14504
rect 10468 14492 10474 14544
rect 10962 14492 10968 14544
rect 11020 14532 11026 14544
rect 12437 14535 12495 14541
rect 12437 14532 12449 14535
rect 11020 14504 12449 14532
rect 11020 14492 11026 14504
rect 12437 14501 12449 14504
rect 12483 14532 12495 14535
rect 12710 14532 12716 14544
rect 12483 14504 12716 14532
rect 12483 14501 12495 14504
rect 12437 14495 12495 14501
rect 12710 14492 12716 14504
rect 12768 14492 12774 14544
rect 8481 14467 8539 14473
rect 8481 14464 8493 14467
rect 8404 14436 8493 14464
rect 8404 14408 8432 14436
rect 8481 14433 8493 14436
rect 8527 14433 8539 14467
rect 11514 14464 11520 14476
rect 11475 14436 11520 14464
rect 8481 14427 8539 14433
rect 11514 14424 11520 14436
rect 11572 14424 11578 14476
rect 11698 14464 11704 14476
rect 11659 14436 11704 14464
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 12856 14467 12914 14473
rect 12856 14433 12868 14467
rect 12902 14464 12914 14467
rect 13262 14464 13268 14476
rect 12902 14436 13268 14464
rect 12902 14433 12914 14436
rect 12856 14427 12914 14433
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 1578 14356 1584 14408
rect 1636 14396 1642 14408
rect 1949 14399 2007 14405
rect 1949 14396 1961 14399
rect 1636 14368 1961 14396
rect 1636 14356 1642 14368
rect 1949 14365 1961 14368
rect 1995 14396 2007 14399
rect 4706 14396 4712 14408
rect 1995 14368 4712 14396
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 4706 14356 4712 14368
rect 4764 14356 4770 14408
rect 4890 14396 4896 14408
rect 4851 14368 4896 14396
rect 4890 14356 4896 14368
rect 4948 14356 4954 14408
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 5000 14368 6837 14396
rect 2501 14331 2559 14337
rect 2501 14297 2513 14331
rect 2547 14328 2559 14331
rect 3142 14328 3148 14340
rect 2547 14300 3148 14328
rect 2547 14297 2559 14300
rect 2501 14291 2559 14297
rect 3142 14288 3148 14300
rect 3200 14288 3206 14340
rect 5000 14328 5028 14368
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 8386 14356 8392 14408
rect 8444 14356 8450 14408
rect 8662 14396 8668 14408
rect 8623 14368 8668 14396
rect 8662 14356 8668 14368
rect 8720 14356 8726 14408
rect 9769 14399 9827 14405
rect 9769 14396 9781 14399
rect 9692 14368 9781 14396
rect 9692 14340 9720 14368
rect 9769 14365 9781 14368
rect 9815 14396 9827 14399
rect 12943 14399 13001 14405
rect 12943 14396 12955 14399
rect 9815 14368 12955 14396
rect 9815 14365 9827 14368
rect 9769 14359 9827 14365
rect 12943 14365 12955 14368
rect 12989 14365 13001 14399
rect 12943 14359 13001 14365
rect 3252 14300 5028 14328
rect 5445 14331 5503 14337
rect 2314 14260 2320 14272
rect 2227 14232 2320 14260
rect 2314 14220 2320 14232
rect 2372 14260 2378 14272
rect 3252 14260 3280 14300
rect 5445 14297 5457 14331
rect 5491 14328 5503 14331
rect 6178 14328 6184 14340
rect 5491 14300 6184 14328
rect 5491 14297 5503 14300
rect 5445 14291 5503 14297
rect 6178 14288 6184 14300
rect 6236 14288 6242 14340
rect 7558 14288 7564 14340
rect 7616 14328 7622 14340
rect 8570 14328 8576 14340
rect 7616 14300 8576 14328
rect 7616 14288 7622 14300
rect 8570 14288 8576 14300
rect 8628 14288 8634 14340
rect 9674 14288 9680 14340
rect 9732 14288 9738 14340
rect 3418 14260 3424 14272
rect 2372 14232 3280 14260
rect 3379 14232 3424 14260
rect 2372 14220 2378 14232
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 4341 14263 4399 14269
rect 4341 14229 4353 14263
rect 4387 14260 4399 14263
rect 4430 14260 4436 14272
rect 4387 14232 4436 14260
rect 4387 14229 4399 14232
rect 4341 14223 4399 14229
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 6822 14220 6828 14272
rect 6880 14260 6886 14272
rect 8478 14260 8484 14272
rect 6880 14232 8484 14260
rect 6880 14220 6886 14232
rect 8478 14220 8484 14232
rect 8536 14220 8542 14272
rect 9125 14263 9183 14269
rect 9125 14229 9137 14263
rect 9171 14260 9183 14263
rect 9950 14260 9956 14272
rect 9171 14232 9956 14260
rect 9171 14229 9183 14232
rect 9125 14223 9183 14229
rect 9950 14220 9956 14232
rect 10008 14260 10014 14272
rect 11606 14260 11612 14272
rect 10008 14232 11612 14260
rect 10008 14220 10014 14232
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 2682 14056 2688 14068
rect 2547 14028 2688 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 2682 14016 2688 14028
rect 2740 14056 2746 14068
rect 4798 14056 4804 14068
rect 2740 14028 4804 14056
rect 2740 14016 2746 14028
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 4982 14016 4988 14068
rect 5040 14056 5046 14068
rect 5261 14059 5319 14065
rect 5261 14056 5273 14059
rect 5040 14028 5273 14056
rect 5040 14016 5046 14028
rect 5261 14025 5273 14028
rect 5307 14025 5319 14059
rect 5261 14019 5319 14025
rect 5445 14059 5503 14065
rect 5445 14025 5457 14059
rect 5491 14056 5503 14059
rect 5721 14059 5779 14065
rect 5721 14056 5733 14059
rect 5491 14028 5733 14056
rect 5491 14025 5503 14028
rect 5445 14019 5503 14025
rect 5721 14025 5733 14028
rect 5767 14056 5779 14059
rect 6086 14056 6092 14068
rect 5767 14028 6092 14056
rect 5767 14025 5779 14028
rect 5721 14019 5779 14025
rect 6086 14016 6092 14028
rect 6144 14016 6150 14068
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 6457 14059 6515 14065
rect 6457 14056 6469 14059
rect 6420 14028 6469 14056
rect 6420 14016 6426 14028
rect 6457 14025 6469 14028
rect 6503 14056 6515 14059
rect 7466 14056 7472 14068
rect 6503 14028 7472 14056
rect 6503 14025 6515 14028
rect 6457 14019 6515 14025
rect 7466 14016 7472 14028
rect 7524 14016 7530 14068
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 7800 14028 7849 14056
rect 7800 14016 7806 14028
rect 7837 14025 7849 14028
rect 7883 14056 7895 14059
rect 7926 14056 7932 14068
rect 7883 14028 7932 14056
rect 7883 14025 7895 14028
rect 7837 14019 7895 14025
rect 7926 14016 7932 14028
rect 7984 14016 7990 14068
rect 9582 14056 9588 14068
rect 9543 14028 9588 14056
rect 9582 14016 9588 14028
rect 9640 14056 9646 14068
rect 9858 14056 9864 14068
rect 9640 14028 9864 14056
rect 9640 14016 9646 14028
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 11146 14016 11152 14068
rect 11204 14056 11210 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 11204 14028 11345 14056
rect 11204 14016 11210 14028
rect 11333 14025 11345 14028
rect 11379 14056 11391 14059
rect 11514 14056 11520 14068
rect 11379 14028 11520 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11514 14016 11520 14028
rect 11572 14016 11578 14068
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 12575 14059 12633 14065
rect 12575 14056 12587 14059
rect 11664 14028 12587 14056
rect 11664 14016 11670 14028
rect 12575 14025 12587 14028
rect 12621 14025 12633 14059
rect 13262 14056 13268 14068
rect 13223 14028 13268 14056
rect 12575 14019 12633 14025
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 2406 13948 2412 14000
rect 2464 13988 2470 14000
rect 4157 13991 4215 13997
rect 4157 13988 4169 13991
rect 2464 13960 4169 13988
rect 2464 13948 2470 13960
rect 4157 13957 4169 13960
rect 4203 13988 4215 13991
rect 6822 13988 6828 14000
rect 4203 13960 6828 13988
rect 4203 13957 4215 13960
rect 4157 13951 4215 13957
rect 6822 13948 6828 13960
rect 6880 13948 6886 14000
rect 6914 13948 6920 14000
rect 6972 13988 6978 14000
rect 7009 13991 7067 13997
rect 7009 13988 7021 13991
rect 6972 13960 7021 13988
rect 6972 13948 6978 13960
rect 7009 13957 7021 13960
rect 7055 13957 7067 13991
rect 7009 13951 7067 13957
rect 7101 13991 7159 13997
rect 7101 13957 7113 13991
rect 7147 13988 7159 13991
rect 7377 13991 7435 13997
rect 7377 13988 7389 13991
rect 7147 13960 7389 13988
rect 7147 13957 7159 13960
rect 7101 13951 7159 13957
rect 7377 13957 7389 13960
rect 7423 13988 7435 13991
rect 8846 13988 8852 14000
rect 7423 13960 8852 13988
rect 7423 13957 7435 13960
rect 7377 13951 7435 13957
rect 8846 13948 8852 13960
rect 8904 13948 8910 14000
rect 9217 13991 9275 13997
rect 9217 13957 9229 13991
rect 9263 13988 9275 13991
rect 13280 13988 13308 14016
rect 9263 13960 9628 13988
rect 9263 13957 9275 13960
rect 9217 13951 9275 13957
rect 2222 13880 2228 13932
rect 2280 13920 2286 13932
rect 2280 13892 2452 13920
rect 2280 13880 2286 13892
rect 2424 13864 2452 13892
rect 2498 13880 2504 13932
rect 2556 13920 2562 13932
rect 4338 13920 4344 13932
rect 2556 13892 2728 13920
rect 4299 13892 4344 13920
rect 2556 13880 2562 13892
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 2314 13852 2320 13864
rect 1719 13824 2320 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 2314 13812 2320 13824
rect 2372 13812 2378 13864
rect 2406 13812 2412 13864
rect 2464 13812 2470 13864
rect 2700 13861 2728 13892
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 4798 13880 4804 13932
rect 4856 13920 4862 13932
rect 4856 13892 5580 13920
rect 4856 13880 4862 13892
rect 5552 13864 5580 13892
rect 5902 13880 5908 13932
rect 5960 13920 5966 13932
rect 8297 13923 8355 13929
rect 8297 13920 8309 13923
rect 5960 13892 8309 13920
rect 5960 13880 5966 13892
rect 8297 13889 8309 13892
rect 8343 13920 8355 13923
rect 8754 13920 8760 13932
rect 8343 13892 8760 13920
rect 8343 13889 8355 13892
rect 8297 13883 8355 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 2685 13855 2743 13861
rect 2685 13821 2697 13855
rect 2731 13852 2743 13855
rect 3050 13852 3056 13864
rect 2731 13824 3056 13852
rect 2731 13821 2743 13824
rect 2685 13815 2743 13821
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 3237 13855 3295 13861
rect 3237 13852 3249 13855
rect 3160 13824 3249 13852
rect 2866 13744 2872 13796
rect 2924 13784 2930 13796
rect 3160 13784 3188 13824
rect 3237 13821 3249 13824
rect 3283 13852 3295 13855
rect 3418 13852 3424 13864
rect 3283 13824 3424 13852
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 5534 13812 5540 13864
rect 5592 13852 5598 13864
rect 5997 13855 6055 13861
rect 5997 13852 6009 13855
rect 5592 13824 6009 13852
rect 5592 13812 5598 13824
rect 5997 13821 6009 13824
rect 6043 13852 6055 13855
rect 6546 13852 6552 13864
rect 6043 13824 6552 13852
rect 6043 13821 6055 13824
rect 5997 13815 6055 13821
rect 6546 13812 6552 13824
rect 6604 13812 6610 13864
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13852 6883 13855
rect 7101 13855 7159 13861
rect 7101 13852 7113 13855
rect 6871 13824 7113 13852
rect 6871 13821 6883 13824
rect 6825 13815 6883 13821
rect 7101 13821 7113 13824
rect 7147 13821 7159 13855
rect 7101 13815 7159 13821
rect 4430 13784 4436 13796
rect 2924 13756 3188 13784
rect 4391 13756 4436 13784
rect 2924 13744 2930 13756
rect 4430 13744 4436 13756
rect 4488 13744 4494 13796
rect 4985 13787 5043 13793
rect 4985 13753 4997 13787
rect 5031 13784 5043 13787
rect 5626 13784 5632 13796
rect 5031 13756 5632 13784
rect 5031 13753 5043 13756
rect 4985 13747 5043 13753
rect 5626 13744 5632 13756
rect 5684 13784 5690 13796
rect 6086 13784 6092 13796
rect 5684 13756 6092 13784
rect 5684 13744 5690 13756
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 7926 13744 7932 13796
rect 7984 13784 7990 13796
rect 8113 13787 8171 13793
rect 8113 13784 8125 13787
rect 7984 13756 8125 13784
rect 7984 13744 7990 13756
rect 8113 13753 8125 13756
rect 8159 13784 8171 13787
rect 8294 13784 8300 13796
rect 8159 13756 8300 13784
rect 8159 13753 8171 13756
rect 8113 13747 8171 13753
rect 8294 13744 8300 13756
rect 8352 13784 8358 13796
rect 8618 13787 8676 13793
rect 8618 13784 8630 13787
rect 8352 13756 8630 13784
rect 8352 13744 8358 13756
rect 8618 13753 8630 13756
rect 8664 13753 8676 13787
rect 9600 13784 9628 13960
rect 11348 13960 13308 13988
rect 11348 13932 11376 13960
rect 10226 13880 10232 13932
rect 10284 13920 10290 13932
rect 10410 13920 10416 13932
rect 10284 13892 10416 13920
rect 10284 13880 10290 13892
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 11330 13880 11336 13932
rect 11388 13880 11394 13932
rect 11698 13920 11704 13932
rect 11659 13892 11704 13920
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 12894 13920 12900 13932
rect 12503 13892 12900 13920
rect 12503 13861 12531 13892
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 12488 13855 12546 13861
rect 12488 13821 12500 13855
rect 12534 13821 12546 13855
rect 12488 13815 12546 13821
rect 13516 13855 13574 13861
rect 13516 13821 13528 13855
rect 13562 13852 13574 13855
rect 13562 13821 13584 13852
rect 13516 13815 13584 13821
rect 9950 13784 9956 13796
rect 9600 13756 9956 13784
rect 8618 13747 8676 13753
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 10134 13784 10140 13796
rect 10095 13756 10140 13784
rect 10134 13744 10140 13756
rect 10192 13744 10198 13796
rect 10229 13787 10287 13793
rect 10229 13753 10241 13787
rect 10275 13753 10287 13787
rect 10229 13747 10287 13753
rect 1854 13716 1860 13728
rect 1815 13688 1860 13716
rect 1854 13676 1860 13688
rect 1912 13676 1918 13728
rect 2958 13716 2964 13728
rect 2919 13688 2964 13716
rect 2958 13676 2964 13688
rect 3016 13676 3022 13728
rect 3142 13676 3148 13728
rect 3200 13716 3206 13728
rect 3697 13719 3755 13725
rect 3697 13716 3709 13719
rect 3200 13688 3709 13716
rect 3200 13676 3206 13688
rect 3697 13685 3709 13688
rect 3743 13716 3755 13719
rect 5445 13719 5503 13725
rect 5445 13716 5457 13719
rect 3743 13688 5457 13716
rect 3743 13685 3755 13688
rect 3697 13679 3755 13685
rect 5445 13685 5457 13688
rect 5491 13685 5503 13719
rect 5445 13679 5503 13685
rect 5994 13676 6000 13728
rect 6052 13716 6058 13728
rect 8018 13716 8024 13728
rect 6052 13688 8024 13716
rect 6052 13676 6058 13688
rect 8018 13676 8024 13688
rect 8076 13676 8082 13728
rect 9858 13676 9864 13728
rect 9916 13716 9922 13728
rect 10244 13716 10272 13747
rect 13078 13744 13084 13796
rect 13136 13784 13142 13796
rect 13556 13784 13584 13815
rect 13909 13787 13967 13793
rect 13909 13784 13921 13787
rect 13136 13756 13921 13784
rect 13136 13744 13142 13756
rect 13909 13753 13921 13756
rect 13955 13753 13967 13787
rect 13909 13747 13967 13753
rect 9916 13688 10272 13716
rect 9916 13676 9922 13688
rect 10594 13676 10600 13728
rect 10652 13716 10658 13728
rect 11330 13716 11336 13728
rect 10652 13688 11336 13716
rect 10652 13676 10658 13688
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 12894 13716 12900 13728
rect 12855 13688 12900 13716
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 12986 13676 12992 13728
rect 13044 13716 13050 13728
rect 13587 13719 13645 13725
rect 13587 13716 13599 13719
rect 13044 13688 13599 13716
rect 13044 13676 13050 13688
rect 13587 13685 13599 13688
rect 13633 13685 13645 13719
rect 13587 13679 13645 13685
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 1854 13472 1860 13524
rect 1912 13512 1918 13524
rect 3605 13515 3663 13521
rect 3605 13512 3617 13515
rect 1912 13484 3617 13512
rect 1912 13472 1918 13484
rect 3605 13481 3617 13484
rect 3651 13481 3663 13515
rect 3605 13475 3663 13481
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4433 13515 4491 13521
rect 4433 13512 4445 13515
rect 4396 13484 4445 13512
rect 4396 13472 4402 13484
rect 4433 13481 4445 13484
rect 4479 13481 4491 13515
rect 4433 13475 4491 13481
rect 5169 13515 5227 13521
rect 5169 13481 5181 13515
rect 5215 13512 5227 13515
rect 7466 13512 7472 13524
rect 5215 13484 7052 13512
rect 7427 13484 7472 13512
rect 5215 13481 5227 13484
rect 5169 13475 5227 13481
rect 3050 13404 3056 13456
rect 3108 13444 3114 13456
rect 3421 13447 3479 13453
rect 3421 13444 3433 13447
rect 3108 13416 3433 13444
rect 3108 13404 3114 13416
rect 3421 13413 3433 13416
rect 3467 13413 3479 13447
rect 3421 13407 3479 13413
rect 5718 13404 5724 13456
rect 5776 13444 5782 13456
rect 5997 13447 6055 13453
rect 5997 13444 6009 13447
rect 5776 13416 6009 13444
rect 5776 13404 5782 13416
rect 5997 13413 6009 13416
rect 6043 13413 6055 13447
rect 5997 13407 6055 13413
rect 6086 13404 6092 13456
rect 6144 13444 6150 13456
rect 6549 13447 6607 13453
rect 6549 13444 6561 13447
rect 6144 13416 6561 13444
rect 6144 13404 6150 13416
rect 6549 13413 6561 13416
rect 6595 13413 6607 13447
rect 7024 13444 7052 13484
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 8754 13512 8760 13524
rect 8715 13484 8760 13512
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 9493 13515 9551 13521
rect 9493 13481 9505 13515
rect 9539 13512 9551 13515
rect 9674 13512 9680 13524
rect 9539 13484 9680 13512
rect 9539 13481 9551 13484
rect 9493 13475 9551 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10781 13515 10839 13521
rect 10781 13512 10793 13515
rect 10192 13484 10793 13512
rect 10192 13472 10198 13484
rect 10781 13481 10793 13484
rect 10827 13512 10839 13515
rect 12986 13512 12992 13524
rect 10827 13484 12992 13512
rect 10827 13481 10839 13484
rect 10781 13475 10839 13481
rect 12986 13472 12992 13484
rect 13044 13472 13050 13524
rect 8386 13444 8392 13456
rect 7024 13416 8392 13444
rect 6549 13407 6607 13413
rect 8386 13404 8392 13416
rect 8444 13404 8450 13456
rect 9858 13444 9864 13456
rect 9819 13416 9864 13444
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 9950 13404 9956 13456
rect 10008 13444 10014 13456
rect 11425 13447 11483 13453
rect 11425 13444 11437 13447
rect 10008 13416 11437 13444
rect 10008 13404 10014 13416
rect 11425 13413 11437 13416
rect 11471 13444 11483 13447
rect 11790 13444 11796 13456
rect 11471 13416 11796 13444
rect 11471 13413 11483 13416
rect 11425 13407 11483 13413
rect 11790 13404 11796 13416
rect 11848 13404 11854 13456
rect 2682 13376 2688 13388
rect 2643 13348 2688 13376
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 2866 13376 2872 13388
rect 2827 13348 2872 13376
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 6822 13336 6828 13388
rect 6880 13376 6886 13388
rect 7377 13379 7435 13385
rect 7377 13376 7389 13379
rect 6880 13348 7389 13376
rect 6880 13336 6886 13348
rect 7377 13345 7389 13348
rect 7423 13376 7435 13379
rect 7650 13376 7656 13388
rect 7423 13348 7656 13376
rect 7423 13345 7435 13348
rect 7377 13339 7435 13345
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 7834 13376 7840 13388
rect 7795 13348 7840 13376
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 3970 13308 3976 13320
rect 3191 13280 3976 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 3970 13268 3976 13280
rect 4028 13308 4034 13320
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 4028 13280 4077 13308
rect 4028 13268 4034 13280
rect 4065 13277 4077 13280
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 4890 13268 4896 13320
rect 4948 13308 4954 13320
rect 5350 13308 5356 13320
rect 4948 13280 5356 13308
rect 4948 13268 4954 13280
rect 5350 13268 5356 13280
rect 5408 13268 5414 13320
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13308 5963 13311
rect 6638 13308 6644 13320
rect 5951 13280 6644 13308
rect 5951 13277 5963 13280
rect 5905 13271 5963 13277
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 9766 13308 9772 13320
rect 9727 13280 9772 13308
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 10410 13308 10416 13320
rect 10323 13280 10416 13308
rect 10410 13268 10416 13280
rect 10468 13308 10474 13320
rect 11330 13308 11336 13320
rect 10468 13280 11336 13308
rect 10468 13268 10474 13280
rect 11330 13268 11336 13280
rect 11388 13268 11394 13320
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 11609 13311 11667 13317
rect 11609 13308 11621 13311
rect 11480 13280 11621 13308
rect 11480 13268 11486 13280
rect 11609 13277 11621 13280
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 11974 13268 11980 13320
rect 12032 13308 12038 13320
rect 12342 13308 12348 13320
rect 12032 13280 12348 13308
rect 12032 13268 12038 13280
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 3234 13200 3240 13252
rect 3292 13240 3298 13252
rect 3789 13243 3847 13249
rect 3789 13240 3801 13243
rect 3292 13212 3801 13240
rect 3292 13200 3298 13212
rect 3789 13209 3801 13212
rect 3835 13209 3847 13243
rect 3789 13203 3847 13209
rect 4430 13200 4436 13252
rect 4488 13240 4494 13252
rect 4985 13243 5043 13249
rect 4985 13240 4997 13243
rect 4488 13212 4997 13240
rect 4488 13200 4494 13212
rect 4985 13209 4997 13212
rect 5031 13240 5043 13243
rect 5994 13240 6000 13252
rect 5031 13212 6000 13240
rect 5031 13209 5043 13212
rect 4985 13203 5043 13209
rect 5994 13200 6000 13212
rect 6052 13200 6058 13252
rect 6730 13200 6736 13252
rect 6788 13240 6794 13252
rect 10226 13240 10232 13252
rect 6788 13212 10232 13240
rect 6788 13200 6794 13212
rect 10226 13200 10232 13212
rect 10284 13200 10290 13252
rect 1762 13132 1768 13184
rect 1820 13172 1826 13184
rect 1857 13175 1915 13181
rect 1857 13172 1869 13175
rect 1820 13144 1869 13172
rect 1820 13132 1826 13144
rect 1857 13141 1869 13144
rect 1903 13141 1915 13175
rect 2314 13172 2320 13184
rect 2275 13144 2320 13172
rect 1857 13135 1915 13141
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 3605 13175 3663 13181
rect 3605 13141 3617 13175
rect 3651 13172 3663 13175
rect 5169 13175 5227 13181
rect 5169 13172 5181 13175
rect 3651 13144 5181 13172
rect 3651 13141 3663 13144
rect 3605 13135 3663 13141
rect 5169 13141 5181 13144
rect 5215 13141 5227 13175
rect 5169 13135 5227 13141
rect 5350 13132 5356 13184
rect 5408 13172 5414 13184
rect 11974 13172 11980 13184
rect 5408 13144 11980 13172
rect 5408 13132 5414 13144
rect 11974 13132 11980 13144
rect 12032 13132 12038 13184
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 8941 12971 8999 12977
rect 8941 12968 8953 12971
rect 8720 12940 8953 12968
rect 8720 12928 8726 12940
rect 8941 12937 8953 12940
rect 8987 12937 8999 12971
rect 8941 12931 8999 12937
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 13587 12971 13645 12977
rect 13587 12968 13599 12971
rect 9824 12940 13599 12968
rect 9824 12928 9830 12940
rect 13587 12937 13599 12940
rect 13633 12937 13645 12971
rect 13906 12968 13912 12980
rect 13867 12940 13912 12968
rect 13587 12931 13645 12937
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12832 5043 12835
rect 5350 12832 5356 12844
rect 5031 12804 5356 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5350 12792 5356 12804
rect 5408 12832 5414 12844
rect 7466 12832 7472 12844
rect 5408 12804 7472 12832
rect 5408 12792 5414 12804
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12832 7803 12835
rect 8680 12832 8708 12928
rect 8757 12903 8815 12909
rect 8757 12869 8769 12903
rect 8803 12900 8815 12903
rect 8803 12872 11468 12900
rect 8803 12869 8815 12872
rect 8757 12863 8815 12869
rect 7791 12804 8708 12832
rect 9585 12835 9643 12841
rect 7791 12801 7803 12804
rect 7745 12795 7803 12801
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 10873 12835 10931 12841
rect 10873 12832 10885 12835
rect 9631 12804 10885 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 10873 12801 10885 12804
rect 10919 12832 10931 12835
rect 11195 12835 11253 12841
rect 11195 12832 11207 12835
rect 10919 12804 11207 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 11195 12801 11207 12804
rect 11241 12801 11253 12835
rect 11440 12832 11468 12872
rect 11790 12860 11796 12912
rect 11848 12900 11854 12912
rect 11885 12903 11943 12909
rect 11885 12900 11897 12903
rect 11848 12872 11897 12900
rect 11848 12860 11854 12872
rect 11885 12869 11897 12872
rect 11931 12869 11943 12903
rect 11885 12863 11943 12869
rect 12575 12835 12633 12841
rect 12575 12832 12587 12835
rect 11440 12804 12587 12832
rect 11195 12795 11253 12801
rect 12575 12801 12587 12804
rect 12621 12801 12633 12835
rect 12575 12795 12633 12801
rect 1765 12767 1823 12773
rect 1765 12733 1777 12767
rect 1811 12764 1823 12767
rect 2041 12767 2099 12773
rect 1811 12736 1992 12764
rect 1811 12733 1823 12736
rect 1765 12727 1823 12733
rect 1964 12628 1992 12736
rect 2041 12733 2053 12767
rect 2087 12764 2099 12767
rect 2314 12764 2320 12776
rect 2087 12736 2320 12764
rect 2087 12733 2099 12736
rect 2041 12727 2099 12733
rect 2314 12724 2320 12736
rect 2372 12764 2378 12776
rect 2866 12764 2872 12776
rect 2372 12736 2872 12764
rect 2372 12724 2378 12736
rect 2866 12724 2872 12736
rect 2924 12724 2930 12776
rect 3053 12767 3111 12773
rect 3053 12733 3065 12767
rect 3099 12764 3111 12767
rect 3142 12764 3148 12776
rect 3099 12736 3148 12764
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 3142 12724 3148 12736
rect 3200 12724 3206 12776
rect 7653 12767 7711 12773
rect 7653 12764 7665 12767
rect 5368 12736 7665 12764
rect 2222 12696 2228 12708
rect 2183 12668 2228 12696
rect 2222 12656 2228 12668
rect 2280 12656 2286 12708
rect 4341 12699 4399 12705
rect 4341 12696 4353 12699
rect 3436 12668 4353 12696
rect 2406 12628 2412 12640
rect 1964 12600 2412 12628
rect 2406 12588 2412 12600
rect 2464 12628 2470 12640
rect 2593 12631 2651 12637
rect 2593 12628 2605 12631
rect 2464 12600 2605 12628
rect 2464 12588 2470 12600
rect 2593 12597 2605 12600
rect 2639 12628 2651 12631
rect 2774 12628 2780 12640
rect 2639 12600 2780 12628
rect 2639 12597 2651 12600
rect 2593 12591 2651 12597
rect 2774 12588 2780 12600
rect 2832 12588 2838 12640
rect 3436 12637 3464 12668
rect 4341 12665 4353 12668
rect 4387 12696 4399 12699
rect 4430 12696 4436 12708
rect 4387 12668 4436 12696
rect 4387 12665 4399 12668
rect 4341 12659 4399 12665
rect 4430 12656 4436 12668
rect 4488 12696 4494 12708
rect 5368 12705 5396 12736
rect 7653 12733 7665 12736
rect 7699 12764 7711 12767
rect 8665 12767 8723 12773
rect 7699 12736 7972 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 7944 12708 7972 12736
rect 8665 12733 8677 12767
rect 8711 12733 8723 12767
rect 8665 12727 8723 12733
rect 4893 12699 4951 12705
rect 4893 12696 4905 12699
rect 4488 12668 4905 12696
rect 4488 12656 4494 12668
rect 4893 12665 4905 12668
rect 4939 12696 4951 12699
rect 5347 12699 5405 12705
rect 5347 12696 5359 12699
rect 4939 12668 5359 12696
rect 4939 12665 4951 12668
rect 4893 12659 4951 12665
rect 5347 12665 5359 12668
rect 5393 12665 5405 12699
rect 6638 12696 6644 12708
rect 6551 12668 6644 12696
rect 5347 12659 5405 12665
rect 6638 12656 6644 12668
rect 6696 12696 6702 12708
rect 6696 12668 7788 12696
rect 6696 12656 6702 12668
rect 2961 12631 3019 12637
rect 2961 12597 2973 12631
rect 3007 12628 3019 12631
rect 3421 12631 3479 12637
rect 3421 12628 3433 12631
rect 3007 12600 3433 12628
rect 3007 12597 3019 12600
rect 2961 12591 3019 12597
rect 3421 12597 3433 12600
rect 3467 12597 3479 12631
rect 3421 12591 3479 12597
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 4062 12628 4068 12640
rect 4019 12600 4068 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 5718 12588 5724 12640
rect 5776 12628 5782 12640
rect 5905 12631 5963 12637
rect 5905 12628 5917 12631
rect 5776 12600 5917 12628
rect 5776 12588 5782 12600
rect 5905 12597 5917 12600
rect 5951 12628 5963 12631
rect 6181 12631 6239 12637
rect 6181 12628 6193 12631
rect 5951 12600 6193 12628
rect 5951 12597 5963 12600
rect 5905 12591 5963 12597
rect 6181 12597 6193 12600
rect 6227 12597 6239 12631
rect 6181 12591 6239 12597
rect 6822 12588 6828 12640
rect 6880 12628 6886 12640
rect 7193 12631 7251 12637
rect 7193 12628 7205 12631
rect 6880 12600 7205 12628
rect 6880 12588 6886 12600
rect 7193 12597 7205 12600
rect 7239 12597 7251 12631
rect 7760 12628 7788 12668
rect 7926 12656 7932 12708
rect 7984 12696 7990 12708
rect 8066 12699 8124 12705
rect 8066 12696 8078 12699
rect 7984 12668 8078 12696
rect 7984 12656 7990 12668
rect 8066 12665 8078 12668
rect 8112 12665 8124 12699
rect 8680 12696 8708 12727
rect 10962 12724 10968 12776
rect 11020 12764 11026 12776
rect 11092 12767 11150 12773
rect 11092 12764 11104 12767
rect 11020 12736 11104 12764
rect 11020 12724 11026 12736
rect 11092 12733 11104 12736
rect 11138 12764 11150 12767
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 11138 12736 11529 12764
rect 11138 12733 11150 12736
rect 11092 12727 11150 12733
rect 11517 12733 11529 12736
rect 11563 12764 11575 12767
rect 12066 12764 12072 12776
rect 11563 12736 12072 12764
rect 11563 12733 11575 12736
rect 11517 12727 11575 12733
rect 12066 12724 12072 12736
rect 12124 12724 12130 12776
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 12472 12767 12530 12773
rect 12472 12764 12484 12767
rect 12216 12736 12484 12764
rect 12216 12724 12222 12736
rect 12472 12733 12484 12736
rect 12518 12764 12530 12767
rect 12894 12764 12900 12776
rect 12518 12736 12900 12764
rect 12518 12733 12530 12736
rect 12472 12727 12530 12733
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 13516 12767 13574 12773
rect 13516 12733 13528 12767
rect 13562 12764 13574 12767
rect 13722 12764 13728 12776
rect 13562 12736 13728 12764
rect 13562 12733 13574 12736
rect 13516 12727 13574 12733
rect 13722 12724 13728 12736
rect 13780 12764 13786 12776
rect 13906 12764 13912 12776
rect 13780 12736 13912 12764
rect 13780 12724 13786 12736
rect 13906 12724 13912 12736
rect 13964 12724 13970 12776
rect 9401 12699 9459 12705
rect 9401 12696 9413 12699
rect 8680 12668 9413 12696
rect 8066 12659 8124 12665
rect 9401 12665 9413 12668
rect 9447 12696 9459 12699
rect 9677 12699 9735 12705
rect 9677 12696 9689 12699
rect 9447 12668 9689 12696
rect 9447 12665 9459 12668
rect 9401 12659 9459 12665
rect 9677 12665 9689 12668
rect 9723 12665 9735 12699
rect 10226 12696 10232 12708
rect 10187 12668 10232 12696
rect 9677 12659 9735 12665
rect 8757 12631 8815 12637
rect 8757 12628 8769 12631
rect 7760 12600 8769 12628
rect 7193 12591 7251 12597
rect 8757 12597 8769 12600
rect 8803 12597 8815 12631
rect 9692 12628 9720 12659
rect 10226 12656 10232 12668
rect 10284 12656 10290 12708
rect 9858 12628 9864 12640
rect 9692 12600 9864 12628
rect 8757 12591 8815 12597
rect 9858 12588 9864 12600
rect 9916 12628 9922 12640
rect 10505 12631 10563 12637
rect 10505 12628 10517 12631
rect 9916 12600 10517 12628
rect 9916 12588 9922 12600
rect 10505 12597 10517 12600
rect 10551 12597 10563 12631
rect 10505 12591 10563 12597
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 2682 12384 2688 12436
rect 2740 12424 2746 12436
rect 2869 12427 2927 12433
rect 2869 12424 2881 12427
rect 2740 12396 2881 12424
rect 2740 12384 2746 12396
rect 2869 12393 2881 12396
rect 2915 12393 2927 12427
rect 2869 12387 2927 12393
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 3970 12424 3976 12436
rect 3927 12396 3976 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4430 12424 4436 12436
rect 4391 12396 4436 12424
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 4982 12424 4988 12436
rect 4943 12396 4988 12424
rect 4982 12384 4988 12396
rect 5040 12384 5046 12436
rect 5350 12424 5356 12436
rect 5311 12396 5356 12424
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 8757 12427 8815 12433
rect 8757 12393 8769 12427
rect 8803 12424 8815 12427
rect 9398 12424 9404 12436
rect 8803 12396 9404 12424
rect 8803 12393 8815 12396
rect 8757 12387 8815 12393
rect 9398 12384 9404 12396
rect 9456 12424 9462 12436
rect 9456 12396 9904 12424
rect 9456 12384 9462 12396
rect 2035 12359 2093 12365
rect 2035 12325 2047 12359
rect 2081 12356 2093 12359
rect 3326 12356 3332 12368
rect 2081 12328 3332 12356
rect 2081 12325 2093 12328
rect 2035 12319 2093 12325
rect 3326 12316 3332 12328
rect 3384 12316 3390 12368
rect 5994 12356 6000 12368
rect 5955 12328 6000 12356
rect 5994 12316 6000 12328
rect 6052 12316 6058 12368
rect 7926 12316 7932 12368
rect 7984 12356 7990 12368
rect 8158 12359 8216 12365
rect 8158 12356 8170 12359
rect 7984 12328 8170 12356
rect 7984 12316 7990 12328
rect 8158 12325 8170 12328
rect 8204 12325 8216 12359
rect 8158 12319 8216 12325
rect 9493 12359 9551 12365
rect 9493 12325 9505 12359
rect 9539 12356 9551 12359
rect 9766 12356 9772 12368
rect 9539 12328 9772 12356
rect 9539 12325 9551 12328
rect 9493 12319 9551 12325
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 9876 12365 9904 12396
rect 11330 12384 11336 12436
rect 11388 12424 11394 12436
rect 11701 12427 11759 12433
rect 11701 12424 11713 12427
rect 11388 12396 11713 12424
rect 11388 12384 11394 12396
rect 11701 12393 11713 12396
rect 11747 12393 11759 12427
rect 11701 12387 11759 12393
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 12391 12427 12449 12433
rect 12391 12424 12403 12427
rect 12032 12396 12403 12424
rect 12032 12384 12038 12396
rect 12391 12393 12403 12396
rect 12437 12393 12449 12427
rect 12391 12387 12449 12393
rect 9861 12359 9919 12365
rect 9861 12325 9873 12359
rect 9907 12325 9919 12359
rect 10410 12356 10416 12368
rect 10323 12328 10416 12356
rect 9861 12319 9919 12325
rect 10410 12316 10416 12328
rect 10468 12356 10474 12368
rect 11422 12356 11428 12368
rect 10468 12328 11428 12356
rect 10468 12316 10474 12328
rect 11422 12316 11428 12328
rect 11480 12316 11486 12368
rect 1486 12248 1492 12300
rect 1544 12288 1550 12300
rect 1762 12288 1768 12300
rect 1544 12260 1768 12288
rect 1544 12248 1550 12260
rect 1762 12248 1768 12260
rect 1820 12248 1826 12300
rect 2222 12248 2228 12300
rect 2280 12288 2286 12300
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 2280 12260 4077 12288
rect 2280 12248 2286 12260
rect 4065 12257 4077 12260
rect 4111 12288 4123 12291
rect 4246 12288 4252 12300
rect 4111 12260 4252 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 10870 12248 10876 12300
rect 10928 12288 10934 12300
rect 11276 12291 11334 12297
rect 11276 12288 11288 12291
rect 10928 12260 11288 12288
rect 10928 12248 10934 12260
rect 11276 12257 11288 12260
rect 11322 12257 11334 12291
rect 11276 12251 11334 12257
rect 12288 12291 12346 12297
rect 12288 12257 12300 12291
rect 12334 12257 12346 12291
rect 12288 12251 12346 12257
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 1854 12220 1860 12232
rect 1719 12192 1860 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 1854 12180 1860 12192
rect 1912 12180 1918 12232
rect 2866 12180 2872 12232
rect 2924 12220 2930 12232
rect 3145 12223 3203 12229
rect 3145 12220 3157 12223
rect 2924 12192 3157 12220
rect 2924 12180 2930 12192
rect 3145 12189 3157 12192
rect 3191 12220 3203 12223
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 3191 12192 3249 12220
rect 3191 12189 3203 12192
rect 3145 12183 3203 12189
rect 3237 12189 3249 12192
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 5905 12223 5963 12229
rect 5905 12189 5917 12223
rect 5951 12189 5963 12223
rect 6178 12220 6184 12232
rect 6139 12192 6184 12220
rect 5905 12183 5963 12189
rect 1762 12112 1768 12164
rect 1820 12152 1826 12164
rect 5629 12155 5687 12161
rect 5629 12152 5641 12155
rect 1820 12124 5641 12152
rect 1820 12112 1826 12124
rect 5629 12121 5641 12124
rect 5675 12152 5687 12155
rect 5920 12152 5948 12183
rect 6178 12180 6184 12192
rect 6236 12220 6242 12232
rect 6825 12223 6883 12229
rect 6825 12220 6837 12223
rect 6236 12192 6837 12220
rect 6236 12180 6242 12192
rect 6825 12189 6837 12192
rect 6871 12220 6883 12223
rect 6914 12220 6920 12232
rect 6871 12192 6920 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 7742 12180 7748 12232
rect 7800 12220 7806 12232
rect 7837 12223 7895 12229
rect 7837 12220 7849 12223
rect 7800 12192 7849 12220
rect 7800 12180 7806 12192
rect 7837 12189 7849 12192
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 9582 12180 9588 12232
rect 9640 12220 9646 12232
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 9640 12192 9781 12220
rect 9640 12180 9646 12192
rect 9769 12189 9781 12192
rect 9815 12220 9827 12223
rect 10226 12220 10232 12232
rect 9815 12192 10232 12220
rect 9815 12189 9827 12192
rect 9769 12183 9827 12189
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12303 12220 12331 12251
rect 12124 12192 12331 12220
rect 12124 12180 12130 12192
rect 5675 12124 5948 12152
rect 5675 12121 5687 12124
rect 5629 12115 5687 12121
rect 6086 12112 6092 12164
rect 6144 12152 6150 12164
rect 11379 12155 11437 12161
rect 11379 12152 11391 12155
rect 6144 12124 11391 12152
rect 6144 12112 6150 12124
rect 11379 12121 11391 12124
rect 11425 12121 11437 12155
rect 11379 12115 11437 12121
rect 2314 12044 2320 12096
rect 2372 12084 2378 12096
rect 2593 12087 2651 12093
rect 2593 12084 2605 12087
rect 2372 12056 2605 12084
rect 2372 12044 2378 12056
rect 2593 12053 2605 12056
rect 2639 12053 2651 12087
rect 2593 12047 2651 12053
rect 3145 12087 3203 12093
rect 3145 12053 3157 12087
rect 3191 12084 3203 12087
rect 7469 12087 7527 12093
rect 7469 12084 7481 12087
rect 3191 12056 7481 12084
rect 3191 12053 3203 12056
rect 3145 12047 3203 12053
rect 7469 12053 7481 12056
rect 7515 12084 7527 12087
rect 7834 12084 7840 12096
rect 7515 12056 7840 12084
rect 7515 12053 7527 12056
rect 7469 12047 7527 12053
rect 7834 12044 7840 12056
rect 7892 12084 7898 12096
rect 9858 12084 9864 12096
rect 7892 12056 9864 12084
rect 7892 12044 7898 12056
rect 9858 12044 9864 12056
rect 9916 12044 9922 12096
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 1578 11840 1584 11892
rect 1636 11880 1642 11892
rect 2038 11880 2044 11892
rect 1636 11852 2044 11880
rect 1636 11840 1642 11852
rect 2038 11840 2044 11852
rect 2096 11840 2102 11892
rect 3053 11883 3111 11889
rect 3053 11849 3065 11883
rect 3099 11880 3111 11883
rect 3326 11880 3332 11892
rect 3099 11852 3332 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 3326 11840 3332 11852
rect 3384 11880 3390 11892
rect 4430 11880 4436 11892
rect 3384 11852 4436 11880
rect 3384 11840 3390 11852
rect 4430 11840 4436 11852
rect 4488 11840 4494 11892
rect 4801 11883 4859 11889
rect 4801 11849 4813 11883
rect 4847 11880 4859 11883
rect 4982 11880 4988 11892
rect 4847 11852 4988 11880
rect 4847 11849 4859 11852
rect 4801 11843 4859 11849
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 5994 11880 6000 11892
rect 5955 11852 6000 11880
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 8478 11840 8484 11892
rect 8536 11880 8542 11892
rect 8665 11883 8723 11889
rect 8665 11880 8677 11883
rect 8536 11852 8677 11880
rect 8536 11840 8542 11852
rect 8665 11849 8677 11852
rect 8711 11849 8723 11883
rect 9490 11880 9496 11892
rect 9451 11852 9496 11880
rect 8665 11843 8723 11849
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 12066 11840 12072 11892
rect 12124 11880 12130 11892
rect 12897 11883 12955 11889
rect 12897 11880 12909 11883
rect 12124 11852 12909 11880
rect 12124 11840 12130 11852
rect 12897 11849 12909 11852
rect 12943 11880 12955 11883
rect 13078 11880 13084 11892
rect 12943 11852 13084 11880
rect 12943 11849 12955 11852
rect 12897 11843 12955 11849
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 4065 11815 4123 11821
rect 4065 11781 4077 11815
rect 4111 11812 4123 11815
rect 6549 11815 6607 11821
rect 6549 11812 6561 11815
rect 4111 11784 6561 11812
rect 4111 11781 4123 11784
rect 4065 11775 4123 11781
rect 6549 11781 6561 11784
rect 6595 11781 6607 11815
rect 6549 11775 6607 11781
rect 1394 11704 1400 11756
rect 1452 11744 1458 11756
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1452 11716 1685 11744
rect 1452 11704 1458 11716
rect 1673 11713 1685 11716
rect 1719 11744 1731 11747
rect 2593 11747 2651 11753
rect 2593 11744 2605 11747
rect 1719 11716 2605 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 2593 11713 2605 11716
rect 2639 11713 2651 11747
rect 2593 11707 2651 11713
rect 2958 11704 2964 11756
rect 3016 11744 3022 11756
rect 3145 11747 3203 11753
rect 3145 11744 3157 11747
rect 3016 11716 3157 11744
rect 3016 11704 3022 11716
rect 3145 11713 3157 11716
rect 3191 11713 3203 11747
rect 3145 11707 3203 11713
rect 4985 11747 5043 11753
rect 4985 11713 4997 11747
rect 5031 11744 5043 11747
rect 5166 11744 5172 11756
rect 5031 11716 5172 11744
rect 5031 11713 5043 11716
rect 4985 11707 5043 11713
rect 5166 11704 5172 11716
rect 5224 11744 5230 11756
rect 6086 11744 6092 11756
rect 5224 11716 6092 11744
rect 5224 11704 5230 11716
rect 6086 11704 6092 11716
rect 6144 11704 6150 11756
rect 2317 11679 2375 11685
rect 2317 11645 2329 11679
rect 2363 11676 2375 11679
rect 4430 11676 4436 11688
rect 2363 11648 4436 11676
rect 2363 11645 2375 11648
rect 2317 11639 2375 11645
rect 4430 11636 4436 11648
rect 4488 11636 4494 11688
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 5684 11648 5729 11676
rect 5684 11636 5690 11648
rect 1765 11611 1823 11617
rect 1765 11577 1777 11611
rect 1811 11608 1823 11611
rect 2130 11608 2136 11620
rect 1811 11580 2136 11608
rect 1811 11577 1823 11580
rect 1765 11571 1823 11577
rect 2130 11568 2136 11580
rect 2188 11568 2194 11620
rect 5074 11568 5080 11620
rect 5132 11608 5138 11620
rect 5132 11580 5177 11608
rect 5132 11568 5138 11580
rect 3326 11500 3332 11552
rect 3384 11540 3390 11552
rect 3513 11543 3571 11549
rect 3513 11540 3525 11543
rect 3384 11512 3525 11540
rect 3384 11500 3390 11512
rect 3513 11509 3525 11512
rect 3559 11509 3571 11543
rect 3513 11503 3571 11509
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 5644 11540 5672 11636
rect 6564 11608 6592 11775
rect 6914 11744 6920 11756
rect 6875 11716 6920 11744
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 7190 11744 7196 11756
rect 7151 11716 7196 11744
rect 7190 11704 7196 11716
rect 7248 11744 7254 11756
rect 8662 11744 8668 11756
rect 7248 11716 8668 11744
rect 7248 11704 7254 11716
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 9508 11744 9536 11840
rect 9508 11716 10456 11744
rect 8110 11636 8116 11688
rect 8168 11676 8174 11688
rect 10428 11685 10456 11716
rect 8481 11679 8539 11685
rect 8481 11676 8493 11679
rect 8168 11648 8493 11676
rect 8168 11636 8174 11648
rect 8481 11645 8493 11648
rect 8527 11645 8539 11679
rect 8481 11639 8539 11645
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 9953 11679 10011 11685
rect 9953 11676 9965 11679
rect 9723 11648 9965 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 9953 11645 9965 11648
rect 9999 11645 10011 11679
rect 9953 11639 10011 11645
rect 10413 11679 10471 11685
rect 10413 11645 10425 11679
rect 10459 11645 10471 11679
rect 10413 11639 10471 11645
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 12472 11679 12530 11685
rect 12472 11676 12484 11679
rect 12124 11648 12484 11676
rect 12124 11636 12130 11648
rect 12472 11645 12484 11648
rect 12518 11676 12530 11679
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 12518 11648 13277 11676
rect 12518 11645 12530 11648
rect 12472 11639 12530 11645
rect 13265 11645 13277 11648
rect 13311 11676 13323 11679
rect 13446 11676 13452 11688
rect 13311 11648 13452 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 7009 11611 7067 11617
rect 7009 11608 7021 11611
rect 6564 11580 7021 11608
rect 7009 11577 7021 11580
rect 7055 11577 7067 11611
rect 7009 11571 7067 11577
rect 7650 11568 7656 11620
rect 7708 11608 7714 11620
rect 12575 11611 12633 11617
rect 12575 11608 12587 11611
rect 7708 11580 12587 11608
rect 7708 11568 7714 11580
rect 12575 11577 12587 11580
rect 12621 11577 12633 11611
rect 12575 11571 12633 11577
rect 7926 11540 7932 11552
rect 4028 11512 5672 11540
rect 7887 11512 7932 11540
rect 4028 11500 4034 11512
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 8168 11512 8217 11540
rect 8168 11500 8174 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 8205 11503 8263 11509
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 9677 11543 9735 11549
rect 9677 11540 9689 11543
rect 9548 11512 9689 11540
rect 9548 11500 9554 11512
rect 9677 11509 9689 11512
rect 9723 11540 9735 11543
rect 9769 11543 9827 11549
rect 9769 11540 9781 11543
rect 9723 11512 9781 11540
rect 9723 11509 9735 11512
rect 9677 11503 9735 11509
rect 9769 11509 9781 11512
rect 9815 11509 9827 11543
rect 10042 11540 10048 11552
rect 10003 11512 10048 11540
rect 9769 11503 9827 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 10928 11512 11253 11540
rect 10928 11500 10934 11512
rect 11241 11509 11253 11512
rect 11287 11509 11299 11543
rect 11241 11503 11299 11509
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1762 11336 1768 11348
rect 1719 11308 1768 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1762 11296 1768 11308
rect 1820 11296 1826 11348
rect 2314 11336 2320 11348
rect 2275 11308 2320 11336
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 2958 11296 2964 11348
rect 3016 11336 3022 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 3016 11308 3433 11336
rect 3016 11296 3022 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 4246 11336 4252 11348
rect 4207 11308 4252 11336
rect 3421 11299 3479 11305
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 4985 11339 5043 11345
rect 4985 11305 4997 11339
rect 5031 11336 5043 11339
rect 5166 11336 5172 11348
rect 5031 11308 5172 11336
rect 5031 11305 5043 11308
rect 4985 11299 5043 11305
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 9398 11336 9404 11348
rect 9359 11308 9404 11336
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 9766 11336 9772 11348
rect 9727 11308 9772 11336
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 9858 11296 9864 11348
rect 9916 11336 9922 11348
rect 11425 11339 11483 11345
rect 11425 11336 11437 11339
rect 9916 11308 11437 11336
rect 9916 11296 9922 11308
rect 11425 11305 11437 11308
rect 11471 11305 11483 11339
rect 11425 11299 11483 11305
rect 3142 11268 3148 11280
rect 3103 11240 3148 11268
rect 3142 11228 3148 11240
rect 3200 11228 3206 11280
rect 5718 11268 5724 11280
rect 5679 11240 5724 11268
rect 5718 11228 5724 11240
rect 5776 11228 5782 11280
rect 6273 11271 6331 11277
rect 6273 11237 6285 11271
rect 6319 11268 6331 11271
rect 6914 11268 6920 11280
rect 6319 11240 6920 11268
rect 6319 11237 6331 11240
rect 6273 11231 6331 11237
rect 6914 11228 6920 11240
rect 6972 11228 6978 11280
rect 7926 11228 7932 11280
rect 7984 11268 7990 11280
rect 8199 11271 8257 11277
rect 8199 11268 8211 11271
rect 7984 11240 8211 11268
rect 7984 11228 7990 11240
rect 8199 11237 8211 11240
rect 8245 11268 8257 11271
rect 8386 11268 8392 11280
rect 8245 11240 8392 11268
rect 8245 11237 8257 11240
rect 8199 11231 8257 11237
rect 8386 11228 8392 11240
rect 8444 11228 8450 11280
rect 9125 11271 9183 11277
rect 9125 11237 9137 11271
rect 9171 11268 9183 11271
rect 9582 11268 9588 11280
rect 9171 11240 9588 11268
rect 9171 11237 9183 11240
rect 9125 11231 9183 11237
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 1464 11203 1522 11209
rect 1464 11169 1476 11203
rect 1510 11200 1522 11203
rect 1946 11200 1952 11212
rect 1510 11172 1952 11200
rect 1510 11169 1522 11172
rect 1464 11163 1522 11169
rect 1946 11160 1952 11172
rect 2004 11160 2010 11212
rect 2498 11200 2504 11212
rect 2459 11172 2504 11200
rect 2498 11160 2504 11172
rect 2556 11160 2562 11212
rect 2866 11200 2872 11212
rect 2827 11172 2872 11200
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 5258 11200 5264 11212
rect 4479 11172 5264 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 9950 11200 9956 11212
rect 9911 11172 9956 11200
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 1854 11092 1860 11144
rect 1912 11132 1918 11144
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 1912 11104 3801 11132
rect 1912 11092 1918 11104
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11132 5687 11135
rect 5994 11132 6000 11144
rect 5675 11104 6000 11132
rect 5675 11101 5687 11104
rect 5629 11095 5687 11101
rect 5994 11092 6000 11104
rect 6052 11132 6058 11144
rect 7650 11132 7656 11144
rect 6052 11104 7656 11132
rect 6052 11092 6058 11104
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 7834 11132 7840 11144
rect 7795 11104 7840 11132
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 9490 11092 9496 11144
rect 9548 11132 9554 11144
rect 10152 11132 10180 11163
rect 11054 11160 11060 11212
rect 11112 11200 11118 11212
rect 11241 11203 11299 11209
rect 11241 11200 11253 11203
rect 11112 11172 11253 11200
rect 11112 11160 11118 11172
rect 11241 11169 11253 11172
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11146 11132 11152 11144
rect 9548 11104 11152 11132
rect 9548 11092 9554 11104
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 2958 11024 2964 11076
rect 3016 11064 3022 11076
rect 4617 11067 4675 11073
rect 4617 11064 4629 11067
rect 3016 11036 4629 11064
rect 3016 11024 3022 11036
rect 4617 11033 4629 11036
rect 4663 11033 4675 11067
rect 4617 11027 4675 11033
rect 6917 11067 6975 11073
rect 6917 11033 6929 11067
rect 6963 11064 6975 11067
rect 7374 11064 7380 11076
rect 6963 11036 7380 11064
rect 6963 11033 6975 11036
rect 6917 11027 6975 11033
rect 7374 11024 7380 11036
rect 7432 11024 7438 11076
rect 7742 11064 7748 11076
rect 7655 11036 7748 11064
rect 7742 11024 7748 11036
rect 7800 11064 7806 11076
rect 10042 11064 10048 11076
rect 7800 11036 10048 11064
rect 7800 11024 7806 11036
rect 10042 11024 10048 11036
rect 10100 11024 10106 11076
rect 1949 10999 2007 11005
rect 1949 10965 1961 10999
rect 1995 10996 2007 10999
rect 3326 10996 3332 11008
rect 1995 10968 3332 10996
rect 1995 10965 2007 10968
rect 1949 10959 2007 10965
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 6822 10956 6828 11008
rect 6880 10996 6886 11008
rect 7193 10999 7251 11005
rect 7193 10996 7205 10999
rect 6880 10968 7205 10996
rect 6880 10956 6886 10968
rect 7193 10965 7205 10968
rect 7239 10965 7251 10999
rect 8754 10996 8760 11008
rect 8715 10968 8760 10996
rect 7193 10959 7251 10965
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 2498 10752 2504 10804
rect 2556 10792 2562 10804
rect 2777 10795 2835 10801
rect 2777 10792 2789 10795
rect 2556 10764 2789 10792
rect 2556 10752 2562 10764
rect 2777 10761 2789 10764
rect 2823 10761 2835 10795
rect 2777 10755 2835 10761
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4062 10792 4068 10804
rect 4019 10764 4068 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 5537 10795 5595 10801
rect 5537 10761 5549 10795
rect 5583 10792 5595 10795
rect 5718 10792 5724 10804
rect 5583 10764 5724 10792
rect 5583 10761 5595 10764
rect 5537 10755 5595 10761
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 9950 10792 9956 10804
rect 7984 10764 9956 10792
rect 7984 10752 7990 10764
rect 9950 10752 9956 10764
rect 10008 10792 10014 10804
rect 10229 10795 10287 10801
rect 10229 10792 10241 10795
rect 10008 10764 10241 10792
rect 10008 10752 10014 10764
rect 10229 10761 10241 10764
rect 10275 10761 10287 10795
rect 10229 10755 10287 10761
rect 10778 10752 10784 10804
rect 10836 10792 10842 10804
rect 10919 10795 10977 10801
rect 10919 10792 10931 10795
rect 10836 10764 10931 10792
rect 10836 10752 10842 10764
rect 10919 10761 10931 10764
rect 10965 10761 10977 10795
rect 10919 10755 10977 10761
rect 4890 10684 4896 10736
rect 4948 10724 4954 10736
rect 5813 10727 5871 10733
rect 5813 10724 5825 10727
rect 4948 10696 5825 10724
rect 4948 10684 4954 10696
rect 5813 10693 5825 10696
rect 5859 10693 5871 10727
rect 5813 10687 5871 10693
rect 8294 10684 8300 10736
rect 8352 10724 8358 10736
rect 10686 10724 10692 10736
rect 8352 10696 10692 10724
rect 8352 10684 8358 10696
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10656 3663 10659
rect 3970 10656 3976 10668
rect 3651 10628 3976 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 4430 10656 4436 10668
rect 4391 10628 4436 10656
rect 4430 10616 4436 10628
rect 4488 10616 4494 10668
rect 7834 10616 7840 10668
rect 7892 10656 7898 10668
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 7892 10628 7941 10656
rect 7892 10616 7898 10628
rect 7929 10625 7941 10628
rect 7975 10656 7987 10659
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 7975 10628 8585 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8573 10625 8585 10628
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 8662 10616 8668 10668
rect 8720 10656 8726 10668
rect 8720 10628 10272 10656
rect 8720 10616 8726 10628
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1636 10560 1777 10588
rect 1636 10548 1642 10560
rect 1765 10557 1777 10560
rect 1811 10557 1823 10591
rect 2222 10588 2228 10600
rect 2183 10560 2228 10588
rect 1765 10551 1823 10557
rect 2222 10548 2228 10560
rect 2280 10588 2286 10600
rect 2866 10588 2872 10600
rect 2280 10560 2872 10588
rect 2280 10548 2286 10560
rect 2866 10548 2872 10560
rect 2924 10588 2930 10600
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 2924 10560 3157 10588
rect 2924 10548 2930 10560
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 3145 10551 3203 10557
rect 1673 10523 1731 10529
rect 1673 10489 1685 10523
rect 1719 10520 1731 10523
rect 1946 10520 1952 10532
rect 1719 10492 1952 10520
rect 1719 10489 1731 10492
rect 1673 10483 1731 10489
rect 1946 10480 1952 10492
rect 2004 10480 2010 10532
rect 3988 10520 4016 10616
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10588 5687 10591
rect 6822 10588 6828 10600
rect 5675 10560 6224 10588
rect 6783 10560 6828 10588
rect 5675 10557 5687 10560
rect 5629 10551 5687 10557
rect 4146 10523 4204 10529
rect 4146 10520 4158 10523
rect 3988 10492 4158 10520
rect 4146 10489 4158 10492
rect 4192 10489 4204 10523
rect 4146 10483 4204 10489
rect 4246 10480 4252 10532
rect 4304 10520 4310 10532
rect 4304 10492 4349 10520
rect 4304 10480 4310 10492
rect 6196 10464 6224 10560
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7285 10591 7343 10597
rect 7285 10588 7297 10591
rect 7208 10560 7297 10588
rect 7208 10464 7236 10560
rect 7285 10557 7297 10560
rect 7331 10557 7343 10591
rect 7285 10551 7343 10557
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 7653 10591 7711 10597
rect 7653 10588 7665 10591
rect 7432 10560 7665 10588
rect 7432 10548 7438 10560
rect 7653 10557 7665 10560
rect 7699 10588 7711 10591
rect 8478 10588 8484 10600
rect 7699 10560 8484 10588
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 8478 10548 8484 10560
rect 8536 10548 8542 10600
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 8812 10560 9873 10588
rect 8812 10548 8818 10560
rect 9861 10557 9873 10560
rect 9907 10588 9919 10591
rect 10134 10588 10140 10600
rect 9907 10560 10140 10588
rect 9907 10557 9919 10560
rect 9861 10551 9919 10557
rect 10134 10548 10140 10560
rect 10192 10548 10198 10600
rect 10244 10588 10272 10628
rect 10848 10591 10906 10597
rect 10848 10588 10860 10591
rect 10244 10560 10860 10588
rect 10848 10557 10860 10560
rect 10894 10588 10906 10591
rect 11609 10591 11667 10597
rect 11609 10588 11621 10591
rect 10894 10560 11621 10588
rect 10894 10557 10906 10560
rect 10848 10551 10906 10557
rect 11609 10557 11621 10560
rect 11655 10557 11667 10591
rect 11609 10551 11667 10557
rect 9950 10520 9956 10532
rect 9911 10492 9956 10520
rect 9950 10480 9956 10492
rect 10008 10480 10014 10532
rect 1854 10452 1860 10464
rect 1815 10424 1860 10452
rect 1854 10412 1860 10424
rect 1912 10412 1918 10464
rect 5169 10455 5227 10461
rect 5169 10421 5181 10455
rect 5215 10452 5227 10455
rect 5258 10452 5264 10464
rect 5215 10424 5264 10452
rect 5215 10421 5227 10424
rect 5169 10415 5227 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 6178 10452 6184 10464
rect 6139 10424 6184 10452
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 6641 10455 6699 10461
rect 6641 10421 6653 10455
rect 6687 10452 6699 10455
rect 7190 10452 7196 10464
rect 6687 10424 7196 10452
rect 6687 10421 6699 10424
rect 6641 10415 6699 10421
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 8297 10455 8355 10461
rect 8297 10421 8309 10455
rect 8343 10452 8355 10455
rect 8386 10452 8392 10464
rect 8343 10424 8392 10452
rect 8343 10421 8355 10424
rect 8297 10415 8355 10421
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 9125 10455 9183 10461
rect 9125 10421 9137 10455
rect 9171 10452 9183 10455
rect 9490 10452 9496 10464
rect 9171 10424 9496 10452
rect 9171 10421 9183 10424
rect 9125 10415 9183 10421
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11241 10455 11299 10461
rect 11241 10452 11253 10455
rect 11112 10424 11253 10452
rect 11112 10412 11118 10424
rect 11241 10421 11253 10424
rect 11287 10421 11299 10455
rect 11241 10415 11299 10421
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 1857 10251 1915 10257
rect 1857 10217 1869 10251
rect 1903 10248 1915 10251
rect 2222 10248 2228 10260
rect 1903 10220 2228 10248
rect 1903 10217 1915 10220
rect 1857 10211 1915 10217
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 2590 10248 2596 10260
rect 2551 10220 2596 10248
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 4028 10220 4169 10248
rect 4028 10208 4034 10220
rect 4157 10217 4169 10220
rect 4203 10217 4215 10251
rect 5994 10248 6000 10260
rect 5955 10220 6000 10248
rect 4157 10211 4215 10217
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 8297 10251 8355 10257
rect 8297 10248 8309 10251
rect 8260 10220 8309 10248
rect 8260 10208 8266 10220
rect 8297 10217 8309 10220
rect 8343 10248 8355 10251
rect 9766 10248 9772 10260
rect 8343 10220 9772 10248
rect 8343 10217 8355 10220
rect 8297 10211 8355 10217
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 12250 10208 12256 10260
rect 12308 10248 12314 10260
rect 12391 10251 12449 10257
rect 12391 10248 12403 10251
rect 12308 10220 12403 10248
rect 12308 10208 12314 10220
rect 12391 10217 12403 10220
rect 12437 10217 12449 10251
rect 12391 10211 12449 10217
rect 1578 10140 1584 10192
rect 1636 10180 1642 10192
rect 2133 10183 2191 10189
rect 2133 10180 2145 10183
rect 1636 10152 2145 10180
rect 1636 10140 1642 10152
rect 2133 10149 2145 10152
rect 2179 10149 2191 10183
rect 2133 10143 2191 10149
rect 7650 10140 7656 10192
rect 7708 10180 7714 10192
rect 9306 10180 9312 10192
rect 7708 10152 9312 10180
rect 7708 10140 7714 10152
rect 9306 10140 9312 10152
rect 9364 10140 9370 10192
rect 9861 10183 9919 10189
rect 9861 10149 9873 10183
rect 9907 10180 9919 10183
rect 9950 10180 9956 10192
rect 9907 10152 9956 10180
rect 9907 10149 9919 10152
rect 9861 10143 9919 10149
rect 9950 10140 9956 10152
rect 10008 10140 10014 10192
rect 2593 10115 2651 10121
rect 2593 10081 2605 10115
rect 2639 10081 2651 10115
rect 2593 10075 2651 10081
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10112 2927 10115
rect 2958 10112 2964 10124
rect 2915 10084 2964 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 2608 10044 2636 10075
rect 2958 10072 2964 10084
rect 3016 10072 3022 10124
rect 4065 10115 4123 10121
rect 4065 10112 4077 10115
rect 3068 10084 4077 10112
rect 3068 10056 3096 10084
rect 4065 10081 4077 10084
rect 4111 10112 4123 10115
rect 4338 10112 4344 10124
rect 4111 10084 4344 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 4617 10115 4675 10121
rect 4617 10081 4629 10115
rect 4663 10081 4675 10115
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 4617 10075 4675 10081
rect 6380 10084 6561 10112
rect 3050 10044 3056 10056
rect 2608 10016 3056 10044
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 3881 10047 3939 10053
rect 3881 10013 3893 10047
rect 3927 10044 3939 10047
rect 4632 10044 4660 10075
rect 4890 10044 4896 10056
rect 3927 10016 4896 10044
rect 3927 10013 3939 10016
rect 3881 10007 3939 10013
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 5166 9908 5172 9920
rect 5127 9880 5172 9908
rect 5166 9868 5172 9880
rect 5224 9868 5230 9920
rect 5629 9911 5687 9917
rect 5629 9877 5641 9911
rect 5675 9908 5687 9911
rect 5902 9908 5908 9920
rect 5675 9880 5908 9908
rect 5675 9877 5687 9880
rect 5629 9871 5687 9877
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 6380 9917 6408 10084
rect 6549 10081 6561 10084
rect 6595 10112 6607 10115
rect 6822 10112 6828 10124
rect 6595 10084 6828 10112
rect 6595 10081 6607 10084
rect 6549 10075 6607 10081
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 7024 10084 7389 10112
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 7024 10044 7052 10084
rect 7377 10081 7389 10084
rect 7423 10112 7435 10115
rect 8110 10112 8116 10124
rect 7423 10084 8116 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 11238 10112 11244 10124
rect 11199 10084 11244 10112
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 12288 10115 12346 10121
rect 12288 10081 12300 10115
rect 12334 10081 12346 10115
rect 12288 10075 12346 10081
rect 6696 10016 7052 10044
rect 6696 10004 6702 10016
rect 7190 10004 7196 10056
rect 7248 10044 7254 10056
rect 7285 10047 7343 10053
rect 7285 10044 7297 10047
rect 7248 10016 7297 10044
rect 7248 10004 7254 10016
rect 7285 10013 7297 10016
rect 7331 10013 7343 10047
rect 7285 10007 7343 10013
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 9582 10044 9588 10056
rect 8619 10016 9588 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 9582 10004 9588 10016
rect 9640 10004 9646 10056
rect 9769 10047 9827 10053
rect 9769 10013 9781 10047
rect 9815 10013 9827 10047
rect 12303 10044 12331 10075
rect 12618 10044 12624 10056
rect 9769 10007 9827 10013
rect 10336 10016 12624 10044
rect 7466 9976 7472 9988
rect 7427 9948 7472 9976
rect 7466 9936 7472 9948
rect 7524 9936 7530 9988
rect 9674 9936 9680 9988
rect 9732 9976 9738 9988
rect 9784 9976 9812 10007
rect 10336 9988 10364 10016
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 10134 9976 10140 9988
rect 9732 9948 9812 9976
rect 9876 9948 10140 9976
rect 9732 9936 9738 9948
rect 6365 9911 6423 9917
rect 6365 9908 6377 9911
rect 6144 9880 6377 9908
rect 6144 9868 6150 9880
rect 6365 9877 6377 9880
rect 6411 9877 6423 9911
rect 6365 9871 6423 9877
rect 9309 9911 9367 9917
rect 9309 9877 9321 9911
rect 9355 9908 9367 9911
rect 9876 9908 9904 9948
rect 10134 9936 10140 9948
rect 10192 9936 10198 9988
rect 10318 9976 10324 9988
rect 10279 9948 10324 9976
rect 10318 9936 10324 9948
rect 10376 9936 10382 9988
rect 9355 9880 9904 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 10042 9868 10048 9920
rect 10100 9908 10106 9920
rect 10689 9911 10747 9917
rect 10689 9908 10701 9911
rect 10100 9880 10701 9908
rect 10100 9868 10106 9880
rect 10689 9877 10701 9880
rect 10735 9877 10747 9911
rect 10689 9871 10747 9877
rect 10778 9868 10784 9920
rect 10836 9908 10842 9920
rect 11379 9911 11437 9917
rect 11379 9908 11391 9911
rect 10836 9880 11391 9908
rect 10836 9868 10842 9880
rect 11379 9877 11391 9880
rect 11425 9877 11437 9911
rect 11379 9871 11437 9877
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 3050 9704 3056 9716
rect 3011 9676 3056 9704
rect 3050 9664 3056 9676
rect 3108 9664 3114 9716
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 4617 9707 4675 9713
rect 4617 9704 4629 9707
rect 4396 9676 4629 9704
rect 4396 9664 4402 9676
rect 4617 9673 4629 9676
rect 4663 9673 4675 9707
rect 4617 9667 4675 9673
rect 4706 9664 4712 9716
rect 4764 9704 4770 9716
rect 7101 9707 7159 9713
rect 7101 9704 7113 9707
rect 4764 9676 7113 9704
rect 4764 9664 4770 9676
rect 7101 9673 7113 9676
rect 7147 9673 7159 9707
rect 7101 9667 7159 9673
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 9950 9704 9956 9716
rect 9815 9676 9956 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 9950 9664 9956 9676
rect 10008 9664 10014 9716
rect 12618 9704 12624 9716
rect 12579 9676 12624 9704
rect 12618 9664 12624 9676
rect 12676 9664 12682 9716
rect 5166 9636 5172 9648
rect 5092 9608 5172 9636
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 2424 9540 3433 9568
rect 2424 9512 2452 9540
rect 3421 9537 3433 9540
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 2317 9503 2375 9509
rect 2317 9500 2329 9503
rect 1995 9472 2329 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2317 9469 2329 9472
rect 2363 9500 2375 9503
rect 2406 9500 2412 9512
rect 2363 9472 2412 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 2593 9503 2651 9509
rect 2593 9469 2605 9503
rect 2639 9500 2651 9503
rect 2958 9500 2964 9512
rect 2639 9472 2964 9500
rect 2639 9469 2651 9472
rect 2593 9463 2651 9469
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 3436 9500 3464 9531
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 3436 9472 3617 9500
rect 3605 9469 3617 9472
rect 3651 9469 3663 9503
rect 4062 9500 4068 9512
rect 4023 9472 4068 9500
rect 3605 9463 3663 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 5092 9500 5120 9608
rect 5166 9596 5172 9608
rect 5224 9636 5230 9648
rect 5997 9639 6055 9645
rect 5224 9596 5257 9636
rect 5997 9605 6009 9639
rect 6043 9636 6055 9639
rect 12526 9636 12532 9648
rect 6043 9608 12532 9636
rect 6043 9605 6055 9608
rect 5997 9599 6055 9605
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 5229 9568 5257 9596
rect 8202 9568 8208 9580
rect 5229 9540 6040 9568
rect 8163 9540 8208 9568
rect 6012 9512 6040 9540
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 10318 9568 10324 9580
rect 10279 9540 10324 9568
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 5157 9503 5215 9509
rect 5157 9500 5169 9503
rect 5092 9472 5169 9500
rect 5157 9469 5169 9472
rect 5203 9469 5215 9503
rect 5157 9463 5215 9469
rect 5261 9503 5319 9509
rect 5261 9469 5273 9503
rect 5307 9500 5319 9503
rect 5350 9500 5356 9512
rect 5307 9472 5356 9500
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 2682 9432 2688 9444
rect 1912 9404 2688 9432
rect 1912 9392 1918 9404
rect 2682 9392 2688 9404
rect 2740 9392 2746 9444
rect 4338 9432 4344 9444
rect 4299 9404 4344 9432
rect 4338 9392 4344 9404
rect 4396 9392 4402 9444
rect 5077 9435 5135 9441
rect 5077 9401 5089 9435
rect 5123 9432 5135 9435
rect 5276 9432 5304 9463
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 5445 9503 5503 9509
rect 5445 9469 5457 9503
rect 5491 9500 5503 9503
rect 5902 9500 5908 9512
rect 5491 9472 5908 9500
rect 5491 9469 5503 9472
rect 5445 9463 5503 9469
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 5994 9460 6000 9512
rect 6052 9500 6058 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 6052 9472 7021 9500
rect 6052 9460 6058 9472
rect 7009 9469 7021 9472
rect 7055 9500 7067 9503
rect 7653 9503 7711 9509
rect 7653 9500 7665 9503
rect 7055 9472 7665 9500
rect 7055 9469 7067 9472
rect 7009 9463 7067 9469
rect 7653 9469 7665 9472
rect 7699 9469 7711 9503
rect 7653 9463 7711 9469
rect 5123 9404 5304 9432
rect 6273 9435 6331 9441
rect 5123 9401 5135 9404
rect 5077 9395 5135 9401
rect 6273 9401 6285 9435
rect 6319 9432 6331 9435
rect 6825 9435 6883 9441
rect 6825 9432 6837 9435
rect 6319 9404 6837 9432
rect 6319 9401 6331 9404
rect 6273 9395 6331 9401
rect 6825 9401 6837 9404
rect 6871 9432 6883 9435
rect 7190 9432 7196 9444
rect 6871 9404 7196 9432
rect 6871 9401 6883 9404
rect 6825 9395 6883 9401
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 8386 9432 8392 9444
rect 8128 9404 8392 9432
rect 8128 9376 8156 9404
rect 8386 9392 8392 9404
rect 8444 9432 8450 9444
rect 8526 9435 8584 9441
rect 8526 9432 8538 9435
rect 8444 9404 8538 9432
rect 8444 9392 8450 9404
rect 8526 9401 8538 9404
rect 8572 9401 8584 9435
rect 10042 9432 10048 9444
rect 10003 9404 10048 9432
rect 8526 9395 8584 9401
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 10134 9392 10140 9444
rect 10192 9432 10198 9444
rect 10686 9432 10692 9444
rect 10192 9404 10692 9432
rect 10192 9392 10198 9404
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 2130 9364 2136 9376
rect 2091 9336 2136 9364
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 6638 9364 6644 9376
rect 6599 9336 6644 9364
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 8110 9364 8116 9376
rect 8071 9336 8116 9364
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 9125 9367 9183 9373
rect 9125 9333 9137 9367
rect 9171 9364 9183 9367
rect 9858 9364 9864 9376
rect 9171 9336 9864 9364
rect 9171 9333 9183 9336
rect 9125 9327 9183 9333
rect 9858 9324 9864 9336
rect 9916 9324 9922 9376
rect 11238 9364 11244 9376
rect 11199 9336 11244 9364
rect 11238 9324 11244 9336
rect 11296 9364 11302 9376
rect 11514 9364 11520 9376
rect 11296 9336 11520 9364
rect 11296 9324 11302 9336
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2498 9160 2504 9172
rect 2087 9132 2504 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 2498 9120 2504 9132
rect 2556 9160 2562 9172
rect 2958 9160 2964 9172
rect 2556 9132 2964 9160
rect 2556 9120 2562 9132
rect 2958 9120 2964 9132
rect 3016 9160 3022 9172
rect 3145 9163 3203 9169
rect 3145 9160 3157 9163
rect 3016 9132 3157 9160
rect 3016 9120 3022 9132
rect 3145 9129 3157 9132
rect 3191 9129 3203 9163
rect 3145 9123 3203 9129
rect 3697 9163 3755 9169
rect 3697 9129 3709 9163
rect 3743 9160 3755 9163
rect 4062 9160 4068 9172
rect 3743 9132 4068 9160
rect 3743 9129 3755 9132
rect 3697 9123 3755 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 7156 9132 7297 9160
rect 7156 9120 7162 9132
rect 7285 9129 7297 9132
rect 7331 9160 7343 9163
rect 7926 9160 7932 9172
rect 7331 9132 7932 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7926 9120 7932 9132
rect 7984 9120 7990 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 9674 9160 9680 9172
rect 9539 9132 9680 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 9674 9120 9680 9132
rect 9732 9160 9738 9172
rect 11241 9163 11299 9169
rect 11241 9160 11253 9163
rect 9732 9132 11253 9160
rect 9732 9120 9738 9132
rect 11241 9129 11253 9132
rect 11287 9129 11299 9163
rect 11241 9123 11299 9129
rect 2317 9095 2375 9101
rect 2317 9061 2329 9095
rect 2363 9092 2375 9095
rect 2682 9092 2688 9104
rect 2363 9064 2688 9092
rect 2363 9061 2375 9064
rect 2317 9055 2375 9061
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 4246 9092 4252 9104
rect 4207 9064 4252 9092
rect 4246 9052 4252 9064
rect 4304 9052 4310 9104
rect 7116 9092 7144 9120
rect 5552 9064 7144 9092
rect 7831 9095 7889 9101
rect 2222 8956 2228 8968
rect 2183 8928 2228 8956
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4430 8956 4436 8968
rect 4212 8928 4257 8956
rect 4391 8928 4436 8956
rect 4212 8916 4218 8928
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 2774 8888 2780 8900
rect 2735 8860 2780 8888
rect 2774 8848 2780 8860
rect 2832 8848 2838 8900
rect 3234 8848 3240 8900
rect 3292 8888 3298 8900
rect 5552 8888 5580 9064
rect 7831 9061 7843 9095
rect 7877 9092 7889 9095
rect 8110 9092 8116 9104
rect 7877 9064 8116 9092
rect 7877 9061 7889 9064
rect 7831 9055 7889 9061
rect 8110 9052 8116 9064
rect 8168 9052 8174 9104
rect 9582 9052 9588 9104
rect 9640 9092 9646 9104
rect 9769 9095 9827 9101
rect 9769 9092 9781 9095
rect 9640 9064 9781 9092
rect 9640 9052 9646 9064
rect 9769 9061 9781 9064
rect 9815 9061 9827 9095
rect 9769 9055 9827 9061
rect 9858 9052 9864 9104
rect 9916 9092 9922 9104
rect 10962 9092 10968 9104
rect 9916 9064 10968 9092
rect 9916 9052 9922 9064
rect 10962 9052 10968 9064
rect 11020 9052 11026 9104
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 8993 5687 9027
rect 5902 9024 5908 9036
rect 5863 8996 5908 9024
rect 5629 8987 5687 8993
rect 5644 8956 5672 8987
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 6365 9027 6423 9033
rect 6365 8993 6377 9027
rect 6411 9024 6423 9027
rect 6730 9024 6736 9036
rect 6411 8996 6736 9024
rect 6411 8993 6423 8996
rect 6365 8987 6423 8993
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 7466 9024 7472 9036
rect 7427 8996 7472 9024
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 10686 9024 10692 9036
rect 10468 8996 10513 9024
rect 10647 8996 10692 9024
rect 10468 8984 10474 8996
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 12288 9027 12346 9033
rect 12288 9024 12300 9027
rect 12216 8996 12300 9024
rect 12216 8984 12222 8996
rect 12288 8993 12300 8996
rect 12334 8993 12346 9027
rect 12288 8987 12346 8993
rect 5994 8956 6000 8968
rect 5644 8928 6000 8956
rect 5994 8916 6000 8928
rect 6052 8916 6058 8968
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 8536 8928 8769 8956
rect 8536 8916 8542 8928
rect 8757 8925 8769 8928
rect 8803 8956 8815 8959
rect 10778 8956 10784 8968
rect 8803 8928 10784 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 10778 8916 10784 8928
rect 10836 8916 10842 8968
rect 12434 8956 12440 8968
rect 12406 8916 12440 8956
rect 12492 8916 12498 8968
rect 5718 8888 5724 8900
rect 3292 8860 5580 8888
rect 5679 8860 5724 8888
rect 3292 8848 3298 8860
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 4890 8820 4896 8832
rect 4120 8792 4896 8820
rect 4120 8780 4126 8792
rect 4890 8780 4896 8792
rect 4948 8820 4954 8832
rect 5166 8820 5172 8832
rect 4948 8792 5172 8820
rect 4948 8780 4954 8792
rect 5166 8780 5172 8792
rect 5224 8780 5230 8832
rect 5350 8820 5356 8832
rect 5311 8792 5356 8820
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 6917 8823 6975 8829
rect 6917 8789 6929 8823
rect 6963 8820 6975 8823
rect 7190 8820 7196 8832
rect 6963 8792 7196 8820
rect 6963 8789 6975 8792
rect 6917 8783 6975 8789
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 8386 8820 8392 8832
rect 8347 8792 8392 8820
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 12406 8829 12434 8916
rect 12391 8823 12449 8829
rect 12391 8789 12403 8823
rect 12437 8789 12449 8823
rect 12391 8783 12449 8789
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 4246 8576 4252 8628
rect 4304 8616 4310 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 4304 8588 4445 8616
rect 4304 8576 4310 8588
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 4433 8579 4491 8585
rect 4893 8619 4951 8625
rect 4893 8585 4905 8619
rect 4939 8616 4951 8619
rect 5902 8616 5908 8628
rect 4939 8588 5908 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 6457 8619 6515 8625
rect 6457 8585 6469 8619
rect 6503 8616 6515 8619
rect 7282 8616 7288 8628
rect 6503 8588 7288 8616
rect 6503 8585 6515 8588
rect 6457 8579 6515 8585
rect 7282 8576 7288 8588
rect 7340 8576 7346 8628
rect 7929 8619 7987 8625
rect 7929 8585 7941 8619
rect 7975 8616 7987 8619
rect 8110 8616 8116 8628
rect 7975 8588 8116 8616
rect 7975 8585 7987 8588
rect 7929 8579 7987 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 9493 8619 9551 8625
rect 9493 8585 9505 8619
rect 9539 8616 9551 8619
rect 9582 8616 9588 8628
rect 9539 8588 9588 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 10962 8616 10968 8628
rect 10923 8588 10968 8616
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 5074 8508 5080 8560
rect 5132 8548 5138 8560
rect 5442 8548 5448 8560
rect 5132 8520 5448 8548
rect 5132 8508 5138 8520
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 5718 8508 5724 8560
rect 5776 8548 5782 8560
rect 6181 8551 6239 8557
rect 6181 8548 6193 8551
rect 5776 8520 6193 8548
rect 5776 8508 5782 8520
rect 6181 8517 6193 8520
rect 6227 8548 6239 8551
rect 7834 8548 7840 8560
rect 6227 8520 7840 8548
rect 6227 8517 6239 8520
rect 6181 8511 6239 8517
rect 7834 8508 7840 8520
rect 7892 8508 7898 8560
rect 11238 8548 11244 8560
rect 8173 8520 11244 8548
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5905 8483 5963 8489
rect 5307 8452 5580 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8412 1823 8415
rect 1946 8412 1952 8424
rect 1811 8384 1952 8412
rect 1811 8381 1823 8384
rect 1765 8375 1823 8381
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2406 8412 2412 8424
rect 2056 8384 2412 8412
rect 1673 8347 1731 8353
rect 1673 8313 1685 8347
rect 1719 8344 1731 8347
rect 2056 8344 2084 8384
rect 2406 8372 2412 8384
rect 2464 8412 2470 8424
rect 3326 8412 3332 8424
rect 2464 8384 3332 8412
rect 2464 8372 2470 8384
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 3510 8412 3516 8424
rect 3423 8384 3516 8412
rect 3510 8372 3516 8384
rect 3568 8412 3574 8424
rect 5552 8421 5580 8452
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 8173 8480 8201 8520
rect 11238 8508 11244 8520
rect 11296 8508 11302 8560
rect 8478 8480 8484 8492
rect 5951 8452 8201 8480
rect 8439 8452 8484 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8480 9183 8483
rect 10042 8480 10048 8492
rect 9171 8452 10048 8480
rect 9171 8449 9183 8452
rect 9125 8443 9183 8449
rect 10042 8440 10048 8452
rect 10100 8480 10106 8492
rect 10321 8483 10379 8489
rect 10321 8480 10333 8483
rect 10100 8452 10333 8480
rect 10100 8440 10106 8452
rect 10321 8449 10333 8452
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 10410 8440 10416 8492
rect 10468 8480 10474 8492
rect 12158 8480 12164 8492
rect 10468 8452 12164 8480
rect 10468 8440 10474 8452
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 5537 8415 5595 8421
rect 3568 8384 5488 8412
rect 3568 8372 3574 8384
rect 1719 8316 2084 8344
rect 1719 8313 1731 8316
rect 1673 8307 1731 8313
rect 2056 8276 2084 8316
rect 2222 8304 2228 8356
rect 2280 8344 2286 8356
rect 2961 8347 3019 8353
rect 2961 8344 2973 8347
rect 2280 8316 2973 8344
rect 2280 8304 2286 8316
rect 2961 8313 2973 8316
rect 3007 8313 3019 8347
rect 3344 8344 3372 8372
rect 3834 8347 3892 8353
rect 3834 8344 3846 8347
rect 3344 8316 3846 8344
rect 2961 8307 3019 8313
rect 3834 8313 3846 8316
rect 3880 8313 3892 8347
rect 5350 8344 5356 8356
rect 5311 8316 5356 8344
rect 3834 8307 3892 8313
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 5460 8344 5488 8384
rect 5537 8381 5549 8415
rect 5583 8412 5595 8415
rect 7098 8412 7104 8424
rect 5583 8384 6960 8412
rect 7059 8384 7104 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 6932 8344 6960 8384
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7282 8412 7288 8424
rect 7243 8384 7288 8412
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 12342 8372 12348 8424
rect 12400 8412 12406 8424
rect 12472 8415 12530 8421
rect 12472 8412 12484 8415
rect 12400 8384 12484 8412
rect 12400 8372 12406 8384
rect 12472 8381 12484 8384
rect 12518 8412 12530 8415
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12518 8384 12909 8412
rect 12518 8381 12530 8384
rect 12472 8375 12530 8381
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 8110 8344 8116 8356
rect 5460 8316 6868 8344
rect 6932 8316 8116 8344
rect 2133 8279 2191 8285
rect 2133 8276 2145 8279
rect 2056 8248 2145 8276
rect 2133 8245 2145 8248
rect 2179 8245 2191 8279
rect 2682 8276 2688 8288
rect 2643 8248 2688 8276
rect 2133 8239 2191 8245
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 4246 8276 4252 8288
rect 4028 8248 4252 8276
rect 4028 8236 4034 8248
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5442 8276 5448 8288
rect 5224 8248 5448 8276
rect 5224 8236 5230 8248
rect 5442 8236 5448 8248
rect 5500 8276 5506 8288
rect 6457 8279 6515 8285
rect 6457 8276 6469 8279
rect 5500 8248 6469 8276
rect 5500 8236 5506 8248
rect 6457 8245 6469 8248
rect 6503 8276 6515 8279
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 6503 8248 6561 8276
rect 6503 8245 6515 8248
rect 6457 8239 6515 8245
rect 6549 8245 6561 8248
rect 6595 8245 6607 8279
rect 6840 8276 6868 8316
rect 8110 8304 8116 8316
rect 8168 8304 8174 8356
rect 8573 8347 8631 8353
rect 8573 8313 8585 8347
rect 8619 8313 8631 8347
rect 10042 8344 10048 8356
rect 10003 8316 10048 8344
rect 8573 8307 8631 8313
rect 6917 8279 6975 8285
rect 6917 8276 6929 8279
rect 6840 8248 6929 8276
rect 6549 8239 6607 8245
rect 6917 8245 6929 8248
rect 6963 8245 6975 8279
rect 6917 8239 6975 8245
rect 7926 8236 7932 8288
rect 7984 8276 7990 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7984 8248 8217 8276
rect 7984 8236 7990 8248
rect 8205 8245 8217 8248
rect 8251 8276 8263 8279
rect 8386 8276 8392 8288
rect 8251 8248 8392 8276
rect 8251 8245 8263 8248
rect 8205 8239 8263 8245
rect 8386 8236 8392 8248
rect 8444 8276 8450 8288
rect 8588 8276 8616 8307
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 10137 8347 10195 8353
rect 10137 8313 10149 8347
rect 10183 8313 10195 8347
rect 10137 8307 10195 8313
rect 9766 8276 9772 8288
rect 8444 8248 8616 8276
rect 9727 8248 9772 8276
rect 8444 8236 8450 8248
rect 9766 8236 9772 8248
rect 9824 8276 9830 8288
rect 10152 8276 10180 8307
rect 9824 8248 10180 8276
rect 9824 8236 9830 8248
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 12575 8279 12633 8285
rect 12575 8276 12587 8279
rect 12308 8248 12587 8276
rect 12308 8236 12314 8248
rect 12575 8245 12587 8248
rect 12621 8245 12633 8279
rect 12575 8239 12633 8245
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 2133 8075 2191 8081
rect 2133 8041 2145 8075
rect 2179 8072 2191 8075
rect 2682 8072 2688 8084
rect 2179 8044 2688 8072
rect 2179 8041 2191 8044
rect 2133 8035 2191 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 3510 8072 3516 8084
rect 3471 8044 3516 8072
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 3970 8072 3976 8084
rect 3927 8044 3976 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 4212 8044 4261 8072
rect 4212 8032 4218 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4890 8072 4896 8084
rect 4851 8044 4896 8072
rect 4249 8035 4307 8041
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 6178 8032 6184 8084
rect 6236 8072 6242 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6236 8044 6745 8072
rect 6236 8032 6242 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 7466 8072 7472 8084
rect 7427 8044 7472 8072
rect 6733 8035 6791 8041
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 7576 8044 9904 8072
rect 2406 7964 2412 8016
rect 2464 8004 2470 8016
rect 2546 8007 2604 8013
rect 2546 8004 2558 8007
rect 2464 7976 2558 8004
rect 2464 7964 2470 7976
rect 2546 7973 2558 7976
rect 2592 7973 2604 8007
rect 2546 7967 2604 7973
rect 5258 7964 5264 8016
rect 5316 8004 5322 8016
rect 7576 8004 7604 8044
rect 5316 7976 7604 8004
rect 8757 8007 8815 8013
rect 5316 7964 5322 7976
rect 8757 7973 8769 8007
rect 8803 8004 8815 8007
rect 9766 8004 9772 8016
rect 8803 7976 9772 8004
rect 8803 7973 8815 7976
rect 8757 7967 8815 7973
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 9876 8004 9904 8044
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10781 8075 10839 8081
rect 10781 8072 10793 8075
rect 10100 8044 10793 8072
rect 10100 8032 10106 8044
rect 10781 8041 10793 8044
rect 10827 8072 10839 8075
rect 12250 8072 12256 8084
rect 10827 8044 12256 8072
rect 10827 8041 10839 8044
rect 10781 8035 10839 8041
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 10413 8007 10471 8013
rect 10413 8004 10425 8007
rect 9876 7976 10425 8004
rect 10413 7973 10425 7976
rect 10459 7973 10471 8007
rect 10413 7967 10471 7973
rect 2130 7896 2136 7948
rect 2188 7936 2194 7948
rect 2225 7939 2283 7945
rect 2225 7936 2237 7939
rect 2188 7908 2237 7936
rect 2188 7896 2194 7908
rect 2225 7905 2237 7908
rect 2271 7905 2283 7939
rect 2225 7899 2283 7905
rect 4062 7896 4068 7948
rect 4120 7936 4126 7948
rect 4525 7939 4583 7945
rect 4525 7936 4537 7939
rect 4120 7908 4537 7936
rect 4120 7896 4126 7908
rect 4525 7905 4537 7908
rect 4571 7905 4583 7939
rect 4525 7899 4583 7905
rect 6086 7896 6092 7948
rect 6144 7936 6150 7948
rect 6273 7939 6331 7945
rect 6273 7936 6285 7939
rect 6144 7908 6285 7936
rect 6144 7896 6150 7908
rect 6273 7905 6285 7908
rect 6319 7905 6331 7939
rect 6546 7936 6552 7948
rect 6507 7908 6552 7936
rect 6273 7899 6331 7905
rect 6546 7896 6552 7908
rect 6604 7896 6610 7948
rect 7926 7896 7932 7948
rect 7984 7936 7990 7948
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 7984 7908 8125 7936
rect 7984 7896 7990 7908
rect 8113 7905 8125 7908
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 9490 7896 9496 7948
rect 9548 7936 9554 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9548 7908 9689 7936
rect 9548 7896 9554 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 9953 7939 10011 7945
rect 9953 7905 9965 7939
rect 9999 7936 10011 7939
rect 10502 7936 10508 7948
rect 9999 7908 10508 7936
rect 9999 7905 10011 7908
rect 9953 7899 10011 7905
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 5408 7840 6408 7868
rect 5408 7828 5414 7840
rect 6380 7812 6408 7840
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 9968 7868 9996 7899
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 11238 7936 11244 7948
rect 11199 7908 11244 7936
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 6788 7840 9996 7868
rect 6788 7828 6794 7840
rect 5445 7803 5503 7809
rect 5445 7769 5457 7803
rect 5491 7800 5503 7803
rect 5491 7772 6316 7800
rect 5491 7769 5503 7772
rect 5445 7763 5503 7769
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7732 1823 7735
rect 1946 7732 1952 7744
rect 1811 7704 1952 7732
rect 1811 7701 1823 7704
rect 1765 7695 1823 7701
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 3142 7732 3148 7744
rect 3103 7704 3148 7732
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7732 5871 7735
rect 5994 7732 6000 7744
rect 5859 7704 6000 7732
rect 5859 7701 5871 7704
rect 5813 7695 5871 7701
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 6178 7732 6184 7744
rect 6139 7704 6184 7732
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 6288 7732 6316 7772
rect 6362 7760 6368 7812
rect 6420 7800 6426 7812
rect 9766 7800 9772 7812
rect 6420 7772 6465 7800
rect 9727 7772 9772 7800
rect 6420 7760 6426 7772
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 7098 7732 7104 7744
rect 6288 7704 7104 7732
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 7190 7692 7196 7744
rect 7248 7732 7254 7744
rect 11425 7735 11483 7741
rect 11425 7732 11437 7735
rect 7248 7704 11437 7732
rect 7248 7692 7254 7704
rect 11425 7701 11437 7704
rect 11471 7701 11483 7735
rect 11425 7695 11483 7701
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 5997 7531 6055 7537
rect 5997 7528 6009 7531
rect 5960 7500 6009 7528
rect 5960 7488 5966 7500
rect 5997 7497 6009 7500
rect 6043 7528 6055 7531
rect 6546 7528 6552 7540
rect 6043 7500 6552 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6546 7488 6552 7500
rect 6604 7528 6610 7540
rect 6730 7528 6736 7540
rect 6604 7500 6736 7528
rect 6604 7488 6610 7500
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7926 7528 7932 7540
rect 7887 7500 7932 7528
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 11238 7528 11244 7540
rect 11199 7500 11244 7528
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 6362 7460 6368 7472
rect 6275 7432 6368 7460
rect 6362 7420 6368 7432
rect 6420 7460 6426 7472
rect 6420 7432 7512 7460
rect 6420 7420 6426 7432
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 2222 7392 2228 7404
rect 1627 7364 2228 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 2590 7392 2596 7404
rect 2551 7364 2596 7392
rect 2590 7352 2596 7364
rect 2648 7392 2654 7404
rect 3789 7395 3847 7401
rect 3789 7392 3801 7395
rect 2648 7364 3801 7392
rect 2648 7352 2654 7364
rect 3789 7361 3801 7364
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 4338 7352 4344 7404
rect 4396 7392 4402 7404
rect 4525 7395 4583 7401
rect 4525 7392 4537 7395
rect 4396 7364 4537 7392
rect 4396 7352 4402 7364
rect 4525 7361 4537 7364
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 6178 7352 6184 7404
rect 6236 7392 6242 7404
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 6236 7364 6929 7392
rect 6236 7352 6242 7364
rect 6917 7361 6929 7364
rect 6963 7392 6975 7395
rect 7374 7392 7380 7404
rect 6963 7364 7380 7392
rect 6963 7361 6975 7364
rect 6917 7355 6975 7361
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 7484 7392 7512 7432
rect 7834 7420 7840 7472
rect 7892 7460 7898 7472
rect 8205 7463 8263 7469
rect 8205 7460 8217 7463
rect 7892 7432 8217 7460
rect 7892 7420 7898 7432
rect 8205 7429 8217 7432
rect 8251 7460 8263 7463
rect 8251 7432 8524 7460
rect 8251 7429 8263 7432
rect 8205 7423 8263 7429
rect 8389 7395 8447 7401
rect 8389 7392 8401 7395
rect 7484 7364 8401 7392
rect 8389 7361 8401 7364
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 8496 7333 8524 7432
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 9677 7327 9735 7333
rect 9677 7324 9689 7327
rect 8527 7296 9689 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 9677 7293 9689 7296
rect 9723 7324 9735 7327
rect 9766 7324 9772 7336
rect 9723 7296 9772 7324
rect 9723 7293 9735 7296
rect 9677 7287 9735 7293
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7293 10103 7327
rect 10045 7287 10103 7293
rect 4890 7265 4896 7268
rect 2914 7259 2972 7265
rect 2914 7256 2926 7259
rect 2424 7228 2926 7256
rect 2424 7200 2452 7228
rect 2914 7225 2926 7228
rect 2960 7225 2972 7259
rect 4846 7259 4896 7265
rect 4846 7256 4858 7259
rect 2914 7219 2972 7225
rect 4356 7228 4858 7256
rect 2133 7191 2191 7197
rect 2133 7157 2145 7191
rect 2179 7188 2191 7191
rect 2406 7188 2412 7200
rect 2179 7160 2412 7188
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 3510 7188 3516 7200
rect 3471 7160 3516 7188
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4356 7197 4384 7228
rect 4846 7225 4858 7228
rect 4892 7225 4896 7259
rect 4846 7219 4896 7225
rect 4890 7216 4896 7219
rect 4948 7216 4954 7268
rect 6178 7216 6184 7268
rect 6236 7256 6242 7268
rect 6638 7256 6644 7268
rect 6236 7228 6644 7256
rect 6236 7216 6242 7228
rect 6638 7216 6644 7228
rect 6696 7216 6702 7268
rect 7009 7259 7067 7265
rect 7009 7225 7021 7259
rect 7055 7256 7067 7259
rect 7098 7256 7104 7268
rect 7055 7228 7104 7256
rect 7055 7225 7067 7228
rect 7009 7219 7067 7225
rect 7098 7216 7104 7228
rect 7156 7216 7162 7268
rect 7282 7216 7288 7268
rect 7340 7256 7346 7268
rect 7561 7259 7619 7265
rect 7561 7256 7573 7259
rect 7340 7228 7573 7256
rect 7340 7216 7346 7228
rect 7561 7225 7573 7228
rect 7607 7225 7619 7259
rect 7561 7219 7619 7225
rect 8110 7216 8116 7268
rect 8168 7256 8174 7268
rect 9306 7256 9312 7268
rect 8168 7228 9312 7256
rect 8168 7216 8174 7228
rect 9306 7216 9312 7228
rect 9364 7256 9370 7268
rect 10060 7256 10088 7287
rect 10134 7256 10140 7268
rect 9364 7228 10140 7256
rect 9364 7216 9370 7228
rect 10134 7216 10140 7228
rect 10192 7216 10198 7268
rect 4341 7191 4399 7197
rect 4341 7188 4353 7191
rect 4304 7160 4353 7188
rect 4304 7148 4310 7160
rect 4341 7157 4353 7160
rect 4387 7157 4399 7191
rect 5442 7188 5448 7200
rect 5403 7160 5448 7188
rect 4341 7151 4399 7157
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 10413 7191 10471 7197
rect 10413 7157 10425 7191
rect 10459 7188 10471 7191
rect 10502 7188 10508 7200
rect 10459 7160 10508 7188
rect 10459 7157 10471 7160
rect 10413 7151 10471 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 2130 6944 2136 6996
rect 2188 6984 2194 6996
rect 2225 6987 2283 6993
rect 2225 6984 2237 6987
rect 2188 6956 2237 6984
rect 2188 6944 2194 6956
rect 2225 6953 2237 6956
rect 2271 6953 2283 6987
rect 3234 6984 3240 6996
rect 2225 6947 2283 6953
rect 2332 6956 3240 6984
rect 1302 6876 1308 6928
rect 1360 6916 1366 6928
rect 1535 6919 1593 6925
rect 1535 6916 1547 6919
rect 1360 6888 1547 6916
rect 1360 6876 1366 6888
rect 1535 6885 1547 6888
rect 1581 6885 1593 6919
rect 1535 6879 1593 6885
rect 1762 6876 1768 6928
rect 1820 6916 1826 6928
rect 1949 6919 2007 6925
rect 1949 6916 1961 6919
rect 1820 6888 1961 6916
rect 1820 6876 1826 6888
rect 1949 6885 1961 6888
rect 1995 6916 2007 6919
rect 2332 6916 2360 6956
rect 3234 6944 3240 6956
rect 3292 6944 3298 6996
rect 4065 6987 4123 6993
rect 4065 6953 4077 6987
rect 4111 6984 4123 6987
rect 4154 6984 4160 6996
rect 4111 6956 4160 6984
rect 4111 6953 4123 6956
rect 4065 6947 4123 6953
rect 4154 6944 4160 6956
rect 4212 6944 4218 6996
rect 4338 6944 4344 6996
rect 4396 6984 4402 6996
rect 4893 6987 4951 6993
rect 4893 6984 4905 6987
rect 4396 6956 4905 6984
rect 4396 6944 4402 6956
rect 4893 6953 4905 6956
rect 4939 6953 4951 6987
rect 4893 6947 4951 6953
rect 6917 6987 6975 6993
rect 6917 6953 6929 6987
rect 6963 6984 6975 6987
rect 7098 6984 7104 6996
rect 6963 6956 7104 6984
rect 6963 6953 6975 6956
rect 6917 6947 6975 6953
rect 7098 6944 7104 6956
rect 7156 6944 7162 6996
rect 9490 6984 9496 6996
rect 9451 6956 9496 6984
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 9861 6987 9919 6993
rect 9861 6984 9873 6987
rect 9640 6956 9873 6984
rect 9640 6944 9646 6956
rect 9861 6953 9873 6956
rect 9907 6953 9919 6987
rect 10134 6984 10140 6996
rect 10095 6956 10140 6984
rect 9861 6947 9919 6953
rect 10134 6944 10140 6956
rect 10192 6944 10198 6996
rect 10502 6984 10508 6996
rect 10463 6956 10508 6984
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 1995 6888 2360 6916
rect 2593 6919 2651 6925
rect 1995 6885 2007 6888
rect 1949 6879 2007 6885
rect 2593 6885 2605 6919
rect 2639 6916 2651 6919
rect 3510 6916 3516 6928
rect 2639 6888 3516 6916
rect 2639 6885 2651 6888
rect 2593 6879 2651 6885
rect 3510 6876 3516 6888
rect 3568 6876 3574 6928
rect 5442 6916 5448 6928
rect 5403 6888 5448 6916
rect 5442 6876 5448 6888
rect 5500 6876 5506 6928
rect 6086 6876 6092 6928
rect 6144 6916 6150 6928
rect 6365 6919 6423 6925
rect 6365 6916 6377 6919
rect 6144 6888 6377 6916
rect 6144 6876 6150 6888
rect 6365 6885 6377 6888
rect 6411 6916 6423 6919
rect 9508 6916 9536 6944
rect 6411 6888 9536 6916
rect 6411 6885 6423 6888
rect 6365 6879 6423 6885
rect 1448 6851 1506 6857
rect 1448 6817 1460 6851
rect 1494 6848 1506 6851
rect 2222 6848 2228 6860
rect 1494 6820 2228 6848
rect 1494 6817 1506 6820
rect 1448 6811 1506 6817
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 4062 6848 4068 6860
rect 3927 6820 4068 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 7377 6851 7435 6857
rect 7377 6817 7389 6851
rect 7423 6848 7435 6851
rect 7466 6848 7472 6860
rect 7423 6820 7472 6848
rect 7423 6817 7435 6820
rect 7377 6811 7435 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7742 6848 7748 6860
rect 7703 6820 7748 6848
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 8294 6848 8300 6860
rect 8251 6820 8300 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 8294 6808 8300 6820
rect 8352 6808 8358 6860
rect 9677 6851 9735 6857
rect 9677 6817 9689 6851
rect 9723 6848 9735 6851
rect 10134 6848 10140 6860
rect 9723 6820 10140 6848
rect 9723 6817 9735 6820
rect 9677 6811 9735 6817
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6780 2559 6783
rect 2774 6780 2780 6792
rect 2547 6752 2636 6780
rect 2735 6752 2780 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2608 6712 2636 6752
rect 2774 6740 2780 6752
rect 2832 6740 2838 6792
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 5810 6780 5816 6792
rect 5399 6752 5816 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 3326 6712 3332 6724
rect 2608 6684 3332 6712
rect 3326 6672 3332 6684
rect 3384 6712 3390 6724
rect 3421 6715 3479 6721
rect 3421 6712 3433 6715
rect 3384 6684 3433 6712
rect 3384 6672 3390 6684
rect 3421 6681 3433 6684
rect 3467 6681 3479 6715
rect 3421 6675 3479 6681
rect 4430 6672 4436 6724
rect 4488 6712 4494 6724
rect 5905 6715 5963 6721
rect 5905 6712 5917 6715
rect 4488 6684 5917 6712
rect 4488 6672 4494 6684
rect 5905 6681 5917 6684
rect 5951 6712 5963 6715
rect 7282 6712 7288 6724
rect 5951 6684 7288 6712
rect 5951 6681 5963 6684
rect 5905 6675 5963 6681
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 7561 6715 7619 6721
rect 7561 6681 7573 6715
rect 7607 6712 7619 6715
rect 8202 6712 8208 6724
rect 7607 6684 8208 6712
rect 7607 6681 7619 6684
rect 7561 6675 7619 6681
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 2406 6604 2412 6656
rect 2464 6644 2470 6656
rect 4246 6644 4252 6656
rect 2464 6616 4252 6644
rect 2464 6604 2470 6616
rect 4246 6604 4252 6616
rect 4304 6644 4310 6656
rect 4617 6647 4675 6653
rect 4617 6644 4629 6647
rect 4304 6616 4629 6644
rect 4304 6604 4310 6616
rect 4617 6613 4629 6616
rect 4663 6644 4675 6647
rect 5074 6644 5080 6656
rect 4663 6616 5080 6644
rect 4663 6613 4675 6616
rect 4617 6607 4675 6613
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 9033 6647 9091 6653
rect 9033 6644 9045 6647
rect 8812 6616 9045 6644
rect 8812 6604 8818 6616
rect 9033 6613 9045 6616
rect 9079 6613 9091 6647
rect 9033 6607 9091 6613
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 2498 6440 2504 6452
rect 2459 6412 2504 6440
rect 2498 6400 2504 6412
rect 2556 6440 2562 6452
rect 3234 6440 3240 6452
rect 2556 6412 3240 6440
rect 2556 6400 2562 6412
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 3418 6400 3424 6452
rect 3476 6440 3482 6452
rect 4062 6440 4068 6452
rect 3476 6412 4068 6440
rect 3476 6400 3482 6412
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 5442 6400 5448 6452
rect 5500 6440 5506 6452
rect 5537 6443 5595 6449
rect 5537 6440 5549 6443
rect 5500 6412 5549 6440
rect 5500 6400 5506 6412
rect 5537 6409 5549 6412
rect 5583 6409 5595 6443
rect 5537 6403 5595 6409
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 10962 6440 10968 6452
rect 5684 6412 10968 6440
rect 5684 6400 5690 6412
rect 10962 6400 10968 6412
rect 11020 6440 11026 6452
rect 13722 6440 13728 6452
rect 11020 6412 13728 6440
rect 11020 6400 11026 6412
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 2774 6332 2780 6384
rect 2832 6372 2838 6384
rect 3605 6375 3663 6381
rect 3605 6372 3617 6375
rect 2832 6344 3617 6372
rect 2832 6332 2838 6344
rect 3605 6341 3617 6344
rect 3651 6341 3663 6375
rect 3605 6335 3663 6341
rect 4433 6375 4491 6381
rect 4433 6341 4445 6375
rect 4479 6372 4491 6375
rect 4706 6372 4712 6384
rect 4479 6344 4712 6372
rect 4479 6341 4491 6344
rect 4433 6335 4491 6341
rect 1946 6304 1952 6316
rect 1907 6276 1952 6304
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 3418 6304 3424 6316
rect 3099 6276 3424 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 3620 6304 3648 6335
rect 4706 6332 4712 6344
rect 4764 6372 4770 6384
rect 6914 6372 6920 6384
rect 4764 6344 6920 6372
rect 4764 6332 4770 6344
rect 6914 6332 6920 6344
rect 6972 6372 6978 6384
rect 10042 6372 10048 6384
rect 6972 6344 10048 6372
rect 6972 6332 6978 6344
rect 10042 6332 10048 6344
rect 10100 6332 10106 6384
rect 3881 6307 3939 6313
rect 3620 6276 3740 6304
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 1762 6236 1768 6248
rect 1719 6208 1768 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 2498 6236 2504 6248
rect 1903 6208 2504 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 2498 6196 2504 6208
rect 2556 6196 2562 6248
rect 3142 6128 3148 6180
rect 3200 6168 3206 6180
rect 3712 6168 3740 6276
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 3927 6276 4844 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 4706 6236 4712 6248
rect 4667 6208 4712 6236
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 4816 6236 4844 6276
rect 8036 6276 9444 6304
rect 4985 6239 5043 6245
rect 4985 6236 4997 6239
rect 4816 6208 4997 6236
rect 4985 6205 4997 6208
rect 5031 6205 5043 6239
rect 4985 6199 5043 6205
rect 8036 6168 8064 6276
rect 8113 6239 8171 6245
rect 8113 6205 8125 6239
rect 8159 6236 8171 6239
rect 8386 6236 8392 6248
rect 8159 6208 8392 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 9033 6239 9091 6245
rect 9033 6236 9045 6239
rect 8812 6208 9045 6236
rect 8812 6196 8818 6208
rect 9033 6205 9045 6208
rect 9079 6205 9091 6239
rect 9033 6199 9091 6205
rect 9122 6196 9128 6248
rect 9180 6236 9186 6248
rect 9309 6239 9367 6245
rect 9180 6208 9225 6236
rect 9180 6196 9186 6208
rect 9309 6205 9321 6239
rect 9355 6205 9367 6239
rect 9416 6236 9444 6276
rect 9490 6264 9496 6316
rect 9548 6304 9554 6316
rect 10735 6307 10793 6313
rect 10735 6304 10747 6307
rect 9548 6276 10747 6304
rect 9548 6264 9554 6276
rect 10735 6273 10747 6276
rect 10781 6273 10793 6307
rect 10735 6267 10793 6273
rect 10632 6239 10690 6245
rect 10632 6236 10644 6239
rect 9416 6208 10644 6236
rect 9309 6199 9367 6205
rect 10632 6205 10644 6208
rect 10678 6236 10690 6239
rect 11057 6239 11115 6245
rect 11057 6236 11069 6239
rect 10678 6208 11069 6236
rect 10678 6205 10690 6208
rect 10632 6199 10690 6205
rect 11057 6205 11069 6208
rect 11103 6205 11115 6239
rect 11057 6199 11115 6205
rect 8202 6168 8208 6180
rect 3200 6140 3245 6168
rect 3712 6140 8064 6168
rect 8115 6140 8208 6168
rect 3200 6128 3206 6140
rect 8202 6128 8208 6140
rect 8260 6168 8266 6180
rect 8481 6171 8539 6177
rect 8481 6168 8493 6171
rect 8260 6140 8493 6168
rect 8260 6128 8266 6140
rect 8481 6137 8493 6140
rect 8527 6137 8539 6171
rect 8846 6168 8852 6180
rect 8759 6140 8852 6168
rect 8481 6131 8539 6137
rect 8846 6128 8852 6140
rect 8904 6168 8910 6180
rect 9324 6168 9352 6199
rect 9950 6168 9956 6180
rect 8904 6140 9956 6168
rect 8904 6128 8910 6140
rect 9950 6128 9956 6140
rect 10008 6128 10014 6180
rect 2869 6103 2927 6109
rect 2869 6069 2881 6103
rect 2915 6100 2927 6103
rect 3160 6100 3188 6128
rect 2915 6072 3188 6100
rect 2915 6069 2927 6072
rect 2869 6063 2927 6069
rect 3234 6060 3240 6112
rect 3292 6100 3298 6112
rect 3881 6103 3939 6109
rect 3881 6100 3893 6103
rect 3292 6072 3893 6100
rect 3292 6060 3298 6072
rect 3881 6069 3893 6072
rect 3927 6100 3939 6103
rect 3973 6103 4031 6109
rect 3973 6100 3985 6103
rect 3927 6072 3985 6100
rect 3927 6069 3939 6072
rect 3881 6063 3939 6069
rect 3973 6069 3985 6072
rect 4019 6069 4031 6103
rect 3973 6063 4031 6069
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 4617 6103 4675 6109
rect 4617 6100 4629 6103
rect 4580 6072 4629 6100
rect 4580 6060 4586 6072
rect 4617 6069 4629 6072
rect 4663 6069 4675 6103
rect 5902 6100 5908 6112
rect 5863 6072 5908 6100
rect 4617 6063 4675 6069
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 6638 6100 6644 6112
rect 6599 6072 6644 6100
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 7377 6103 7435 6109
rect 7377 6069 7389 6103
rect 7423 6100 7435 6103
rect 7742 6100 7748 6112
rect 7423 6072 7748 6100
rect 7423 6069 7435 6072
rect 7377 6063 7435 6069
rect 7742 6060 7748 6072
rect 7800 6100 7806 6112
rect 7926 6100 7932 6112
rect 7800 6072 7932 6100
rect 7800 6060 7806 6072
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 8938 6060 8944 6112
rect 8996 6100 9002 6112
rect 9493 6103 9551 6109
rect 9493 6100 9505 6103
rect 8996 6072 9505 6100
rect 8996 6060 9002 6072
rect 9493 6069 9505 6072
rect 9539 6069 9551 6103
rect 10134 6100 10140 6112
rect 10095 6072 10140 6100
rect 9493 6063 9551 6069
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 1765 5899 1823 5905
rect 1765 5865 1777 5899
rect 1811 5896 1823 5899
rect 1854 5896 1860 5908
rect 1811 5868 1860 5896
rect 1811 5865 1823 5868
rect 1765 5859 1823 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 2314 5896 2320 5908
rect 2275 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 3145 5899 3203 5905
rect 3145 5865 3157 5899
rect 3191 5896 3203 5899
rect 3510 5896 3516 5908
rect 3191 5868 3516 5896
rect 3191 5865 3203 5868
rect 3145 5859 3203 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 6086 5856 6092 5908
rect 6144 5896 6150 5908
rect 6273 5899 6331 5905
rect 6273 5896 6285 5899
rect 6144 5868 6285 5896
rect 6144 5856 6150 5868
rect 6273 5865 6285 5868
rect 6319 5865 6331 5899
rect 6273 5859 6331 5865
rect 7558 5856 7564 5908
rect 7616 5896 7622 5908
rect 7745 5899 7803 5905
rect 7745 5896 7757 5899
rect 7616 5868 7757 5896
rect 7616 5856 7622 5868
rect 7745 5865 7757 5868
rect 7791 5865 7803 5899
rect 10134 5896 10140 5908
rect 10095 5868 10140 5896
rect 7745 5859 7803 5865
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 2222 5788 2228 5840
rect 2280 5828 2286 5840
rect 3789 5831 3847 5837
rect 3789 5828 3801 5831
rect 2280 5800 3801 5828
rect 2280 5788 2286 5800
rect 3789 5797 3801 5800
rect 3835 5797 3847 5831
rect 8938 5828 8944 5840
rect 3789 5791 3847 5797
rect 6104 5800 8944 5828
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5729 2375 5763
rect 2498 5760 2504 5772
rect 2459 5732 2504 5760
rect 2317 5723 2375 5729
rect 2332 5692 2360 5723
rect 2498 5720 2504 5732
rect 2556 5720 2562 5772
rect 2774 5692 2780 5704
rect 2332 5664 2780 5692
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 3804 5692 3832 5791
rect 6104 5772 6132 5800
rect 8938 5788 8944 5800
rect 8996 5788 9002 5840
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 4065 5763 4123 5769
rect 4065 5760 4077 5763
rect 4028 5732 4077 5760
rect 4028 5720 4034 5732
rect 4065 5729 4077 5732
rect 4111 5760 4123 5763
rect 4246 5760 4252 5772
rect 4111 5732 4252 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4246 5720 4252 5732
rect 4304 5720 4310 5772
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5760 4675 5763
rect 6086 5760 6092 5772
rect 4663 5732 5212 5760
rect 5999 5732 6092 5760
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 4430 5692 4436 5704
rect 3804 5664 4436 5692
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 4706 5692 4712 5704
rect 4667 5664 4712 5692
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 2866 5584 2872 5636
rect 2924 5624 2930 5636
rect 4982 5624 4988 5636
rect 2924 5596 4988 5624
rect 2924 5584 2930 5596
rect 4982 5584 4988 5596
rect 5040 5584 5046 5636
rect 3418 5556 3424 5568
rect 3379 5528 3424 5556
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 5184 5565 5212 5732
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 6270 5720 6276 5772
rect 6328 5760 6334 5772
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 6328 5732 7113 5760
rect 6328 5720 6334 5732
rect 7101 5729 7113 5732
rect 7147 5760 7159 5763
rect 7190 5760 7196 5772
rect 7147 5732 7196 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 7392 5732 8401 5760
rect 7392 5692 7420 5732
rect 8389 5729 8401 5732
rect 8435 5760 8447 5763
rect 8662 5760 8668 5772
rect 8435 5732 8668 5760
rect 8435 5729 8447 5732
rect 8389 5723 8447 5729
rect 8662 5720 8668 5732
rect 8720 5720 8726 5772
rect 9398 5720 9404 5772
rect 9456 5760 9462 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9456 5732 9689 5760
rect 9456 5720 9462 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9950 5760 9956 5772
rect 9911 5732 9956 5760
rect 9677 5723 9735 5729
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 7116 5664 7420 5692
rect 7469 5695 7527 5701
rect 7116 5568 7144 5664
rect 7469 5661 7481 5695
rect 7515 5692 7527 5695
rect 7926 5692 7932 5704
rect 7515 5664 7932 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 7377 5627 7435 5633
rect 7377 5593 7389 5627
rect 7423 5624 7435 5627
rect 7742 5624 7748 5636
rect 7423 5596 7748 5624
rect 7423 5593 7435 5596
rect 7377 5587 7435 5593
rect 7742 5584 7748 5596
rect 7800 5624 7806 5636
rect 8202 5624 8208 5636
rect 7800 5596 8208 5624
rect 7800 5584 7806 5596
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 8478 5584 8484 5636
rect 8536 5624 8542 5636
rect 9122 5624 9128 5636
rect 8536 5596 9128 5624
rect 8536 5584 8542 5596
rect 9122 5584 9128 5596
rect 9180 5624 9186 5636
rect 9769 5627 9827 5633
rect 9769 5624 9781 5627
rect 9180 5596 9781 5624
rect 9180 5584 9186 5596
rect 9769 5593 9781 5596
rect 9815 5624 9827 5627
rect 10134 5624 10140 5636
rect 9815 5596 10140 5624
rect 9815 5593 9827 5596
rect 9769 5587 9827 5593
rect 10134 5584 10140 5596
rect 10192 5584 10198 5636
rect 5169 5559 5227 5565
rect 5169 5525 5181 5559
rect 5215 5556 5227 5559
rect 5350 5556 5356 5568
rect 5215 5528 5356 5556
rect 5215 5525 5227 5528
rect 5169 5519 5227 5525
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 6917 5559 6975 5565
rect 6917 5525 6929 5559
rect 6963 5556 6975 5559
rect 7098 5556 7104 5568
rect 6963 5528 7104 5556
rect 6963 5525 6975 5528
rect 6917 5519 6975 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7263 5556 7269 5568
rect 7224 5528 7269 5556
rect 7263 5516 7269 5528
rect 7321 5516 7327 5568
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 10226 5556 10232 5568
rect 9364 5528 10232 5556
rect 9364 5516 9370 5528
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 12066 5556 12072 5568
rect 10376 5528 12072 5556
rect 10376 5516 10382 5528
rect 12066 5516 12072 5528
rect 12124 5516 12130 5568
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 1854 5312 1860 5364
rect 1912 5352 1918 5364
rect 3970 5352 3976 5364
rect 1912 5324 3976 5352
rect 1912 5312 1918 5324
rect 3970 5312 3976 5324
rect 4028 5312 4034 5364
rect 4246 5352 4252 5364
rect 4207 5324 4252 5352
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 6270 5352 6276 5364
rect 6231 5324 6276 5352
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 9306 5312 9312 5364
rect 9364 5352 9370 5364
rect 9401 5355 9459 5361
rect 9401 5352 9413 5355
rect 9364 5324 9413 5352
rect 9364 5312 9370 5324
rect 9401 5321 9413 5324
rect 9447 5321 9459 5355
rect 9766 5352 9772 5364
rect 9727 5324 9772 5352
rect 9401 5315 9459 5321
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 10965 5355 11023 5361
rect 10965 5352 10977 5355
rect 10008 5324 10977 5352
rect 10008 5312 10014 5324
rect 10965 5321 10977 5324
rect 11011 5321 11023 5355
rect 10965 5315 11023 5321
rect 2774 5284 2780 5296
rect 2687 5256 2780 5284
rect 2774 5244 2780 5256
rect 2832 5284 2838 5296
rect 4617 5287 4675 5293
rect 4617 5284 4629 5287
rect 2832 5256 4629 5284
rect 2832 5244 2838 5256
rect 4617 5253 4629 5256
rect 4663 5253 4675 5287
rect 6638 5284 6644 5296
rect 6551 5256 6644 5284
rect 4617 5247 4675 5253
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 3605 5219 3663 5225
rect 3605 5216 3617 5219
rect 3384 5188 3617 5216
rect 3384 5176 3390 5188
rect 3605 5185 3617 5188
rect 3651 5216 3663 5219
rect 3651 5188 4154 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 1854 5148 1860 5160
rect 1815 5120 1860 5148
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 2225 5151 2283 5157
rect 2225 5117 2237 5151
rect 2271 5148 2283 5151
rect 2498 5148 2504 5160
rect 2271 5120 2504 5148
rect 2271 5117 2283 5120
rect 2225 5111 2283 5117
rect 2498 5108 2504 5120
rect 2556 5108 2562 5160
rect 2406 5080 2412 5092
rect 2367 5052 2412 5080
rect 2406 5040 2412 5052
rect 2464 5040 2470 5092
rect 3326 5080 3332 5092
rect 3287 5052 3332 5080
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 3421 5083 3479 5089
rect 3421 5049 3433 5083
rect 3467 5049 3479 5083
rect 4126 5080 4154 5188
rect 4632 5148 4660 5247
rect 6638 5244 6644 5256
rect 6696 5284 6702 5296
rect 6917 5287 6975 5293
rect 6917 5284 6929 5287
rect 6696 5256 6929 5284
rect 6696 5244 6702 5256
rect 6917 5253 6929 5256
rect 6963 5284 6975 5287
rect 8297 5287 8355 5293
rect 8297 5284 8309 5287
rect 6963 5256 8309 5284
rect 6963 5253 6975 5256
rect 6917 5247 6975 5253
rect 8297 5253 8309 5256
rect 8343 5284 8355 5287
rect 8478 5284 8484 5296
rect 8343 5256 8484 5284
rect 8343 5253 8355 5256
rect 8297 5247 8355 5253
rect 8478 5244 8484 5256
rect 8536 5244 8542 5296
rect 9784 5284 9812 5312
rect 10045 5287 10103 5293
rect 10045 5284 10057 5287
rect 9784 5256 10057 5284
rect 10045 5253 10057 5256
rect 10091 5253 10103 5287
rect 10045 5247 10103 5253
rect 10134 5244 10140 5296
rect 10192 5284 10198 5296
rect 11333 5287 11391 5293
rect 11333 5284 11345 5287
rect 10192 5256 11345 5284
rect 10192 5244 10198 5256
rect 11333 5253 11345 5256
rect 11379 5253 11391 5287
rect 11333 5247 11391 5253
rect 7282 5216 7288 5228
rect 6840 5188 7288 5216
rect 4801 5151 4859 5157
rect 4801 5148 4813 5151
rect 4632 5120 4813 5148
rect 4801 5117 4813 5120
rect 4847 5117 4859 5151
rect 5350 5148 5356 5160
rect 5311 5120 5356 5148
rect 4801 5111 4859 5117
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5148 5963 5151
rect 6638 5148 6644 5160
rect 5951 5120 6644 5148
rect 5951 5117 5963 5120
rect 5905 5111 5963 5117
rect 6638 5108 6644 5120
rect 6696 5148 6702 5160
rect 6840 5157 6868 5188
rect 7282 5176 7288 5188
rect 7340 5216 7346 5228
rect 7340 5188 8800 5216
rect 7340 5176 7346 5188
rect 8772 5160 8800 5188
rect 9398 5176 9404 5228
rect 9456 5216 9462 5228
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 9456 5188 10425 5216
rect 9456 5176 9462 5188
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 10413 5179 10471 5185
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6696 5120 6837 5148
rect 6696 5108 6702 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 7098 5148 7104 5160
rect 7059 5120 7104 5148
rect 6825 5111 6883 5117
rect 7098 5108 7104 5120
rect 7156 5108 7162 5160
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 8386 5148 8392 5160
rect 7524 5120 8392 5148
rect 7524 5108 7530 5120
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 8662 5148 8668 5160
rect 8623 5120 8668 5148
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 8754 5108 8760 5160
rect 8812 5148 8818 5160
rect 9950 5148 9956 5160
rect 8812 5120 9956 5148
rect 8812 5108 8818 5120
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 10226 5148 10232 5160
rect 10187 5120 10232 5148
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 7650 5080 7656 5092
rect 4126 5052 7656 5080
rect 3421 5043 3479 5049
rect 2958 4972 2964 5024
rect 3016 5012 3022 5024
rect 3053 5015 3111 5021
rect 3053 5012 3065 5015
rect 3016 4984 3065 5012
rect 3016 4972 3022 4984
rect 3053 4981 3065 4984
rect 3099 5012 3111 5015
rect 3436 5012 3464 5043
rect 7650 5040 7656 5052
rect 7708 5040 7714 5092
rect 9125 5083 9183 5089
rect 9125 5049 9137 5083
rect 9171 5080 9183 5083
rect 11054 5080 11060 5092
rect 9171 5052 11060 5080
rect 9171 5049 9183 5052
rect 9125 5043 9183 5049
rect 11054 5040 11060 5052
rect 11112 5040 11118 5092
rect 3099 4984 3464 5012
rect 3099 4981 3111 4984
rect 3053 4975 3111 4981
rect 4338 4972 4344 5024
rect 4396 5012 4402 5024
rect 4614 5012 4620 5024
rect 4396 4984 4620 5012
rect 4396 4972 4402 4984
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 4890 5012 4896 5024
rect 4851 4984 4896 5012
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 7285 5015 7343 5021
rect 7285 5012 7297 5015
rect 6052 4984 7297 5012
rect 6052 4972 6058 4984
rect 7285 4981 7297 4984
rect 7331 4981 7343 5015
rect 7926 5012 7932 5024
rect 7887 4984 7932 5012
rect 7285 4975 7343 4981
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 9306 5012 9312 5024
rect 8536 4984 9312 5012
rect 8536 4972 8542 4984
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2317 4811 2375 4817
rect 2317 4808 2329 4811
rect 1995 4780 2329 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2317 4777 2329 4780
rect 2363 4808 2375 4811
rect 2498 4808 2504 4820
rect 2363 4780 2504 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 4706 4808 4712 4820
rect 4667 4780 4712 4808
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 5718 4808 5724 4820
rect 4816 4780 5724 4808
rect 2590 4740 2596 4752
rect 2551 4712 2596 4740
rect 2590 4700 2596 4712
rect 2648 4700 2654 4752
rect 3142 4700 3148 4752
rect 3200 4740 3206 4752
rect 4816 4740 4844 4780
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 6086 4808 6092 4820
rect 6047 4780 6092 4808
rect 6086 4768 6092 4780
rect 6144 4768 6150 4820
rect 7742 4808 7748 4820
rect 6564 4780 7512 4808
rect 7703 4780 7748 4808
rect 3200 4712 4844 4740
rect 3200 4700 3206 4712
rect 5074 4700 5080 4752
rect 5132 4740 5138 4752
rect 5214 4743 5272 4749
rect 5214 4740 5226 4743
rect 5132 4712 5226 4740
rect 5132 4700 5138 4712
rect 5214 4709 5226 4712
rect 5260 4709 5272 4743
rect 5214 4703 5272 4709
rect 1464 4675 1522 4681
rect 1464 4641 1476 4675
rect 1510 4672 1522 4675
rect 1670 4672 1676 4684
rect 1510 4644 1676 4672
rect 1510 4641 1522 4644
rect 1464 4635 1522 4641
rect 1670 4632 1676 4644
rect 1728 4632 1734 4684
rect 4893 4675 4951 4681
rect 4893 4641 4905 4675
rect 4939 4672 4951 4675
rect 5718 4672 5724 4684
rect 4939 4644 5724 4672
rect 4939 4641 4951 4644
rect 4893 4635 4951 4641
rect 5718 4632 5724 4644
rect 5776 4672 5782 4684
rect 6564 4672 6592 4780
rect 6822 4740 6828 4752
rect 6783 4712 6828 4740
rect 6822 4700 6828 4712
rect 6880 4700 6886 4752
rect 7374 4740 7380 4752
rect 7335 4712 7380 4740
rect 7374 4700 7380 4712
rect 7432 4700 7438 4752
rect 7484 4740 7512 4780
rect 7742 4768 7748 4780
rect 7800 4768 7806 4820
rect 9769 4811 9827 4817
rect 9769 4808 9781 4811
rect 7852 4780 9781 4808
rect 7852 4740 7880 4780
rect 9769 4777 9781 4780
rect 9815 4777 9827 4811
rect 9769 4771 9827 4777
rect 7484 4712 7880 4740
rect 8018 4700 8024 4752
rect 8076 4740 8082 4752
rect 8076 4712 8248 4740
rect 8076 4700 8082 4712
rect 8220 4681 8248 4712
rect 8386 4700 8392 4752
rect 8444 4740 8450 4752
rect 8757 4743 8815 4749
rect 8757 4740 8769 4743
rect 8444 4712 8769 4740
rect 8444 4700 8450 4712
rect 8757 4709 8769 4712
rect 8803 4740 8815 4743
rect 9398 4740 9404 4752
rect 8803 4712 9404 4740
rect 8803 4709 8815 4712
rect 8757 4703 8815 4709
rect 9398 4700 9404 4712
rect 9456 4700 9462 4752
rect 5776 4644 6592 4672
rect 8205 4675 8263 4681
rect 5776 4632 5782 4644
rect 8205 4641 8217 4675
rect 8251 4641 8263 4675
rect 8205 4635 8263 4641
rect 9953 4675 10011 4681
rect 9953 4641 9965 4675
rect 9999 4672 10011 4675
rect 10042 4672 10048 4684
rect 9999 4644 10048 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10226 4672 10232 4684
rect 10187 4644 10232 4672
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 11238 4672 11244 4684
rect 11199 4644 11244 4672
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 2038 4564 2044 4616
rect 2096 4604 2102 4616
rect 2501 4607 2559 4613
rect 2501 4604 2513 4607
rect 2096 4576 2513 4604
rect 2096 4564 2102 4576
rect 2501 4573 2513 4576
rect 2547 4573 2559 4607
rect 2501 4567 2559 4573
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4604 3203 4607
rect 3234 4604 3240 4616
rect 3191 4576 3240 4604
rect 3191 4573 3203 4576
rect 3145 4567 3203 4573
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 5350 4604 5356 4616
rect 4387 4576 5356 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 6733 4607 6791 4613
rect 6733 4573 6745 4607
rect 6779 4604 6791 4607
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 6779 4576 8033 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 8021 4573 8033 4576
rect 8067 4604 8079 4607
rect 8110 4604 8116 4616
rect 8067 4576 8116 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 4798 4496 4804 4548
rect 4856 4536 4862 4548
rect 7558 4536 7564 4548
rect 4856 4508 7564 4536
rect 4856 4496 4862 4508
rect 7558 4496 7564 4508
rect 7616 4496 7622 4548
rect 1535 4471 1593 4477
rect 1535 4437 1547 4471
rect 1581 4468 1593 4471
rect 1762 4468 1768 4480
rect 1581 4440 1768 4468
rect 1581 4437 1593 4440
rect 1535 4431 1593 4437
rect 1762 4428 1768 4440
rect 1820 4428 1826 4480
rect 3326 4428 3332 4480
rect 3384 4468 3390 4480
rect 3513 4471 3571 4477
rect 3513 4468 3525 4471
rect 3384 4440 3525 4468
rect 3384 4428 3390 4440
rect 3513 4437 3525 4440
rect 3559 4468 3571 4471
rect 3970 4468 3976 4480
rect 3559 4440 3976 4468
rect 3559 4437 3571 4440
rect 3513 4431 3571 4437
rect 3970 4428 3976 4440
rect 4028 4428 4034 4480
rect 5810 4468 5816 4480
rect 5771 4440 5816 4468
rect 5810 4428 5816 4440
rect 5868 4428 5874 4480
rect 6549 4471 6607 4477
rect 6549 4437 6561 4471
rect 6595 4468 6607 4471
rect 6638 4468 6644 4480
rect 6595 4440 6644 4468
rect 6595 4437 6607 4440
rect 6549 4431 6607 4437
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 8386 4468 8392 4480
rect 8347 4440 8392 4468
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 10689 4471 10747 4477
rect 10689 4468 10701 4471
rect 10008 4440 10701 4468
rect 10008 4428 10014 4440
rect 10689 4437 10701 4440
rect 10735 4437 10747 4471
rect 10689 4431 10747 4437
rect 10778 4428 10784 4480
rect 10836 4468 10842 4480
rect 11379 4471 11437 4477
rect 11379 4468 11391 4471
rect 10836 4440 11391 4468
rect 10836 4428 10842 4440
rect 11379 4437 11391 4440
rect 11425 4437 11437 4471
rect 11379 4431 11437 4437
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 6181 4267 6239 4273
rect 6181 4264 6193 4267
rect 5868 4236 6193 4264
rect 5868 4224 5874 4236
rect 6181 4233 6193 4236
rect 6227 4264 6239 4267
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6227 4236 6561 4264
rect 6227 4233 6239 4236
rect 6181 4227 6239 4233
rect 6549 4233 6561 4236
rect 6595 4264 6607 4267
rect 6822 4264 6828 4276
rect 6595 4236 6828 4264
rect 6595 4233 6607 4236
rect 6549 4227 6607 4233
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 7837 4267 7895 4273
rect 7837 4233 7849 4267
rect 7883 4264 7895 4267
rect 8018 4264 8024 4276
rect 7883 4236 8024 4264
rect 7883 4233 7895 4236
rect 7837 4227 7895 4233
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 8662 4264 8668 4276
rect 8623 4236 8668 4264
rect 8662 4224 8668 4236
rect 8720 4224 8726 4276
rect 9769 4267 9827 4273
rect 9769 4233 9781 4267
rect 9815 4264 9827 4267
rect 10042 4264 10048 4276
rect 9815 4236 10048 4264
rect 9815 4233 9827 4236
rect 9769 4227 9827 4233
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 10137 4267 10195 4273
rect 10137 4233 10149 4267
rect 10183 4264 10195 4267
rect 11330 4264 11336 4276
rect 10183 4236 11336 4264
rect 10183 4233 10195 4236
rect 10137 4227 10195 4233
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 1903 4199 1961 4205
rect 1903 4165 1915 4199
rect 1949 4196 1961 4199
rect 7558 4196 7564 4208
rect 1949 4168 7564 4196
rect 1949 4165 1961 4168
rect 1903 4159 1961 4165
rect 7558 4156 7564 4168
rect 7616 4156 7622 4208
rect 7926 4156 7932 4208
rect 7984 4196 7990 4208
rect 8846 4196 8852 4208
rect 7984 4168 8852 4196
rect 7984 4156 7990 4168
rect 8846 4156 8852 4168
rect 8904 4156 8910 4208
rect 10597 4199 10655 4205
rect 10597 4196 10609 4199
rect 10060 4168 10609 4196
rect 1670 4128 1676 4140
rect 1631 4100 1676 4128
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 3326 4128 3332 4140
rect 3287 4100 3332 4128
rect 3326 4088 3332 4100
rect 3384 4088 3390 4140
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4128 4491 4131
rect 4614 4128 4620 4140
rect 4479 4100 4620 4128
rect 4479 4097 4491 4100
rect 4433 4091 4491 4097
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 6917 4131 6975 4137
rect 6917 4097 6929 4131
rect 6963 4128 6975 4131
rect 7006 4128 7012 4140
rect 6963 4100 7012 4128
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7098 4088 7104 4140
rect 7156 4128 7162 4140
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 7156 4100 7205 4128
rect 7156 4088 7162 4100
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 1832 4063 1890 4069
rect 1832 4029 1844 4063
rect 1878 4060 1890 4063
rect 8297 4063 8355 4069
rect 1878 4032 2360 4060
rect 1878 4029 1890 4032
rect 1832 4023 1890 4029
rect 2332 4001 2360 4032
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8754 4060 8760 4072
rect 8343 4032 8760 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8754 4020 8760 4032
rect 8812 4060 8818 4072
rect 8864 4060 8892 4156
rect 8812 4032 8892 4060
rect 9953 4063 10011 4069
rect 8812 4020 8818 4032
rect 9953 4029 9965 4063
rect 9999 4060 10011 4063
rect 10060 4060 10088 4168
rect 10597 4165 10609 4168
rect 10643 4196 10655 4199
rect 12158 4196 12164 4208
rect 10643 4168 12164 4196
rect 10643 4165 10655 4168
rect 10597 4159 10655 4165
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 9999 4032 10088 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 10410 4020 10416 4072
rect 10468 4060 10474 4072
rect 11146 4069 11152 4072
rect 11092 4063 11152 4069
rect 11092 4060 11104 4063
rect 10468 4032 11104 4060
rect 10468 4020 10474 4032
rect 11092 4029 11104 4032
rect 11138 4029 11152 4063
rect 11092 4023 11152 4029
rect 11146 4020 11152 4023
rect 11204 4020 11210 4072
rect 11238 4020 11244 4072
rect 11296 4020 11302 4072
rect 11422 4020 11428 4072
rect 11480 4060 11486 4072
rect 12472 4063 12530 4069
rect 12472 4060 12484 4063
rect 11480 4032 12484 4060
rect 11480 4020 11486 4032
rect 12472 4029 12484 4032
rect 12518 4060 12530 4063
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12518 4032 12909 4060
rect 12518 4029 12530 4032
rect 12472 4023 12530 4029
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 2317 3995 2375 4001
rect 2317 3961 2329 3995
rect 2363 3992 2375 3995
rect 2682 3992 2688 4004
rect 2363 3964 2688 3992
rect 2363 3961 2375 3964
rect 2317 3955 2375 3961
rect 2682 3952 2688 3964
rect 2740 3952 2746 4004
rect 2869 3995 2927 4001
rect 2869 3961 2881 3995
rect 2915 3961 2927 3995
rect 2869 3955 2927 3961
rect 2590 3924 2596 3936
rect 2551 3896 2596 3924
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2884 3924 2912 3955
rect 2958 3952 2964 4004
rect 3016 3992 3022 4004
rect 4795 3995 4853 4001
rect 3016 3964 3109 3992
rect 3016 3952 3022 3964
rect 4795 3961 4807 3995
rect 4841 3961 4853 3995
rect 5629 3995 5687 4001
rect 5629 3992 5641 3995
rect 4795 3955 4853 3961
rect 5092 3964 5641 3992
rect 2832 3896 2912 3924
rect 2976 3924 3004 3952
rect 3789 3927 3847 3933
rect 3789 3924 3801 3927
rect 2976 3896 3801 3924
rect 2832 3884 2838 3896
rect 3789 3893 3801 3896
rect 3835 3893 3847 3927
rect 3789 3887 3847 3893
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3924 4399 3927
rect 4810 3924 4838 3955
rect 5092 3936 5120 3964
rect 5629 3961 5641 3964
rect 5675 3961 5687 3995
rect 5629 3955 5687 3961
rect 7009 3995 7067 4001
rect 7009 3961 7021 3995
rect 7055 3961 7067 3995
rect 7009 3955 7067 3961
rect 5074 3924 5080 3936
rect 4387 3896 5080 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5350 3924 5356 3936
rect 5311 3896 5356 3924
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 6822 3884 6828 3936
rect 6880 3924 6886 3936
rect 7024 3924 7052 3955
rect 8110 3952 8116 4004
rect 8168 3992 8174 4004
rect 8168 3964 8524 3992
rect 8168 3952 8174 3964
rect 6880 3896 7052 3924
rect 8496 3924 8524 3964
rect 10686 3952 10692 4004
rect 10744 3992 10750 4004
rect 11256 3992 11284 4020
rect 11885 3995 11943 4001
rect 10744 3964 11319 3992
rect 10744 3952 10750 3964
rect 11195 3927 11253 3933
rect 11195 3924 11207 3927
rect 8496 3896 11207 3924
rect 6880 3884 6886 3896
rect 11195 3893 11207 3896
rect 11241 3893 11253 3927
rect 11291 3924 11319 3964
rect 11885 3961 11897 3995
rect 11931 3992 11943 3995
rect 12066 3992 12072 4004
rect 11931 3964 12072 3992
rect 11931 3961 11943 3964
rect 11885 3955 11943 3961
rect 12066 3952 12072 3964
rect 12124 3952 12130 4004
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11291 3896 11529 3924
rect 11195 3887 11253 3893
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12575 3927 12633 3933
rect 12575 3924 12587 3927
rect 12032 3896 12587 3924
rect 12032 3884 12038 3896
rect 12575 3893 12587 3896
rect 12621 3893 12633 3927
rect 12575 3887 12633 3893
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 2498 3720 2504 3732
rect 2459 3692 2504 3720
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 4341 3723 4399 3729
rect 4341 3689 4353 3723
rect 4387 3720 4399 3723
rect 4430 3720 4436 3732
rect 4387 3692 4436 3720
rect 4387 3689 4399 3692
rect 4341 3683 4399 3689
rect 4430 3680 4436 3692
rect 4488 3720 4494 3732
rect 4890 3720 4896 3732
rect 4488 3692 4896 3720
rect 4488 3680 4494 3692
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 5718 3720 5724 3732
rect 5679 3692 5724 3720
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 7558 3720 7564 3732
rect 7519 3692 7564 3720
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 9858 3720 9864 3732
rect 7668 3692 8524 3720
rect 9819 3692 9864 3720
rect 2038 3652 2044 3664
rect 1999 3624 2044 3652
rect 2038 3612 2044 3624
rect 2096 3612 2102 3664
rect 4795 3655 4853 3661
rect 4795 3621 4807 3655
rect 4841 3652 4853 3655
rect 5074 3652 5080 3664
rect 4841 3624 5080 3652
rect 4841 3621 4853 3624
rect 4795 3615 4853 3621
rect 5074 3612 5080 3624
rect 5132 3612 5138 3664
rect 5350 3612 5356 3664
rect 5408 3652 5414 3664
rect 6270 3652 6276 3664
rect 5408 3624 6276 3652
rect 5408 3612 5414 3624
rect 6270 3612 6276 3624
rect 6328 3652 6334 3664
rect 6365 3655 6423 3661
rect 6365 3652 6377 3655
rect 6328 3624 6377 3652
rect 6328 3612 6334 3624
rect 6365 3621 6377 3624
rect 6411 3621 6423 3655
rect 6365 3615 6423 3621
rect 1762 3544 1768 3596
rect 1820 3584 1826 3596
rect 3789 3587 3847 3593
rect 3789 3584 3801 3587
rect 1820 3556 3801 3584
rect 1820 3544 1826 3556
rect 3789 3553 3801 3556
rect 3835 3584 3847 3587
rect 5258 3584 5264 3596
rect 3835 3556 5264 3584
rect 3835 3553 3847 3556
rect 3789 3547 3847 3553
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3516 2191 3519
rect 2406 3516 2412 3528
rect 2179 3488 2412 3516
rect 2179 3485 2191 3488
rect 2133 3479 2191 3485
rect 2406 3476 2412 3488
rect 2464 3516 2470 3528
rect 3510 3516 3516 3528
rect 2464 3488 3516 3516
rect 2464 3476 2470 3488
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 4430 3516 4436 3528
rect 4391 3488 4436 3516
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3516 6147 3519
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 6135 3488 6285 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 6273 3485 6285 3488
rect 6319 3516 6331 3519
rect 7668 3516 7696 3692
rect 7926 3652 7932 3664
rect 7887 3624 7932 3652
rect 7926 3612 7932 3624
rect 7984 3612 7990 3664
rect 8496 3584 8524 3692
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 10229 3723 10287 3729
rect 10229 3689 10241 3723
rect 10275 3720 10287 3723
rect 15746 3720 15752 3732
rect 10275 3692 15752 3720
rect 10275 3689 10287 3692
rect 10229 3683 10287 3689
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 8573 3655 8631 3661
rect 8573 3621 8585 3655
rect 8619 3652 8631 3655
rect 8849 3655 8907 3661
rect 8849 3652 8861 3655
rect 8619 3624 8861 3652
rect 8619 3621 8631 3624
rect 8573 3615 8631 3621
rect 8849 3621 8861 3624
rect 8895 3652 8907 3655
rect 11974 3652 11980 3664
rect 8895 3624 11980 3652
rect 8895 3621 8907 3624
rect 8849 3615 8907 3621
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 10045 3587 10103 3593
rect 8496 3556 9674 3584
rect 6319 3488 7696 3516
rect 7837 3519 7895 3525
rect 6319 3485 6331 3488
rect 6273 3479 6331 3485
rect 7837 3485 7849 3519
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 2774 3408 2780 3460
rect 2832 3448 2838 3460
rect 2832 3420 3464 3448
rect 2832 3408 2838 3420
rect 3436 3392 3464 3420
rect 5902 3408 5908 3460
rect 5960 3448 5966 3460
rect 6825 3451 6883 3457
rect 6825 3448 6837 3451
rect 5960 3420 6837 3448
rect 5960 3408 5966 3420
rect 6825 3417 6837 3420
rect 6871 3448 6883 3451
rect 7098 3448 7104 3460
rect 6871 3420 7104 3448
rect 6871 3417 6883 3420
rect 6825 3411 6883 3417
rect 7098 3408 7104 3420
rect 7156 3408 7162 3460
rect 7742 3408 7748 3460
rect 7800 3448 7806 3460
rect 7852 3448 7880 3479
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 8573 3519 8631 3525
rect 8573 3516 8585 3519
rect 8352 3488 8585 3516
rect 8352 3476 8358 3488
rect 8573 3485 8585 3488
rect 8619 3485 8631 3519
rect 9646 3516 9674 3556
rect 10045 3553 10057 3587
rect 10091 3584 10103 3587
rect 10318 3584 10324 3596
rect 10091 3556 10324 3584
rect 10091 3553 10103 3556
rect 10045 3547 10103 3553
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 11146 3584 11152 3596
rect 11107 3556 11152 3584
rect 11146 3544 11152 3556
rect 11204 3584 11210 3596
rect 12066 3584 12072 3596
rect 11204 3556 12072 3584
rect 11204 3544 11210 3556
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 12158 3544 12164 3596
rect 12216 3584 12222 3596
rect 12288 3587 12346 3593
rect 12288 3584 12300 3587
rect 12216 3556 12300 3584
rect 12216 3544 12222 3556
rect 12288 3553 12300 3556
rect 12334 3553 12346 3587
rect 13262 3584 13268 3596
rect 13223 3556 13268 3584
rect 12288 3547 12346 3553
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 13403 3519 13461 3525
rect 13403 3516 13415 3519
rect 9646 3488 13415 3516
rect 8573 3479 8631 3485
rect 13403 3485 13415 3488
rect 13449 3485 13461 3519
rect 13403 3479 13461 3485
rect 7800 3420 7880 3448
rect 8389 3451 8447 3457
rect 7800 3408 7806 3420
rect 8389 3417 8401 3451
rect 8435 3417 8447 3451
rect 8389 3411 8447 3417
rect 11333 3451 11391 3457
rect 11333 3417 11345 3451
rect 11379 3448 11391 3451
rect 15194 3448 15200 3460
rect 11379 3420 15200 3448
rect 11379 3417 11391 3420
rect 11333 3411 11391 3417
rect 2590 3340 2596 3392
rect 2648 3380 2654 3392
rect 3053 3383 3111 3389
rect 3053 3380 3065 3383
rect 2648 3352 3065 3380
rect 2648 3340 2654 3352
rect 3053 3349 3065 3352
rect 3099 3349 3111 3383
rect 3418 3380 3424 3392
rect 3379 3352 3424 3380
rect 3053 3343 3111 3349
rect 3418 3340 3424 3352
rect 3476 3340 3482 3392
rect 5350 3380 5356 3392
rect 5263 3352 5356 3380
rect 5350 3340 5356 3352
rect 5408 3380 5414 3392
rect 6638 3380 6644 3392
rect 5408 3352 6644 3380
rect 5408 3340 5414 3352
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 7006 3340 7012 3392
rect 7064 3380 7070 3392
rect 7193 3383 7251 3389
rect 7193 3380 7205 3383
rect 7064 3352 7205 3380
rect 7064 3340 7070 3352
rect 7193 3349 7205 3352
rect 7239 3349 7251 3383
rect 7193 3343 7251 3349
rect 7374 3340 7380 3392
rect 7432 3380 7438 3392
rect 8404 3380 8432 3411
rect 15194 3408 15200 3420
rect 15252 3408 15258 3460
rect 7432 3352 8432 3380
rect 7432 3340 7438 3352
rect 9306 3340 9312 3392
rect 9364 3380 9370 3392
rect 12391 3383 12449 3389
rect 12391 3380 12403 3383
rect 9364 3352 12403 3380
rect 9364 3340 9370 3352
rect 12391 3349 12403 3352
rect 12437 3349 12449 3383
rect 12391 3343 12449 3349
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 2958 3136 2964 3188
rect 3016 3176 3022 3188
rect 3237 3179 3295 3185
rect 3237 3176 3249 3179
rect 3016 3148 3249 3176
rect 3016 3136 3022 3148
rect 3237 3145 3249 3148
rect 3283 3145 3295 3179
rect 3510 3176 3516 3188
rect 3471 3148 3516 3176
rect 3237 3139 3295 3145
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 4709 3179 4767 3185
rect 4709 3176 4721 3179
rect 4126 3148 4721 3176
rect 1670 3068 1676 3120
rect 1728 3108 1734 3120
rect 4126 3108 4154 3148
rect 4709 3145 4721 3148
rect 4755 3176 4767 3179
rect 4890 3176 4896 3188
rect 4755 3148 4896 3176
rect 4755 3145 4767 3148
rect 4709 3139 4767 3145
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 6270 3176 6276 3188
rect 6231 3148 6276 3176
rect 6270 3136 6276 3148
rect 6328 3176 6334 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6328 3148 6561 3176
rect 6328 3136 6334 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 1728 3080 4154 3108
rect 1728 3068 1734 3080
rect 2314 3040 2320 3052
rect 2227 3012 2320 3040
rect 2314 3000 2320 3012
rect 2372 3040 2378 3052
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 2372 3012 3893 3040
rect 2372 3000 2378 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 4080 2981 4108 3080
rect 5258 3040 5264 3052
rect 5219 3012 5264 3040
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 5902 3040 5908 3052
rect 5863 3012 5908 3040
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 4065 2975 4123 2981
rect 4065 2941 4077 2975
rect 4111 2941 4123 2975
rect 4065 2935 4123 2941
rect 1857 2907 1915 2913
rect 1857 2873 1869 2907
rect 1903 2904 1915 2907
rect 2225 2907 2283 2913
rect 2225 2904 2237 2907
rect 1903 2876 2237 2904
rect 1903 2873 1915 2876
rect 1857 2867 1915 2873
rect 2225 2873 2237 2876
rect 2271 2904 2283 2907
rect 2498 2904 2504 2916
rect 2271 2876 2504 2904
rect 2271 2873 2283 2876
rect 2225 2867 2283 2873
rect 2498 2864 2504 2876
rect 2556 2904 2562 2916
rect 2679 2907 2737 2913
rect 2679 2904 2691 2907
rect 2556 2876 2691 2904
rect 2556 2864 2562 2876
rect 2679 2873 2691 2876
rect 2725 2873 2737 2907
rect 2679 2867 2737 2873
rect 2694 2836 2722 2867
rect 2774 2864 2780 2916
rect 2832 2904 2838 2916
rect 4338 2904 4344 2916
rect 2832 2876 4344 2904
rect 2832 2864 2838 2876
rect 4338 2864 4344 2876
rect 4396 2864 4402 2916
rect 5350 2904 5356 2916
rect 5311 2876 5356 2904
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 6564 2904 6592 3139
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 7926 3176 7932 3188
rect 6696 3148 7932 3176
rect 6696 3136 6702 3148
rect 7926 3136 7932 3148
rect 7984 3136 7990 3188
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3176 9919 3179
rect 10318 3176 10324 3188
rect 9907 3148 10324 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 10594 3176 10600 3188
rect 10555 3148 10600 3176
rect 10594 3136 10600 3148
rect 10652 3136 10658 3188
rect 11057 3179 11115 3185
rect 11057 3145 11069 3179
rect 11103 3176 11115 3179
rect 11146 3176 11152 3188
rect 11103 3148 11152 3176
rect 11103 3145 11115 3148
rect 11057 3139 11115 3145
rect 11146 3136 11152 3148
rect 11204 3136 11210 3188
rect 12158 3176 12164 3188
rect 12119 3148 12164 3176
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 12250 3136 12256 3188
rect 12308 3176 12314 3188
rect 13587 3179 13645 3185
rect 13587 3176 13599 3179
rect 12308 3148 13599 3176
rect 12308 3136 12314 3148
rect 13587 3145 13599 3148
rect 13633 3145 13645 3179
rect 13587 3139 13645 3145
rect 7374 3068 7380 3120
rect 7432 3108 7438 3120
rect 7469 3111 7527 3117
rect 7469 3108 7481 3111
rect 7432 3080 7481 3108
rect 7432 3068 7438 3080
rect 7469 3077 7481 3080
rect 7515 3077 7527 3111
rect 7469 3071 7527 3077
rect 7650 3068 7656 3120
rect 7708 3108 7714 3120
rect 10137 3111 10195 3117
rect 7708 3080 8800 3108
rect 7708 3068 7714 3080
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3040 6975 3043
rect 7558 3040 7564 3052
rect 6963 3012 7564 3040
rect 6963 3009 6975 3012
rect 6917 3003 6975 3009
rect 7558 3000 7564 3012
rect 7616 3000 7622 3052
rect 8772 3049 8800 3080
rect 10137 3077 10149 3111
rect 10183 3108 10195 3111
rect 10686 3108 10692 3120
rect 10183 3080 10692 3108
rect 10183 3077 10195 3080
rect 10137 3071 10195 3077
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 11333 3111 11391 3117
rect 11333 3077 11345 3111
rect 11379 3108 11391 3111
rect 12434 3108 12440 3120
rect 11379 3080 12440 3108
rect 11379 3077 11391 3080
rect 11333 3071 11391 3077
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 8757 3043 8815 3049
rect 8757 3009 8769 3043
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 10870 3000 10876 3052
rect 10928 3040 10934 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 10928 3012 11713 3040
rect 10928 3000 10934 3012
rect 11164 2984 11192 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 9953 2975 10011 2981
rect 9953 2941 9965 2975
rect 9999 2972 10011 2975
rect 10594 2972 10600 2984
rect 9999 2944 10600 2972
rect 9999 2941 10011 2944
rect 9953 2935 10011 2941
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 11146 2972 11152 2984
rect 11107 2944 11152 2972
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 12472 2975 12530 2981
rect 12472 2972 12484 2975
rect 11572 2944 12484 2972
rect 11572 2932 11578 2944
rect 12472 2941 12484 2944
rect 12518 2972 12530 2975
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 12518 2944 12909 2972
rect 12518 2941 12530 2944
rect 12472 2935 12530 2941
rect 12897 2941 12909 2944
rect 12943 2941 12955 2975
rect 12897 2935 12955 2941
rect 13516 2975 13574 2981
rect 13516 2941 13528 2975
rect 13562 2972 13574 2975
rect 13814 2972 13820 2984
rect 13562 2944 13820 2972
rect 13562 2941 13574 2944
rect 13516 2935 13574 2941
rect 13814 2932 13820 2944
rect 13872 2972 13878 2984
rect 13909 2975 13967 2981
rect 13909 2972 13921 2975
rect 13872 2944 13921 2972
rect 13872 2932 13878 2944
rect 13909 2941 13921 2944
rect 13955 2941 13967 2975
rect 13909 2935 13967 2941
rect 7009 2907 7067 2913
rect 7009 2904 7021 2907
rect 6564 2876 7021 2904
rect 7009 2873 7021 2876
rect 7055 2873 7067 2907
rect 7009 2867 7067 2873
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 8481 2907 8539 2913
rect 8481 2904 8493 2907
rect 8352 2876 8493 2904
rect 8352 2864 8358 2876
rect 8481 2873 8493 2876
rect 8527 2873 8539 2907
rect 8481 2867 8539 2873
rect 8573 2907 8631 2913
rect 8573 2873 8585 2907
rect 8619 2873 8631 2907
rect 8573 2867 8631 2873
rect 3234 2836 3240 2848
rect 2694 2808 3240 2836
rect 3234 2796 3240 2808
rect 3292 2796 3298 2848
rect 4246 2836 4252 2848
rect 4207 2808 4252 2836
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 5074 2836 5080 2848
rect 5035 2808 5080 2836
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 5534 2796 5540 2848
rect 5592 2836 5598 2848
rect 6638 2836 6644 2848
rect 5592 2808 6644 2836
rect 5592 2796 5598 2808
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 7156 2808 8217 2836
rect 7156 2796 7162 2808
rect 8205 2805 8217 2808
rect 8251 2836 8263 2839
rect 8588 2836 8616 2867
rect 8251 2808 8616 2836
rect 8251 2805 8263 2808
rect 8205 2799 8263 2805
rect 11974 2796 11980 2848
rect 12032 2836 12038 2848
rect 12575 2839 12633 2845
rect 12575 2836 12587 2839
rect 12032 2808 12587 2836
rect 12032 2796 12038 2808
rect 12575 2805 12587 2808
rect 12621 2805 12633 2839
rect 13262 2836 13268 2848
rect 13223 2808 13268 2836
rect 12575 2799 12633 2805
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2774 2632 2780 2644
rect 1995 2604 2780 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 1464 2499 1522 2505
rect 1464 2465 1476 2499
rect 1510 2496 1522 2499
rect 1964 2496 1992 2595
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 3326 2632 3332 2644
rect 3160 2604 3332 2632
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 2590 2564 2596 2576
rect 2363 2536 2596 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 2590 2524 2596 2536
rect 2648 2524 2654 2576
rect 3160 2573 3188 2604
rect 3326 2592 3332 2604
rect 3384 2632 3390 2644
rect 7745 2635 7803 2641
rect 7745 2632 7757 2635
rect 3384 2604 7757 2632
rect 3384 2592 3390 2604
rect 7745 2601 7757 2604
rect 7791 2601 7803 2635
rect 10042 2632 10048 2644
rect 10003 2604 10048 2632
rect 7745 2595 7803 2601
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 3145 2567 3203 2573
rect 3145 2533 3157 2567
rect 3191 2533 3203 2567
rect 3145 2527 3203 2533
rect 3234 2524 3240 2576
rect 3292 2564 3298 2576
rect 3881 2567 3939 2573
rect 3881 2564 3893 2567
rect 3292 2536 3893 2564
rect 3292 2524 3298 2536
rect 3881 2533 3893 2536
rect 3927 2564 3939 2567
rect 4427 2567 4485 2573
rect 4427 2564 4439 2567
rect 3927 2536 4439 2564
rect 3927 2533 3939 2536
rect 3881 2527 3939 2533
rect 4427 2533 4439 2536
rect 4473 2564 4485 2567
rect 5074 2564 5080 2576
rect 4473 2536 5080 2564
rect 4473 2533 4485 2536
rect 4427 2527 4485 2533
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 5350 2564 5356 2576
rect 5311 2536 5356 2564
rect 5350 2524 5356 2536
rect 5408 2524 5414 2576
rect 5951 2567 6009 2573
rect 5951 2533 5963 2567
rect 5997 2564 6009 2567
rect 7006 2564 7012 2576
rect 5997 2536 7012 2564
rect 5997 2533 6009 2536
rect 5951 2527 6009 2533
rect 7006 2524 7012 2536
rect 7064 2524 7070 2576
rect 7098 2524 7104 2576
rect 7156 2564 7162 2576
rect 7156 2536 7201 2564
rect 7156 2524 7162 2536
rect 1510 2468 1992 2496
rect 3513 2499 3571 2505
rect 1510 2465 1522 2468
rect 1464 2459 1522 2465
rect 3513 2465 3525 2499
rect 3559 2496 3571 2499
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3559 2468 4077 2496
rect 3559 2465 3571 2468
rect 3513 2459 3571 2465
rect 4065 2465 4077 2468
rect 4111 2496 4123 2499
rect 4522 2496 4528 2508
rect 4111 2468 4528 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 5848 2499 5906 2505
rect 5848 2496 5860 2499
rect 5592 2468 5860 2496
rect 5592 2456 5598 2468
rect 5848 2465 5860 2468
rect 5894 2496 5906 2499
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5894 2468 6285 2496
rect 5894 2465 5906 2468
rect 5848 2459 5906 2465
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2496 8539 2499
rect 8570 2496 8576 2508
rect 8527 2468 8576 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 8570 2456 8576 2468
rect 8628 2496 8634 2508
rect 9033 2499 9091 2505
rect 9033 2496 9045 2499
rect 8628 2468 9045 2496
rect 8628 2456 8634 2468
rect 9033 2465 9045 2468
rect 9079 2465 9091 2499
rect 9858 2496 9864 2508
rect 9819 2468 9864 2496
rect 9033 2459 9091 2465
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 10962 2456 10968 2508
rect 11020 2496 11026 2508
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 11020 2468 11437 2496
rect 11020 2456 11026 2468
rect 11425 2465 11437 2468
rect 11471 2496 11483 2499
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11471 2468 11989 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12656 2499 12714 2505
rect 12656 2496 12668 2499
rect 12584 2468 12668 2496
rect 12584 2456 12590 2468
rect 12656 2465 12668 2468
rect 12702 2496 12714 2499
rect 13081 2499 13139 2505
rect 13081 2496 13093 2499
rect 12702 2468 13093 2496
rect 12702 2465 12714 2468
rect 12656 2459 12714 2465
rect 13081 2465 13093 2468
rect 13127 2496 13139 2499
rect 13262 2496 13268 2508
rect 13127 2468 13268 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 13262 2456 13268 2468
rect 13320 2456 13326 2508
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 5718 2428 5724 2440
rect 2547 2400 5724 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7055 2400 8033 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 8021 2397 8033 2400
rect 8067 2428 8079 2431
rect 12759 2431 12817 2437
rect 12759 2428 12771 2431
rect 8067 2400 12771 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 12759 2397 12771 2400
rect 12805 2397 12817 2431
rect 12759 2391 12817 2397
rect 5994 2320 6000 2372
rect 6052 2360 6058 2372
rect 9493 2363 9551 2369
rect 9493 2360 9505 2363
rect 6052 2332 9505 2360
rect 6052 2320 6058 2332
rect 9493 2329 9505 2332
rect 9539 2360 9551 2363
rect 9858 2360 9864 2372
rect 9539 2332 9864 2360
rect 9539 2329 9551 2332
rect 9493 2323 9551 2329
rect 9858 2320 9864 2332
rect 9916 2320 9922 2372
rect 11609 2363 11667 2369
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 13354 2360 13360 2372
rect 11655 2332 13360 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 13354 2320 13360 2332
rect 13412 2320 13418 2372
rect 1535 2295 1593 2301
rect 1535 2261 1547 2295
rect 1581 2292 1593 2295
rect 1762 2292 1768 2304
rect 1581 2264 1768 2292
rect 1581 2261 1593 2264
rect 1535 2255 1593 2261
rect 1762 2252 1768 2264
rect 1820 2252 1826 2304
rect 4985 2295 5043 2301
rect 4985 2261 4997 2295
rect 5031 2292 5043 2295
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 5031 2264 6653 2292
rect 5031 2261 5043 2264
rect 4985 2255 5043 2261
rect 6641 2261 6653 2264
rect 6687 2292 6699 2295
rect 7098 2292 7104 2304
rect 6687 2264 7104 2292
rect 6687 2261 6699 2264
rect 6641 2255 6699 2261
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 8294 2292 8300 2304
rect 8255 2264 8300 2292
rect 8294 2252 8300 2264
rect 8352 2252 8358 2304
rect 8662 2292 8668 2304
rect 8623 2264 8668 2292
rect 8662 2252 8668 2264
rect 8720 2252 8726 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 1762 2048 1768 2100
rect 1820 2088 1826 2100
rect 7742 2088 7748 2100
rect 1820 2060 7748 2088
rect 1820 2048 1826 2060
rect 7742 2048 7748 2060
rect 7800 2088 7806 2100
rect 8294 2088 8300 2100
rect 7800 2060 8300 2088
rect 7800 2048 7806 2060
rect 8294 2048 8300 2060
rect 8352 2048 8358 2100
rect 1486 1980 1492 2032
rect 1544 2020 1550 2032
rect 5534 2020 5540 2032
rect 1544 1992 5540 2020
rect 1544 1980 1550 1992
rect 5534 1980 5540 1992
rect 5592 1980 5598 2032
rect 5074 1912 5080 1964
rect 5132 1952 5138 1964
rect 10226 1952 10232 1964
rect 5132 1924 10232 1952
rect 5132 1912 5138 1924
rect 10226 1912 10232 1924
rect 10284 1912 10290 1964
rect 4062 1776 4068 1828
rect 4120 1816 4126 1828
rect 4120 1776 4154 1816
rect 4126 1748 4154 1776
rect 5258 1748 5264 1760
rect 4126 1720 5264 1748
rect 5258 1708 5264 1720
rect 5316 1708 5322 1760
rect 8662 1164 8668 1216
rect 8720 1204 8726 1216
rect 13722 1204 13728 1216
rect 8720 1176 13728 1204
rect 8720 1164 8726 1176
rect 13722 1164 13728 1176
rect 13780 1164 13786 1216
rect 290 76 296 128
rect 348 116 354 128
rect 1026 116 1032 128
rect 348 88 1032 116
rect 348 76 354 88
rect 1026 76 1032 88
rect 1084 76 1090 128
rect 1486 76 1492 128
rect 1544 116 1550 128
rect 2038 116 2044 128
rect 1544 88 2044 116
rect 1544 76 1550 88
rect 2038 76 2044 88
rect 2096 76 2102 128
rect 4246 76 4252 128
rect 4304 116 4310 128
rect 12066 116 12072 128
rect 4304 88 12072 116
rect 4304 76 4310 88
rect 12066 76 12072 88
rect 12124 76 12130 128
rect 842 8 848 60
rect 900 48 906 60
rect 5166 48 5172 60
rect 900 20 5172 48
rect 900 8 906 20
rect 5166 8 5172 20
rect 5224 8 5230 60
<< via1 >>
rect 388 39652 440 39704
rect 6184 39720 6236 39772
rect 5540 39652 5592 39704
rect 6552 39652 6604 39704
rect 1492 39584 1544 39636
rect 2136 39584 2188 39636
rect 3056 39584 3108 39636
rect 3884 39584 3936 39636
rect 5080 39584 5132 39636
rect 5724 39584 5776 39636
rect 7472 39584 7524 39636
rect 8024 39584 8076 39636
rect 13820 39584 13872 39636
rect 15476 39584 15528 39636
rect 9404 39516 9456 39568
rect 5816 39448 5868 39500
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 8116 35232 8168 35284
rect 7656 35139 7708 35148
rect 7656 35105 7665 35139
rect 7665 35105 7699 35139
rect 7699 35105 7708 35139
rect 7656 35096 7708 35105
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 9772 34688 9824 34740
rect 10692 34688 10744 34740
rect 14648 34688 14700 34740
rect 4620 34552 4672 34604
rect 13452 34620 13504 34672
rect 12532 34552 12584 34604
rect 8300 34527 8352 34536
rect 8300 34493 8309 34527
rect 8309 34493 8343 34527
rect 8343 34493 8352 34527
rect 8300 34484 8352 34493
rect 9312 34484 9364 34536
rect 11980 34484 12032 34536
rect 5264 34348 5316 34400
rect 7656 34348 7708 34400
rect 10508 34348 10560 34400
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 8852 34144 8904 34196
rect 8116 34051 8168 34060
rect 8116 34017 8125 34051
rect 8125 34017 8159 34051
rect 8159 34017 8168 34051
rect 8116 34008 8168 34017
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 5632 33260 5684 33312
rect 8116 33303 8168 33312
rect 8116 33269 8125 33303
rect 8125 33269 8159 33303
rect 8159 33269 8168 33303
rect 8116 33260 8168 33269
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 1032 30336 1084 30388
rect 3148 29996 3200 30048
rect 10048 29996 10100 30048
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 7104 29792 7156 29844
rect 6092 29767 6144 29776
rect 6092 29733 6101 29767
rect 6101 29733 6135 29767
rect 6135 29733 6144 29767
rect 6092 29724 6144 29733
rect 7840 29656 7892 29708
rect 6000 29631 6052 29640
rect 6000 29597 6009 29631
rect 6009 29597 6043 29631
rect 6043 29597 6052 29631
rect 6000 29588 6052 29597
rect 7196 29588 7248 29640
rect 6276 29452 6328 29504
rect 8300 29452 8352 29504
rect 8484 29495 8536 29504
rect 8484 29461 8493 29495
rect 8493 29461 8527 29495
rect 8527 29461 8536 29495
rect 8484 29452 8536 29461
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 5908 29248 5960 29300
rect 6276 29291 6328 29300
rect 6276 29257 6285 29291
rect 6285 29257 6319 29291
rect 6319 29257 6328 29291
rect 6276 29248 6328 29257
rect 7840 29291 7892 29300
rect 7840 29257 7849 29291
rect 7849 29257 7883 29291
rect 7883 29257 7892 29291
rect 7840 29248 7892 29257
rect 6184 29180 6236 29232
rect 7104 29180 7156 29232
rect 7288 29112 7340 29164
rect 10600 29112 10652 29164
rect 6276 29044 6328 29096
rect 6920 29019 6972 29028
rect 6920 28985 6929 29019
rect 6929 28985 6963 29019
rect 6963 28985 6972 29019
rect 6920 28976 6972 28985
rect 5080 28908 5132 28960
rect 6092 28908 6144 28960
rect 6644 28951 6696 28960
rect 6644 28917 6653 28951
rect 6653 28917 6687 28951
rect 6687 28917 6696 28951
rect 7196 28976 7248 29028
rect 8484 29019 8536 29028
rect 8484 28985 8493 29019
rect 8493 28985 8527 29019
rect 8527 28985 8536 29019
rect 8484 28976 8536 28985
rect 8576 29019 8628 29028
rect 8576 28985 8585 29019
rect 8585 28985 8619 29019
rect 8619 28985 8628 29019
rect 8576 28976 8628 28985
rect 6644 28908 6696 28917
rect 7656 28908 7708 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 6000 28704 6052 28756
rect 6920 28747 6972 28756
rect 6920 28713 6929 28747
rect 6929 28713 6963 28747
rect 6963 28713 6972 28747
rect 6920 28704 6972 28713
rect 7288 28747 7340 28756
rect 7288 28713 7297 28747
rect 7297 28713 7331 28747
rect 7331 28713 7340 28747
rect 7288 28704 7340 28713
rect 6092 28679 6144 28688
rect 6092 28645 6101 28679
rect 6101 28645 6135 28679
rect 6135 28645 6144 28679
rect 6092 28636 6144 28645
rect 7656 28679 7708 28688
rect 7656 28645 7665 28679
rect 7665 28645 7699 28679
rect 7699 28645 7708 28679
rect 7656 28636 7708 28645
rect 1492 28568 1544 28620
rect 4988 28568 5040 28620
rect 9588 28611 9640 28620
rect 9588 28577 9597 28611
rect 9597 28577 9631 28611
rect 9631 28577 9640 28611
rect 9588 28568 9640 28577
rect 4436 28500 4488 28552
rect 6000 28543 6052 28552
rect 6000 28509 6009 28543
rect 6009 28509 6043 28543
rect 6043 28509 6052 28543
rect 6000 28500 6052 28509
rect 7012 28500 7064 28552
rect 5356 28407 5408 28416
rect 5356 28373 5365 28407
rect 5365 28373 5399 28407
rect 5399 28373 5408 28407
rect 5356 28364 5408 28373
rect 8208 28364 8260 28416
rect 9312 28364 9364 28416
rect 9680 28364 9732 28416
rect 10416 28364 10468 28416
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 4436 28160 4488 28212
rect 4620 28203 4672 28212
rect 4620 28169 4629 28203
rect 4629 28169 4663 28203
rect 4663 28169 4672 28203
rect 4620 28160 4672 28169
rect 4988 28203 5040 28212
rect 4988 28169 4997 28203
rect 4997 28169 5031 28203
rect 5031 28169 5040 28203
rect 4988 28160 5040 28169
rect 7656 28160 7708 28212
rect 10048 28203 10100 28212
rect 10048 28169 10057 28203
rect 10057 28169 10091 28203
rect 10091 28169 10100 28203
rect 10048 28160 10100 28169
rect 3976 28092 4028 28144
rect 5540 28092 5592 28144
rect 5724 28092 5776 28144
rect 10416 28092 10468 28144
rect 10048 28024 10100 28076
rect 10600 28067 10652 28076
rect 10600 28033 10609 28067
rect 10609 28033 10643 28067
rect 10643 28033 10652 28067
rect 10600 28024 10652 28033
rect 6920 27999 6972 28008
rect 3332 27888 3384 27940
rect 6920 27965 6929 27999
rect 6929 27965 6963 27999
rect 6963 27965 6972 27999
rect 6920 27956 6972 27965
rect 4620 27888 4672 27940
rect 4988 27888 5040 27940
rect 5356 27931 5408 27940
rect 5356 27897 5365 27931
rect 5365 27897 5399 27931
rect 5399 27897 5408 27931
rect 5356 27888 5408 27897
rect 7012 27888 7064 27940
rect 8760 27931 8812 27940
rect 5540 27820 5592 27872
rect 6092 27820 6144 27872
rect 6736 27820 6788 27872
rect 8760 27897 8769 27931
rect 8769 27897 8803 27931
rect 8803 27897 8812 27931
rect 8760 27888 8812 27897
rect 9404 27931 9456 27940
rect 8300 27820 8352 27872
rect 9404 27897 9413 27931
rect 9413 27897 9447 27931
rect 9447 27897 9456 27931
rect 9404 27888 9456 27897
rect 9864 27888 9916 27940
rect 10416 27931 10468 27940
rect 10416 27897 10425 27931
rect 10425 27897 10459 27931
rect 10459 27897 10468 27931
rect 10416 27888 10468 27897
rect 9588 27820 9640 27872
rect 12072 27820 12124 27872
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 4988 27659 5040 27668
rect 4988 27625 4997 27659
rect 4997 27625 5031 27659
rect 5031 27625 5040 27659
rect 4988 27616 5040 27625
rect 6000 27616 6052 27668
rect 8300 27659 8352 27668
rect 8300 27625 8309 27659
rect 8309 27625 8343 27659
rect 8343 27625 8352 27659
rect 8300 27616 8352 27625
rect 9680 27616 9732 27668
rect 5172 27548 5224 27600
rect 8116 27548 8168 27600
rect 9864 27591 9916 27600
rect 9864 27557 9873 27591
rect 9873 27557 9907 27591
rect 9907 27557 9916 27591
rect 9864 27548 9916 27557
rect 3240 27480 3292 27532
rect 4344 27480 4396 27532
rect 6644 27480 6696 27532
rect 10508 27480 10560 27532
rect 11244 27523 11296 27532
rect 11244 27489 11288 27523
rect 11288 27489 11296 27523
rect 11244 27480 11296 27489
rect 4988 27412 5040 27464
rect 7380 27455 7432 27464
rect 2964 27344 3016 27396
rect 7380 27421 7389 27455
rect 7389 27421 7423 27455
rect 7423 27421 7432 27455
rect 7380 27412 7432 27421
rect 8760 27455 8812 27464
rect 8760 27421 8769 27455
rect 8769 27421 8803 27455
rect 8803 27421 8812 27455
rect 8760 27412 8812 27421
rect 6184 27344 6236 27396
rect 8484 27344 8536 27396
rect 9956 27344 10008 27396
rect 3516 27319 3568 27328
rect 3516 27285 3525 27319
rect 3525 27285 3559 27319
rect 3559 27285 3568 27319
rect 3516 27276 3568 27285
rect 4068 27276 4120 27328
rect 6920 27276 6972 27328
rect 7564 27276 7616 27328
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 3240 27115 3292 27124
rect 3240 27081 3249 27115
rect 3249 27081 3283 27115
rect 3283 27081 3292 27115
rect 3240 27072 3292 27081
rect 4344 27072 4396 27124
rect 6092 27072 6144 27124
rect 9864 27072 9916 27124
rect 11244 27115 11296 27124
rect 11244 27081 11253 27115
rect 11253 27081 11287 27115
rect 11287 27081 11296 27115
rect 11244 27072 11296 27081
rect 12348 27072 12400 27124
rect 5724 27004 5776 27056
rect 10416 27004 10468 27056
rect 3516 26979 3568 26988
rect 3516 26945 3525 26979
rect 3525 26945 3559 26979
rect 3559 26945 3568 26979
rect 3516 26936 3568 26945
rect 6184 26979 6236 26988
rect 6184 26945 6193 26979
rect 6193 26945 6227 26979
rect 6227 26945 6236 26979
rect 6184 26936 6236 26945
rect 6736 26936 6788 26988
rect 2412 26732 2464 26784
rect 3608 26843 3660 26852
rect 3608 26809 3617 26843
rect 3617 26809 3651 26843
rect 3651 26809 3660 26843
rect 3608 26800 3660 26809
rect 4896 26800 4948 26852
rect 5172 26800 5224 26852
rect 3332 26732 3384 26784
rect 4988 26732 5040 26784
rect 6920 26732 6972 26784
rect 8116 26936 8168 26988
rect 10600 26936 10652 26988
rect 8760 26775 8812 26784
rect 8760 26741 8769 26775
rect 8769 26741 8803 26775
rect 8803 26741 8812 26775
rect 8760 26732 8812 26741
rect 9404 26843 9456 26852
rect 9404 26809 9413 26843
rect 9413 26809 9447 26843
rect 9447 26809 9456 26843
rect 9404 26800 9456 26809
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 2412 26528 2464 26580
rect 3516 26528 3568 26580
rect 5356 26528 5408 26580
rect 6644 26528 6696 26580
rect 8576 26528 8628 26580
rect 9680 26528 9732 26580
rect 3148 26460 3200 26512
rect 4988 26460 5040 26512
rect 8116 26460 8168 26512
rect 4160 26435 4212 26444
rect 4160 26401 4178 26435
rect 4178 26401 4212 26435
rect 4160 26392 4212 26401
rect 5540 26392 5592 26444
rect 6736 26392 6788 26444
rect 4436 26324 4488 26376
rect 6000 26324 6052 26376
rect 9312 26324 9364 26376
rect 3516 26231 3568 26240
rect 3516 26197 3525 26231
rect 3525 26197 3559 26231
rect 3559 26197 3568 26231
rect 3516 26188 3568 26197
rect 4712 26188 4764 26240
rect 4988 26188 5040 26240
rect 7380 26188 7432 26240
rect 8484 26188 8536 26240
rect 9404 26231 9456 26240
rect 9404 26197 9413 26231
rect 9413 26197 9447 26231
rect 9447 26197 9456 26231
rect 9404 26188 9456 26197
rect 10692 26188 10744 26240
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 4160 26027 4212 26036
rect 4160 25993 4169 26027
rect 4169 25993 4203 26027
rect 4203 25993 4212 26027
rect 4160 25984 4212 25993
rect 5172 25984 5224 26036
rect 5632 25984 5684 26036
rect 6644 26027 6696 26036
rect 6644 25993 6653 26027
rect 6653 25993 6687 26027
rect 6687 25993 6696 26027
rect 6644 25984 6696 25993
rect 3148 25916 3200 25968
rect 4896 25891 4948 25900
rect 1308 25780 1360 25832
rect 2320 25780 2372 25832
rect 3424 25780 3476 25832
rect 3516 25780 3568 25832
rect 4252 25780 4304 25832
rect 4896 25857 4905 25891
rect 4905 25857 4939 25891
rect 4939 25857 4948 25891
rect 4896 25848 4948 25857
rect 6736 25848 6788 25900
rect 7196 25848 7248 25900
rect 8852 25848 8904 25900
rect 4620 25755 4672 25764
rect 2596 25687 2648 25696
rect 2596 25653 2605 25687
rect 2605 25653 2639 25687
rect 2639 25653 2648 25687
rect 4620 25721 4629 25755
rect 4629 25721 4663 25755
rect 4663 25721 4672 25755
rect 4620 25712 4672 25721
rect 4712 25755 4764 25764
rect 4712 25721 4721 25755
rect 4721 25721 4755 25755
rect 4755 25721 4764 25755
rect 4712 25712 4764 25721
rect 8668 25755 8720 25764
rect 2596 25644 2648 25653
rect 4988 25644 5040 25696
rect 6000 25687 6052 25696
rect 6000 25653 6009 25687
rect 6009 25653 6043 25687
rect 6043 25653 6052 25687
rect 6000 25644 6052 25653
rect 6644 25644 6696 25696
rect 8668 25721 8677 25755
rect 8677 25721 8711 25755
rect 8711 25721 8720 25755
rect 8668 25712 8720 25721
rect 9864 25712 9916 25764
rect 8116 25644 8168 25696
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 2596 25483 2648 25492
rect 2596 25449 2605 25483
rect 2605 25449 2639 25483
rect 2639 25449 2648 25483
rect 2596 25440 2648 25449
rect 4620 25440 4672 25492
rect 6000 25440 6052 25492
rect 13820 25440 13872 25492
rect 4252 25415 4304 25424
rect 4252 25381 4261 25415
rect 4261 25381 4295 25415
rect 4295 25381 4304 25415
rect 4252 25372 4304 25381
rect 4988 25372 5040 25424
rect 5448 25372 5500 25424
rect 7656 25347 7708 25356
rect 2228 25279 2280 25288
rect 2228 25245 2237 25279
rect 2237 25245 2271 25279
rect 2271 25245 2280 25279
rect 2228 25236 2280 25245
rect 4160 25279 4212 25288
rect 4160 25245 4169 25279
rect 4169 25245 4203 25279
rect 4203 25245 4212 25279
rect 4160 25236 4212 25245
rect 4436 25279 4488 25288
rect 4436 25245 4445 25279
rect 4445 25245 4479 25279
rect 4479 25245 4488 25279
rect 4436 25236 4488 25245
rect 3148 25211 3200 25220
rect 3148 25177 3157 25211
rect 3157 25177 3191 25211
rect 3191 25177 3200 25211
rect 3148 25168 3200 25177
rect 4620 25168 4672 25220
rect 5540 25236 5592 25288
rect 7656 25313 7665 25347
rect 7665 25313 7699 25347
rect 7699 25313 7708 25347
rect 7656 25304 7708 25313
rect 8392 25304 8444 25356
rect 10968 25304 11020 25356
rect 7840 25236 7892 25288
rect 3424 25143 3476 25152
rect 3424 25109 3433 25143
rect 3433 25109 3467 25143
rect 3467 25109 3476 25143
rect 3424 25100 3476 25109
rect 3516 25100 3568 25152
rect 7288 25100 7340 25152
rect 7656 25100 7708 25152
rect 8300 25100 8352 25152
rect 8852 25143 8904 25152
rect 8852 25109 8861 25143
rect 8861 25109 8895 25143
rect 8895 25109 8904 25143
rect 8852 25100 8904 25109
rect 10048 25143 10100 25152
rect 10048 25109 10057 25143
rect 10057 25109 10091 25143
rect 10091 25109 10100 25143
rect 10048 25100 10100 25109
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 2964 24803 3016 24812
rect 2964 24769 2973 24803
rect 2973 24769 3007 24803
rect 3007 24769 3016 24803
rect 2964 24760 3016 24769
rect 1952 24692 2004 24744
rect 3516 24896 3568 24948
rect 4988 24939 5040 24948
rect 4988 24905 4997 24939
rect 4997 24905 5031 24939
rect 5031 24905 5040 24939
rect 4988 24896 5040 24905
rect 5448 24939 5500 24948
rect 5448 24905 5457 24939
rect 5457 24905 5491 24939
rect 5491 24905 5500 24939
rect 5448 24896 5500 24905
rect 10968 24939 11020 24948
rect 10968 24905 10977 24939
rect 10977 24905 11011 24939
rect 11011 24905 11020 24939
rect 10968 24896 11020 24905
rect 4252 24828 4304 24880
rect 4344 24760 4396 24812
rect 4988 24760 5040 24812
rect 5264 24760 5316 24812
rect 3884 24692 3936 24744
rect 6736 24760 6788 24812
rect 10048 24803 10100 24812
rect 10048 24769 10057 24803
rect 10057 24769 10091 24803
rect 10091 24769 10100 24803
rect 10048 24760 10100 24769
rect 7288 24735 7340 24744
rect 4528 24624 4580 24676
rect 7288 24701 7297 24735
rect 7297 24701 7331 24735
rect 7331 24701 7340 24735
rect 7288 24692 7340 24701
rect 8300 24692 8352 24744
rect 2596 24556 2648 24608
rect 3976 24556 4028 24608
rect 4160 24599 4212 24608
rect 4160 24565 4169 24599
rect 4169 24565 4203 24599
rect 4203 24565 4212 24599
rect 4160 24556 4212 24565
rect 4344 24556 4396 24608
rect 4804 24556 4856 24608
rect 6920 24599 6972 24608
rect 6920 24565 6929 24599
rect 6929 24565 6963 24599
rect 6963 24565 6972 24599
rect 6920 24556 6972 24565
rect 7840 24599 7892 24608
rect 7840 24565 7849 24599
rect 7849 24565 7883 24599
rect 7883 24565 7892 24599
rect 7840 24556 7892 24565
rect 7932 24556 7984 24608
rect 8484 24599 8536 24608
rect 8484 24565 8493 24599
rect 8493 24565 8527 24599
rect 8527 24565 8536 24599
rect 8484 24556 8536 24565
rect 9588 24556 9640 24608
rect 10692 24667 10744 24676
rect 10692 24633 10701 24667
rect 10701 24633 10735 24667
rect 10735 24633 10744 24667
rect 10692 24624 10744 24633
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 2228 24352 2280 24404
rect 4712 24352 4764 24404
rect 7288 24395 7340 24404
rect 7288 24361 7297 24395
rect 7297 24361 7331 24395
rect 7331 24361 7340 24395
rect 7288 24352 7340 24361
rect 7564 24395 7616 24404
rect 7564 24361 7573 24395
rect 7573 24361 7607 24395
rect 7607 24361 7616 24395
rect 7564 24352 7616 24361
rect 11520 24352 11572 24404
rect 4252 24327 4304 24336
rect 4252 24293 4261 24327
rect 4261 24293 4295 24327
rect 4295 24293 4304 24327
rect 4252 24284 4304 24293
rect 4896 24284 4948 24336
rect 6092 24327 6144 24336
rect 6092 24293 6101 24327
rect 6101 24293 6135 24327
rect 6135 24293 6144 24327
rect 6092 24284 6144 24293
rect 9588 24284 9640 24336
rect 2688 24259 2740 24268
rect 2688 24225 2697 24259
rect 2697 24225 2731 24259
rect 2731 24225 2740 24259
rect 2688 24216 2740 24225
rect 7472 24259 7524 24268
rect 7472 24225 7481 24259
rect 7481 24225 7515 24259
rect 7515 24225 7524 24259
rect 7472 24216 7524 24225
rect 7932 24259 7984 24268
rect 7932 24225 7941 24259
rect 7941 24225 7975 24259
rect 7975 24225 7984 24259
rect 7932 24216 7984 24225
rect 11244 24259 11296 24268
rect 11244 24225 11253 24259
rect 11253 24225 11287 24259
rect 11287 24225 11296 24259
rect 11244 24216 11296 24225
rect 3148 24148 3200 24200
rect 4344 24148 4396 24200
rect 5724 24148 5776 24200
rect 7380 24148 7432 24200
rect 9772 24191 9824 24200
rect 9772 24157 9781 24191
rect 9781 24157 9815 24191
rect 9815 24157 9824 24191
rect 9772 24148 9824 24157
rect 9864 24148 9916 24200
rect 4528 24080 4580 24132
rect 5264 24080 5316 24132
rect 7196 24080 7248 24132
rect 3976 24012 4028 24064
rect 4160 24012 4212 24064
rect 4620 24012 4672 24064
rect 5540 24012 5592 24064
rect 8484 24055 8536 24064
rect 8484 24021 8493 24055
rect 8493 24021 8527 24055
rect 8527 24021 8536 24055
rect 8484 24012 8536 24021
rect 11520 24012 11572 24064
rect 12716 24012 12768 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 1952 23851 2004 23860
rect 1952 23817 1961 23851
rect 1961 23817 1995 23851
rect 1995 23817 2004 23851
rect 1952 23808 2004 23817
rect 4252 23808 4304 23860
rect 6092 23808 6144 23860
rect 7932 23808 7984 23860
rect 8668 23851 8720 23860
rect 8668 23817 8677 23851
rect 8677 23817 8711 23851
rect 8711 23817 8720 23851
rect 8668 23808 8720 23817
rect 9772 23808 9824 23860
rect 3424 23672 3476 23724
rect 1952 23604 2004 23656
rect 2136 23604 2188 23656
rect 2688 23604 2740 23656
rect 7840 23740 7892 23792
rect 4160 23715 4212 23724
rect 4160 23681 4169 23715
rect 4169 23681 4203 23715
rect 4203 23681 4212 23715
rect 4160 23672 4212 23681
rect 5632 23672 5684 23724
rect 8484 23672 8536 23724
rect 1584 23536 1636 23588
rect 3976 23604 4028 23656
rect 5264 23579 5316 23588
rect 5264 23545 5273 23579
rect 5273 23545 5307 23579
rect 5307 23545 5316 23579
rect 5264 23536 5316 23545
rect 5632 23536 5684 23588
rect 6000 23536 6052 23588
rect 7380 23536 7432 23588
rect 7932 23536 7984 23588
rect 8116 23536 8168 23588
rect 3148 23511 3200 23520
rect 3148 23477 3157 23511
rect 3157 23477 3191 23511
rect 3191 23477 3200 23511
rect 3148 23468 3200 23477
rect 5724 23468 5776 23520
rect 7748 23468 7800 23520
rect 10048 23604 10100 23656
rect 11244 23604 11296 23656
rect 9404 23468 9456 23520
rect 9680 23468 9732 23520
rect 10968 23468 11020 23520
rect 12164 23468 12216 23520
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 1124 23264 1176 23316
rect 4620 23264 4672 23316
rect 4804 23307 4856 23316
rect 4804 23273 4813 23307
rect 4813 23273 4847 23307
rect 4847 23273 4856 23307
rect 4804 23264 4856 23273
rect 5264 23307 5316 23316
rect 5264 23273 5273 23307
rect 5273 23273 5307 23307
rect 5307 23273 5316 23307
rect 5264 23264 5316 23273
rect 6092 23264 6144 23316
rect 7012 23264 7064 23316
rect 7472 23307 7524 23316
rect 7472 23273 7481 23307
rect 7481 23273 7515 23307
rect 7515 23273 7524 23307
rect 7472 23264 7524 23273
rect 9588 23264 9640 23316
rect 10968 23264 11020 23316
rect 4068 23196 4120 23248
rect 5540 23196 5592 23248
rect 7840 23196 7892 23248
rect 2044 23128 2096 23180
rect 3056 23128 3108 23180
rect 2596 23060 2648 23112
rect 3976 23060 4028 23112
rect 5080 23128 5132 23180
rect 8300 23128 8352 23180
rect 9404 23128 9456 23180
rect 9772 23171 9824 23180
rect 9772 23137 9781 23171
rect 9781 23137 9815 23171
rect 9815 23137 9824 23171
rect 9772 23128 9824 23137
rect 10048 23128 10100 23180
rect 11336 23128 11388 23180
rect 6644 23060 6696 23112
rect 7748 23103 7800 23112
rect 7748 23069 7757 23103
rect 7757 23069 7791 23103
rect 7791 23069 7800 23103
rect 7748 23060 7800 23069
rect 8576 23060 8628 23112
rect 2136 22992 2188 23044
rect 2780 22992 2832 23044
rect 6000 22992 6052 23044
rect 8852 22992 8904 23044
rect 1768 22924 1820 22976
rect 2688 22924 2740 22976
rect 5816 22924 5868 22976
rect 13268 22924 13320 22976
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 2044 22763 2096 22772
rect 2044 22729 2053 22763
rect 2053 22729 2087 22763
rect 2087 22729 2096 22763
rect 2044 22720 2096 22729
rect 2780 22720 2832 22772
rect 3056 22763 3108 22772
rect 3056 22729 3065 22763
rect 3065 22729 3099 22763
rect 3099 22729 3108 22763
rect 3056 22720 3108 22729
rect 4068 22720 4120 22772
rect 4436 22720 4488 22772
rect 5908 22720 5960 22772
rect 7288 22720 7340 22772
rect 5540 22652 5592 22704
rect 7840 22695 7892 22704
rect 7840 22661 7849 22695
rect 7849 22661 7883 22695
rect 7883 22661 7892 22695
rect 7840 22652 7892 22661
rect 4068 22627 4120 22636
rect 4068 22593 4077 22627
rect 4077 22593 4111 22627
rect 4111 22593 4120 22627
rect 4068 22584 4120 22593
rect 4252 22584 4304 22636
rect 5724 22627 5776 22636
rect 5724 22593 5733 22627
rect 5733 22593 5767 22627
rect 5767 22593 5776 22627
rect 5724 22584 5776 22593
rect 7012 22584 7064 22636
rect 7380 22627 7432 22636
rect 7380 22593 7389 22627
rect 7389 22593 7423 22627
rect 7423 22593 7432 22627
rect 7380 22584 7432 22593
rect 8760 22584 8812 22636
rect 10968 22652 11020 22704
rect 10692 22627 10744 22636
rect 10692 22593 10701 22627
rect 10701 22593 10735 22627
rect 10735 22593 10744 22627
rect 10692 22584 10744 22593
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 6092 22516 6144 22568
rect 8576 22559 8628 22568
rect 8576 22525 8585 22559
rect 8585 22525 8619 22559
rect 8619 22525 8628 22559
rect 8576 22516 8628 22525
rect 8852 22559 8904 22568
rect 8852 22525 8861 22559
rect 8861 22525 8895 22559
rect 8895 22525 8904 22559
rect 8852 22516 8904 22525
rect 4160 22491 4212 22500
rect 4160 22457 4169 22491
rect 4169 22457 4203 22491
rect 4203 22457 4212 22491
rect 4160 22448 4212 22457
rect 5908 22448 5960 22500
rect 8668 22448 8720 22500
rect 10508 22448 10560 22500
rect 1676 22423 1728 22432
rect 1676 22389 1685 22423
rect 1685 22389 1719 22423
rect 1719 22389 1728 22423
rect 1676 22380 1728 22389
rect 2228 22423 2280 22432
rect 2228 22389 2237 22423
rect 2237 22389 2271 22423
rect 2271 22389 2280 22423
rect 2228 22380 2280 22389
rect 5540 22423 5592 22432
rect 5540 22389 5549 22423
rect 5549 22389 5583 22423
rect 5583 22389 5592 22423
rect 5540 22380 5592 22389
rect 6644 22380 6696 22432
rect 8852 22380 8904 22432
rect 10048 22380 10100 22432
rect 11336 22423 11388 22432
rect 11336 22389 11345 22423
rect 11345 22389 11379 22423
rect 11379 22389 11388 22423
rect 11336 22380 11388 22389
rect 12440 22380 12492 22432
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 5540 22219 5592 22228
rect 5540 22185 5549 22219
rect 5549 22185 5583 22219
rect 5583 22185 5592 22219
rect 5540 22176 5592 22185
rect 5632 22176 5684 22228
rect 6644 22176 6696 22228
rect 7104 22176 7156 22228
rect 1308 22108 1360 22160
rect 2228 22108 2280 22160
rect 2596 22151 2648 22160
rect 2596 22117 2605 22151
rect 2605 22117 2639 22151
rect 2639 22117 2648 22151
rect 2596 22108 2648 22117
rect 4344 22040 4396 22092
rect 7472 22108 7524 22160
rect 1676 21972 1728 22024
rect 4252 21972 4304 22024
rect 5172 22015 5224 22024
rect 5172 21981 5181 22015
rect 5181 21981 5215 22015
rect 5215 21981 5224 22015
rect 5172 21972 5224 21981
rect 7196 21904 7248 21956
rect 8208 22040 8260 22092
rect 8392 22040 8444 22092
rect 9956 22176 10008 22228
rect 10508 22219 10560 22228
rect 10508 22185 10517 22219
rect 10517 22185 10551 22219
rect 10551 22185 10560 22219
rect 10508 22176 10560 22185
rect 9680 22083 9732 22092
rect 9680 22049 9724 22083
rect 9724 22049 9732 22083
rect 10692 22083 10744 22092
rect 9680 22040 9732 22049
rect 10692 22049 10701 22083
rect 10701 22049 10735 22083
rect 10735 22049 10744 22083
rect 10692 22040 10744 22049
rect 9864 21972 9916 22024
rect 10048 21904 10100 21956
rect 1768 21836 1820 21888
rect 3056 21836 3108 21888
rect 5080 21879 5132 21888
rect 5080 21845 5089 21879
rect 5089 21845 5123 21879
rect 5123 21845 5132 21879
rect 5080 21836 5132 21845
rect 7748 21836 7800 21888
rect 8484 21836 8536 21888
rect 8576 21836 8628 21888
rect 9312 21836 9364 21888
rect 9496 21836 9548 21888
rect 9772 21836 9824 21888
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 2228 21632 2280 21684
rect 4344 21632 4396 21684
rect 5908 21675 5960 21684
rect 5908 21641 5917 21675
rect 5917 21641 5951 21675
rect 5951 21641 5960 21675
rect 5908 21632 5960 21641
rect 7656 21632 7708 21684
rect 9680 21675 9732 21684
rect 9680 21641 9689 21675
rect 9689 21641 9723 21675
rect 9723 21641 9732 21675
rect 9680 21632 9732 21641
rect 7380 21564 7432 21616
rect 1676 21471 1728 21480
rect 1676 21437 1685 21471
rect 1685 21437 1719 21471
rect 1719 21437 1728 21471
rect 1676 21428 1728 21437
rect 1768 21428 1820 21480
rect 3148 21428 3200 21480
rect 5080 21428 5132 21480
rect 5908 21428 5960 21480
rect 7196 21428 7248 21480
rect 8576 21496 8628 21548
rect 10692 21539 10744 21548
rect 10692 21505 10701 21539
rect 10701 21505 10735 21539
rect 10735 21505 10744 21539
rect 10692 21496 10744 21505
rect 8668 21428 8720 21480
rect 8852 21471 8904 21480
rect 8852 21437 8861 21471
rect 8861 21437 8895 21471
rect 8895 21437 8904 21471
rect 8852 21428 8904 21437
rect 2872 21403 2924 21412
rect 2872 21369 2881 21403
rect 2881 21369 2915 21403
rect 2915 21369 2924 21403
rect 2872 21360 2924 21369
rect 3976 21292 4028 21344
rect 4620 21292 4672 21344
rect 5540 21360 5592 21412
rect 6000 21360 6052 21412
rect 6184 21335 6236 21344
rect 6184 21301 6193 21335
rect 6193 21301 6227 21335
rect 6227 21301 6236 21335
rect 6184 21292 6236 21301
rect 6920 21335 6972 21344
rect 6920 21301 6929 21335
rect 6929 21301 6963 21335
rect 6963 21301 6972 21335
rect 6920 21292 6972 21301
rect 8208 21335 8260 21344
rect 8208 21301 8217 21335
rect 8217 21301 8251 21335
rect 8251 21301 8260 21335
rect 8208 21292 8260 21301
rect 8484 21335 8536 21344
rect 8484 21301 8493 21335
rect 8493 21301 8527 21335
rect 8527 21301 8536 21335
rect 8484 21292 8536 21301
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 1676 21131 1728 21140
rect 1676 21097 1685 21131
rect 1685 21097 1719 21131
rect 1719 21097 1728 21131
rect 1676 21088 1728 21097
rect 2596 21088 2648 21140
rect 3148 21088 3200 21140
rect 4160 21088 4212 21140
rect 5908 21131 5960 21140
rect 5908 21097 5917 21131
rect 5917 21097 5951 21131
rect 5951 21097 5960 21131
rect 5908 21088 5960 21097
rect 7472 21088 7524 21140
rect 8852 21088 8904 21140
rect 2872 21020 2924 21072
rect 4620 21020 4672 21072
rect 5172 21020 5224 21072
rect 6920 21020 6972 21072
rect 8668 21020 8720 21072
rect 9864 21063 9916 21072
rect 9864 21029 9873 21063
rect 9873 21029 9907 21063
rect 9907 21029 9916 21063
rect 9864 21020 9916 21029
rect 4160 20952 4212 21004
rect 4712 20952 4764 21004
rect 5816 20995 5868 21004
rect 5816 20961 5825 20995
rect 5825 20961 5859 20995
rect 5859 20961 5868 20995
rect 5816 20952 5868 20961
rect 6184 20952 6236 21004
rect 2596 20884 2648 20936
rect 4068 20927 4120 20936
rect 4068 20893 4077 20927
rect 4077 20893 4111 20927
rect 4111 20893 4120 20927
rect 4068 20884 4120 20893
rect 7196 20952 7248 21004
rect 7656 20995 7708 21004
rect 7656 20961 7665 20995
rect 7665 20961 7699 20995
rect 7699 20961 7708 20995
rect 7656 20952 7708 20961
rect 7748 20952 7800 21004
rect 11060 20952 11112 21004
rect 7932 20927 7984 20936
rect 7932 20893 7941 20927
rect 7941 20893 7975 20927
rect 7975 20893 7984 20927
rect 7932 20884 7984 20893
rect 9956 20884 10008 20936
rect 10600 20884 10652 20936
rect 5356 20791 5408 20800
rect 5356 20757 5365 20791
rect 5365 20757 5399 20791
rect 5399 20757 5408 20791
rect 5356 20748 5408 20757
rect 6920 20791 6972 20800
rect 6920 20757 6929 20791
rect 6929 20757 6963 20791
rect 6963 20757 6972 20791
rect 6920 20748 6972 20757
rect 10416 20748 10468 20800
rect 10784 20748 10836 20800
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 2872 20587 2924 20596
rect 2872 20553 2881 20587
rect 2881 20553 2915 20587
rect 2915 20553 2924 20587
rect 2872 20544 2924 20553
rect 4620 20544 4672 20596
rect 5356 20544 5408 20596
rect 6644 20544 6696 20596
rect 7472 20544 7524 20596
rect 9864 20544 9916 20596
rect 4160 20476 4212 20528
rect 6920 20476 6972 20528
rect 12992 20476 13044 20528
rect 1768 20451 1820 20460
rect 1768 20417 1777 20451
rect 1777 20417 1811 20451
rect 1811 20417 1820 20451
rect 1768 20408 1820 20417
rect 1860 20383 1912 20392
rect 1860 20349 1869 20383
rect 1869 20349 1903 20383
rect 1903 20349 1912 20383
rect 1860 20340 1912 20349
rect 4252 20451 4304 20460
rect 4252 20417 4261 20451
rect 4261 20417 4295 20451
rect 4295 20417 4304 20451
rect 4252 20408 4304 20417
rect 10416 20408 10468 20460
rect 2964 20340 3016 20392
rect 5908 20340 5960 20392
rect 2596 20315 2648 20324
rect 2596 20281 2605 20315
rect 2605 20281 2639 20315
rect 2639 20281 2648 20315
rect 2596 20272 2648 20281
rect 3976 20272 4028 20324
rect 4160 20272 4212 20324
rect 5816 20272 5868 20324
rect 5540 20204 5592 20256
rect 8024 20340 8076 20392
rect 9772 20340 9824 20392
rect 8300 20272 8352 20324
rect 10600 20315 10652 20324
rect 8116 20204 8168 20256
rect 8760 20204 8812 20256
rect 10600 20281 10609 20315
rect 10609 20281 10643 20315
rect 10643 20281 10652 20315
rect 10600 20272 10652 20281
rect 11060 20204 11112 20256
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 1584 20043 1636 20052
rect 1584 20009 1593 20043
rect 1593 20009 1627 20043
rect 1627 20009 1636 20043
rect 1584 20000 1636 20009
rect 2596 20000 2648 20052
rect 4068 19932 4120 19984
rect 4896 20000 4948 20052
rect 6000 20000 6052 20052
rect 8116 20000 8168 20052
rect 8760 20043 8812 20052
rect 8760 20009 8769 20043
rect 8769 20009 8803 20043
rect 8803 20009 8812 20043
rect 8760 20000 8812 20009
rect 9772 20043 9824 20052
rect 9772 20009 9781 20043
rect 9781 20009 9815 20043
rect 9815 20009 9824 20043
rect 9772 20000 9824 20009
rect 12992 20043 13044 20052
rect 12992 20009 13001 20043
rect 13001 20009 13035 20043
rect 13035 20009 13044 20043
rect 12992 20000 13044 20009
rect 5264 19932 5316 19984
rect 5356 19932 5408 19984
rect 6368 19975 6420 19984
rect 6368 19941 6377 19975
rect 6377 19941 6411 19975
rect 6411 19941 6420 19975
rect 6368 19932 6420 19941
rect 8300 19932 8352 19984
rect 10048 19932 10100 19984
rect 11428 19975 11480 19984
rect 11428 19941 11437 19975
rect 11437 19941 11471 19975
rect 11471 19941 11480 19975
rect 11428 19932 11480 19941
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 2412 19728 2464 19780
rect 7932 19864 7984 19916
rect 9312 19864 9364 19916
rect 9680 19907 9732 19916
rect 9680 19873 9689 19907
rect 9689 19873 9723 19907
rect 9723 19873 9732 19907
rect 9680 19864 9732 19873
rect 9772 19864 9824 19916
rect 12624 19864 12676 19916
rect 2964 19796 3016 19848
rect 3240 19796 3292 19848
rect 3976 19728 4028 19780
rect 4160 19728 4212 19780
rect 5632 19796 5684 19848
rect 7748 19796 7800 19848
rect 11704 19796 11756 19848
rect 10600 19728 10652 19780
rect 11612 19728 11664 19780
rect 4068 19660 4120 19712
rect 5264 19660 5316 19712
rect 8024 19660 8076 19712
rect 9956 19660 10008 19712
rect 10784 19660 10836 19712
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 1768 19499 1820 19508
rect 1768 19465 1777 19499
rect 1777 19465 1811 19499
rect 1811 19465 1820 19499
rect 1768 19456 1820 19465
rect 4896 19499 4948 19508
rect 4896 19465 4905 19499
rect 4905 19465 4939 19499
rect 4939 19465 4948 19499
rect 4896 19456 4948 19465
rect 5264 19499 5316 19508
rect 5264 19465 5273 19499
rect 5273 19465 5307 19499
rect 5307 19465 5316 19499
rect 5264 19456 5316 19465
rect 6644 19499 6696 19508
rect 6644 19465 6653 19499
rect 6653 19465 6687 19499
rect 6687 19465 6696 19499
rect 6644 19456 6696 19465
rect 7932 19456 7984 19508
rect 9680 19456 9732 19508
rect 9956 19456 10008 19508
rect 11704 19499 11756 19508
rect 11704 19465 11713 19499
rect 11713 19465 11747 19499
rect 11747 19465 11756 19499
rect 11704 19456 11756 19465
rect 1584 19388 1636 19440
rect 7196 19388 7248 19440
rect 7472 19388 7524 19440
rect 3976 19320 4028 19372
rect 6368 19320 6420 19372
rect 10600 19388 10652 19440
rect 2596 19252 2648 19304
rect 2780 19295 2832 19304
rect 2780 19261 2789 19295
rect 2789 19261 2823 19295
rect 2823 19261 2832 19295
rect 2780 19252 2832 19261
rect 4804 19252 4856 19304
rect 6184 19252 6236 19304
rect 6644 19252 6696 19304
rect 7840 19320 7892 19372
rect 8116 19363 8168 19372
rect 8116 19329 8125 19363
rect 8125 19329 8159 19363
rect 8159 19329 8168 19363
rect 8116 19320 8168 19329
rect 8024 19252 8076 19304
rect 3424 19184 3476 19236
rect 3884 19227 3936 19236
rect 3884 19193 3893 19227
rect 3893 19193 3927 19227
rect 3927 19193 3936 19227
rect 3884 19184 3936 19193
rect 10048 19363 10100 19372
rect 10048 19329 10057 19363
rect 10057 19329 10091 19363
rect 10091 19329 10100 19363
rect 10048 19320 10100 19329
rect 10784 19252 10836 19304
rect 11520 19252 11572 19304
rect 12256 19252 12308 19304
rect 8760 19184 8812 19236
rect 10508 19184 10560 19236
rect 4160 19116 4212 19168
rect 5632 19159 5684 19168
rect 5632 19125 5641 19159
rect 5641 19125 5675 19159
rect 5675 19125 5684 19159
rect 5632 19116 5684 19125
rect 5724 19116 5776 19168
rect 7564 19116 7616 19168
rect 9312 19116 9364 19168
rect 9772 19159 9824 19168
rect 9772 19125 9781 19159
rect 9781 19125 9815 19159
rect 9815 19125 9824 19159
rect 9772 19116 9824 19125
rect 11428 19184 11480 19236
rect 12624 19184 12676 19236
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 1676 18912 1728 18964
rect 5632 18912 5684 18964
rect 8116 18912 8168 18964
rect 2228 18844 2280 18896
rect 2320 18776 2372 18828
rect 3056 18844 3108 18896
rect 4528 18844 4580 18896
rect 1952 18751 2004 18760
rect 1952 18717 1961 18751
rect 1961 18717 1995 18751
rect 1995 18717 2004 18751
rect 1952 18708 2004 18717
rect 2780 18776 2832 18828
rect 6184 18819 6236 18828
rect 6184 18785 6193 18819
rect 6193 18785 6227 18819
rect 6227 18785 6236 18819
rect 6184 18776 6236 18785
rect 6736 18819 6788 18828
rect 6736 18785 6745 18819
rect 6745 18785 6779 18819
rect 6779 18785 6788 18819
rect 6736 18776 6788 18785
rect 8484 18776 8536 18828
rect 10508 18912 10560 18964
rect 8760 18819 8812 18828
rect 8760 18785 8769 18819
rect 8769 18785 8803 18819
rect 8803 18785 8812 18819
rect 8760 18776 8812 18785
rect 9404 18776 9456 18828
rect 10968 18844 11020 18896
rect 11428 18887 11480 18896
rect 11428 18853 11437 18887
rect 11437 18853 11471 18887
rect 11471 18853 11480 18887
rect 11428 18844 11480 18853
rect 9772 18776 9824 18828
rect 13268 18776 13320 18828
rect 2964 18751 3016 18760
rect 2044 18572 2096 18624
rect 2964 18717 2973 18751
rect 2973 18717 3007 18751
rect 3007 18717 3016 18751
rect 2964 18708 3016 18717
rect 3976 18708 4028 18760
rect 4712 18708 4764 18760
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 8760 18640 8812 18692
rect 10876 18708 10928 18760
rect 10416 18640 10468 18692
rect 11520 18640 11572 18692
rect 8852 18572 8904 18624
rect 11336 18572 11388 18624
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 2412 18368 2464 18420
rect 4160 18411 4212 18420
rect 4160 18377 4169 18411
rect 4169 18377 4203 18411
rect 4203 18377 4212 18411
rect 4160 18368 4212 18377
rect 4804 18368 4856 18420
rect 6184 18368 6236 18420
rect 10876 18368 10928 18420
rect 13268 18411 13320 18420
rect 13268 18377 13277 18411
rect 13277 18377 13311 18411
rect 13311 18377 13320 18411
rect 13268 18368 13320 18377
rect 1768 18300 1820 18352
rect 5540 18300 5592 18352
rect 6736 18300 6788 18352
rect 7472 18300 7524 18352
rect 8392 18300 8444 18352
rect 11428 18300 11480 18352
rect 2964 18232 3016 18284
rect 4712 18232 4764 18284
rect 1952 18164 2004 18216
rect 6184 18164 6236 18216
rect 8116 18232 8168 18284
rect 8852 18232 8904 18284
rect 10692 18232 10744 18284
rect 12072 18232 12124 18284
rect 4712 18139 4764 18148
rect 4712 18105 4721 18139
rect 4721 18105 4755 18139
rect 4755 18105 4764 18139
rect 4712 18096 4764 18105
rect 4804 18139 4856 18148
rect 4804 18105 4813 18139
rect 4813 18105 4847 18139
rect 4847 18105 4856 18139
rect 9772 18164 9824 18216
rect 4804 18096 4856 18105
rect 1952 18028 2004 18080
rect 2228 18028 2280 18080
rect 2780 18071 2832 18080
rect 2780 18037 2789 18071
rect 2789 18037 2823 18071
rect 2823 18037 2832 18071
rect 2780 18028 2832 18037
rect 4528 18071 4580 18080
rect 4528 18037 4537 18071
rect 4537 18037 4571 18071
rect 4571 18037 4580 18071
rect 4528 18028 4580 18037
rect 8392 18096 8444 18148
rect 9312 18096 9364 18148
rect 9864 18096 9916 18148
rect 10876 18164 10928 18216
rect 10968 18207 11020 18216
rect 10968 18173 10977 18207
rect 10977 18173 11011 18207
rect 11011 18173 11020 18207
rect 10968 18164 11020 18173
rect 12348 18164 12400 18216
rect 13912 18232 13964 18284
rect 8208 18028 8260 18080
rect 9404 18028 9456 18080
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 9772 18028 9824 18080
rect 12072 18096 12124 18148
rect 13360 18028 13412 18080
rect 13912 18071 13964 18080
rect 13912 18037 13921 18071
rect 13921 18037 13955 18071
rect 13955 18037 13964 18071
rect 13912 18028 13964 18037
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 2964 17824 3016 17876
rect 4344 17824 4396 17876
rect 2688 17756 2740 17808
rect 4528 17824 4580 17876
rect 8484 17867 8536 17876
rect 4620 17756 4672 17808
rect 8484 17833 8493 17867
rect 8493 17833 8527 17867
rect 8527 17833 8536 17867
rect 8484 17824 8536 17833
rect 9588 17824 9640 17876
rect 6000 17799 6052 17808
rect 6000 17765 6009 17799
rect 6009 17765 6043 17799
rect 6043 17765 6052 17799
rect 6000 17756 6052 17765
rect 8116 17799 8168 17808
rect 8116 17765 8125 17799
rect 8125 17765 8159 17799
rect 8159 17765 8168 17799
rect 8116 17756 8168 17765
rect 8392 17756 8444 17808
rect 9496 17756 9548 17808
rect 9864 17799 9916 17808
rect 9864 17765 9873 17799
rect 9873 17765 9907 17799
rect 9907 17765 9916 17799
rect 9864 17756 9916 17765
rect 11336 17799 11388 17808
rect 11336 17765 11345 17799
rect 11345 17765 11379 17799
rect 11379 17765 11388 17799
rect 11336 17756 11388 17765
rect 11428 17799 11480 17808
rect 11428 17765 11437 17799
rect 11437 17765 11471 17799
rect 11471 17765 11480 17799
rect 11428 17756 11480 17765
rect 3424 17688 3476 17740
rect 7380 17731 7432 17740
rect 7380 17697 7389 17731
rect 7389 17697 7423 17731
rect 7423 17697 7432 17731
rect 7380 17688 7432 17697
rect 7840 17688 7892 17740
rect 9588 17688 9640 17740
rect 10416 17731 10468 17740
rect 10416 17697 10425 17731
rect 10425 17697 10459 17731
rect 10459 17697 10468 17731
rect 10416 17688 10468 17697
rect 13268 17688 13320 17740
rect 2044 17663 2096 17672
rect 2044 17629 2053 17663
rect 2053 17629 2087 17663
rect 2087 17629 2096 17663
rect 2044 17620 2096 17629
rect 2320 17620 2372 17672
rect 5632 17620 5684 17672
rect 6184 17663 6236 17672
rect 6184 17629 6193 17663
rect 6193 17629 6227 17663
rect 6227 17629 6236 17663
rect 6184 17620 6236 17629
rect 7564 17620 7616 17672
rect 10048 17620 10100 17672
rect 13360 17620 13412 17672
rect 1952 17484 2004 17536
rect 2320 17484 2372 17536
rect 10876 17552 10928 17604
rect 4712 17484 4764 17536
rect 7380 17484 7432 17536
rect 9312 17484 9364 17536
rect 10784 17484 10836 17536
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 5724 17280 5776 17332
rect 6000 17323 6052 17332
rect 6000 17289 6009 17323
rect 6009 17289 6043 17323
rect 6043 17289 6052 17323
rect 6000 17280 6052 17289
rect 9864 17323 9916 17332
rect 9864 17289 9873 17323
rect 9873 17289 9907 17323
rect 9907 17289 9916 17323
rect 9864 17280 9916 17289
rect 10048 17280 10100 17332
rect 11336 17280 11388 17332
rect 13268 17323 13320 17332
rect 13268 17289 13277 17323
rect 13277 17289 13311 17323
rect 13311 17289 13320 17323
rect 13268 17280 13320 17289
rect 6644 17212 6696 17264
rect 6736 17144 6788 17196
rect 8024 17187 8076 17196
rect 8024 17153 8033 17187
rect 8033 17153 8067 17187
rect 8067 17153 8076 17187
rect 8024 17144 8076 17153
rect 9220 17144 9272 17196
rect 10692 17144 10744 17196
rect 11428 17144 11480 17196
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 3148 17076 3200 17128
rect 4804 17119 4856 17128
rect 4804 17085 4813 17119
rect 4813 17085 4847 17119
rect 4847 17085 4856 17119
rect 4804 17076 4856 17085
rect 5816 17076 5868 17128
rect 6828 17076 6880 17128
rect 7564 17119 7616 17128
rect 7564 17085 7573 17119
rect 7573 17085 7607 17119
rect 7607 17085 7616 17119
rect 7564 17076 7616 17085
rect 7840 17119 7892 17128
rect 7840 17085 7849 17119
rect 7849 17085 7883 17119
rect 7883 17085 7892 17119
rect 7840 17076 7892 17085
rect 8668 17076 8720 17128
rect 9312 17076 9364 17128
rect 9956 17076 10008 17128
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 12164 17076 12216 17128
rect 12900 17119 12952 17128
rect 12900 17085 12909 17119
rect 12909 17085 12943 17119
rect 12943 17085 12952 17119
rect 12900 17076 12952 17085
rect 13728 17076 13780 17128
rect 2136 17008 2188 17060
rect 2780 17051 2832 17060
rect 2780 17017 2789 17051
rect 2789 17017 2823 17051
rect 2823 17017 2832 17051
rect 2780 17008 2832 17017
rect 4344 17008 4396 17060
rect 5540 17008 5592 17060
rect 1676 16983 1728 16992
rect 1676 16949 1685 16983
rect 1685 16949 1719 16983
rect 1719 16949 1728 16983
rect 1676 16940 1728 16949
rect 1860 16940 1912 16992
rect 3884 16983 3936 16992
rect 3884 16949 3893 16983
rect 3893 16949 3927 16983
rect 3927 16949 3936 16983
rect 3884 16940 3936 16949
rect 5724 16983 5776 16992
rect 5724 16949 5733 16983
rect 5733 16949 5767 16983
rect 5767 16949 5776 16983
rect 5724 16940 5776 16949
rect 7564 16940 7616 16992
rect 8392 16983 8444 16992
rect 8392 16949 8401 16983
rect 8401 16949 8435 16983
rect 8435 16949 8444 16983
rect 8392 16940 8444 16949
rect 8852 16940 8904 16992
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 2688 16736 2740 16788
rect 3424 16736 3476 16788
rect 4804 16736 4856 16788
rect 7380 16736 7432 16788
rect 2136 16668 2188 16720
rect 3884 16668 3936 16720
rect 4252 16711 4304 16720
rect 4252 16677 4261 16711
rect 4261 16677 4295 16711
rect 4295 16677 4304 16711
rect 4252 16668 4304 16677
rect 5540 16711 5592 16720
rect 5540 16677 5549 16711
rect 5549 16677 5583 16711
rect 5583 16677 5592 16711
rect 5540 16668 5592 16677
rect 5724 16668 5776 16720
rect 7472 16668 7524 16720
rect 10968 16668 11020 16720
rect 11520 16668 11572 16720
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 7196 16643 7248 16652
rect 7196 16609 7205 16643
rect 7205 16609 7239 16643
rect 7239 16609 7248 16643
rect 7196 16600 7248 16609
rect 8208 16600 8260 16652
rect 9680 16643 9732 16652
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 11244 16643 11296 16652
rect 11244 16609 11253 16643
rect 11253 16609 11287 16643
rect 11287 16609 11296 16643
rect 11244 16600 11296 16609
rect 12624 16600 12676 16652
rect 3976 16532 4028 16584
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 6000 16532 6052 16584
rect 6184 16575 6236 16584
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 6184 16532 6236 16541
rect 6736 16532 6788 16584
rect 10876 16532 10928 16584
rect 13176 16532 13228 16584
rect 8668 16464 8720 16516
rect 9312 16464 9364 16516
rect 9864 16464 9916 16516
rect 3056 16439 3108 16448
rect 3056 16405 3065 16439
rect 3065 16405 3099 16439
rect 3099 16405 3108 16439
rect 3056 16396 3108 16405
rect 3148 16396 3200 16448
rect 6828 16439 6880 16448
rect 6828 16405 6837 16439
rect 6837 16405 6871 16439
rect 6871 16405 6880 16439
rect 6828 16396 6880 16405
rect 9588 16396 9640 16448
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 2044 16192 2096 16244
rect 4252 16235 4304 16244
rect 4252 16201 4261 16235
rect 4261 16201 4295 16235
rect 4295 16201 4304 16235
rect 4252 16192 4304 16201
rect 4988 16192 5040 16244
rect 5724 16192 5776 16244
rect 6000 16192 6052 16244
rect 6644 16192 6696 16244
rect 7196 16192 7248 16244
rect 7656 16192 7708 16244
rect 9956 16192 10008 16244
rect 10968 16192 11020 16244
rect 12624 16235 12676 16244
rect 12624 16201 12633 16235
rect 12633 16201 12667 16235
rect 12667 16201 12676 16235
rect 12624 16192 12676 16201
rect 3240 16124 3292 16176
rect 1308 16056 1360 16108
rect 4896 16056 4948 16108
rect 5908 16056 5960 16108
rect 9220 16099 9272 16108
rect 9220 16065 9229 16099
rect 9229 16065 9263 16099
rect 9263 16065 9272 16099
rect 9220 16056 9272 16065
rect 9588 16056 9640 16108
rect 9680 16056 9732 16108
rect 2320 15988 2372 16040
rect 3056 15988 3108 16040
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 6920 16031 6972 16040
rect 6920 15997 6929 16031
rect 6929 15997 6963 16031
rect 6963 15997 6972 16031
rect 6920 15988 6972 15997
rect 2136 15920 2188 15972
rect 4252 15920 4304 15972
rect 3884 15895 3936 15904
rect 3884 15861 3893 15895
rect 3893 15861 3927 15895
rect 3927 15861 3936 15895
rect 3884 15852 3936 15861
rect 4988 15963 5040 15972
rect 4988 15929 4997 15963
rect 4997 15929 5031 15963
rect 5031 15929 5040 15963
rect 4988 15920 5040 15929
rect 7564 15988 7616 16040
rect 9496 15963 9548 15972
rect 9496 15929 9505 15963
rect 9505 15929 9539 15963
rect 9539 15929 9548 15963
rect 9496 15920 9548 15929
rect 10232 15920 10284 15972
rect 10692 15920 10744 15972
rect 11244 15920 11296 15972
rect 5540 15852 5592 15904
rect 8208 15895 8260 15904
rect 8208 15861 8217 15895
rect 8217 15861 8251 15895
rect 8251 15861 8260 15895
rect 8208 15852 8260 15861
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 1676 15648 1728 15700
rect 3976 15648 4028 15700
rect 4068 15648 4120 15700
rect 5264 15691 5316 15700
rect 5264 15657 5273 15691
rect 5273 15657 5307 15691
rect 5307 15657 5316 15691
rect 5264 15648 5316 15657
rect 9588 15648 9640 15700
rect 2044 15580 2096 15632
rect 3148 15623 3200 15632
rect 3148 15589 3157 15623
rect 3157 15589 3191 15623
rect 3191 15589 3200 15623
rect 3148 15580 3200 15589
rect 3884 15580 3936 15632
rect 4620 15580 4672 15632
rect 4804 15623 4856 15632
rect 4804 15589 4813 15623
rect 4813 15589 4847 15623
rect 4847 15589 4856 15623
rect 4804 15580 4856 15589
rect 2412 15555 2464 15564
rect 2412 15521 2421 15555
rect 2421 15521 2455 15555
rect 2455 15521 2464 15555
rect 2412 15512 2464 15521
rect 2964 15555 3016 15564
rect 2964 15521 2973 15555
rect 2973 15521 3007 15555
rect 3007 15521 3016 15555
rect 2964 15512 3016 15521
rect 6276 15512 6328 15564
rect 9220 15580 9272 15632
rect 9496 15580 9548 15632
rect 9864 15623 9916 15632
rect 9864 15589 9873 15623
rect 9873 15589 9907 15623
rect 9907 15589 9916 15623
rect 9864 15580 9916 15589
rect 9956 15580 10008 15632
rect 4896 15444 4948 15496
rect 2320 15419 2372 15428
rect 2320 15385 2329 15419
rect 2329 15385 2363 15419
rect 2363 15385 2372 15419
rect 2320 15376 2372 15385
rect 4068 15376 4120 15428
rect 7564 15555 7616 15564
rect 7564 15521 7573 15555
rect 7573 15521 7607 15555
rect 7607 15521 7616 15555
rect 11428 15555 11480 15564
rect 7564 15512 7616 15521
rect 11428 15521 11437 15555
rect 11437 15521 11471 15555
rect 11471 15521 11480 15555
rect 11428 15512 11480 15521
rect 12440 15512 12492 15564
rect 13452 15512 13504 15564
rect 7748 15487 7800 15496
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 9956 15444 10008 15496
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 6920 15419 6972 15428
rect 6920 15385 6929 15419
rect 6929 15385 6963 15419
rect 6963 15385 6972 15419
rect 7380 15419 7432 15428
rect 6920 15376 6972 15385
rect 7380 15385 7389 15419
rect 7389 15385 7423 15419
rect 7423 15385 7432 15419
rect 7380 15376 7432 15385
rect 7472 15376 7524 15428
rect 8116 15376 8168 15428
rect 9680 15376 9732 15428
rect 8300 15351 8352 15360
rect 8300 15317 8309 15351
rect 8309 15317 8343 15351
rect 8343 15317 8352 15351
rect 8300 15308 8352 15317
rect 8760 15351 8812 15360
rect 8760 15317 8769 15351
rect 8769 15317 8803 15351
rect 8803 15317 8812 15351
rect 8760 15308 8812 15317
rect 11336 15308 11388 15360
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 1952 15104 2004 15156
rect 2964 15104 3016 15156
rect 6736 15104 6788 15156
rect 7472 15104 7524 15156
rect 7564 15104 7616 15156
rect 1584 15036 1636 15088
rect 2412 15079 2464 15088
rect 1584 14900 1636 14952
rect 2412 15045 2421 15079
rect 2421 15045 2455 15079
rect 2455 15045 2464 15079
rect 2412 15036 2464 15045
rect 3056 15011 3108 15020
rect 3056 14977 3065 15011
rect 3065 14977 3099 15011
rect 3099 14977 3108 15011
rect 3056 14968 3108 14977
rect 2780 14900 2832 14952
rect 2964 14943 3016 14952
rect 2964 14909 2973 14943
rect 2973 14909 3007 14943
rect 3007 14909 3016 14943
rect 8208 15036 8260 15088
rect 9864 15104 9916 15156
rect 11428 15104 11480 15156
rect 6276 15011 6328 15020
rect 6276 14977 6285 15011
rect 6285 14977 6319 15011
rect 6319 14977 6328 15011
rect 6276 14968 6328 14977
rect 8760 14968 8812 15020
rect 2964 14900 3016 14909
rect 5264 14900 5316 14952
rect 5724 14943 5776 14952
rect 5724 14909 5733 14943
rect 5733 14909 5767 14943
rect 5767 14909 5776 14943
rect 5724 14900 5776 14909
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 5908 14900 5960 14909
rect 7748 14900 7800 14952
rect 9772 14943 9824 14952
rect 9772 14909 9781 14943
rect 9781 14909 9815 14943
rect 9815 14909 9824 14943
rect 9772 14900 9824 14909
rect 11520 14900 11572 14952
rect 12716 14900 12768 14952
rect 7932 14832 7984 14884
rect 4436 14764 4488 14816
rect 5724 14764 5776 14816
rect 8300 14764 8352 14816
rect 8944 14807 8996 14816
rect 8944 14773 8953 14807
rect 8953 14773 8987 14807
rect 8987 14773 8996 14807
rect 8944 14764 8996 14773
rect 11336 14764 11388 14816
rect 13452 14807 13504 14816
rect 13452 14773 13461 14807
rect 13461 14773 13495 14807
rect 13495 14773 13504 14807
rect 13452 14764 13504 14773
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 4620 14603 4672 14612
rect 4620 14569 4629 14603
rect 4629 14569 4663 14603
rect 4663 14569 4672 14603
rect 4620 14560 4672 14569
rect 7380 14603 7432 14612
rect 7380 14569 7389 14603
rect 7389 14569 7423 14603
rect 7423 14569 7432 14603
rect 7380 14560 7432 14569
rect 9772 14560 9824 14612
rect 4344 14492 4396 14544
rect 4988 14535 5040 14544
rect 4988 14501 4997 14535
rect 4997 14501 5031 14535
rect 5031 14501 5040 14535
rect 4988 14492 5040 14501
rect 6184 14492 6236 14544
rect 1768 14424 1820 14476
rect 2412 14467 2464 14476
rect 2412 14433 2421 14467
rect 2421 14433 2455 14467
rect 2455 14433 2464 14467
rect 2412 14424 2464 14433
rect 2688 14467 2740 14476
rect 2688 14433 2697 14467
rect 2697 14433 2731 14467
rect 2731 14433 2740 14467
rect 2688 14424 2740 14433
rect 3240 14424 3292 14476
rect 6368 14467 6420 14476
rect 6368 14433 6377 14467
rect 6377 14433 6411 14467
rect 6411 14433 6420 14467
rect 6368 14424 6420 14433
rect 7012 14492 7064 14544
rect 6552 14424 6604 14476
rect 7564 14424 7616 14476
rect 7932 14467 7984 14476
rect 7932 14433 7941 14467
rect 7941 14433 7975 14467
rect 7975 14433 7984 14467
rect 7932 14424 7984 14433
rect 8668 14492 8720 14544
rect 8944 14492 8996 14544
rect 9588 14492 9640 14544
rect 10416 14535 10468 14544
rect 10416 14501 10425 14535
rect 10425 14501 10459 14535
rect 10459 14501 10468 14535
rect 10416 14492 10468 14501
rect 10968 14492 11020 14544
rect 12716 14492 12768 14544
rect 11520 14467 11572 14476
rect 11520 14433 11529 14467
rect 11529 14433 11563 14467
rect 11563 14433 11572 14467
rect 11520 14424 11572 14433
rect 11704 14467 11756 14476
rect 11704 14433 11713 14467
rect 11713 14433 11747 14467
rect 11747 14433 11756 14467
rect 11704 14424 11756 14433
rect 13268 14424 13320 14476
rect 1584 14356 1636 14408
rect 4712 14356 4764 14408
rect 4896 14399 4948 14408
rect 4896 14365 4905 14399
rect 4905 14365 4939 14399
rect 4939 14365 4948 14399
rect 4896 14356 4948 14365
rect 3148 14288 3200 14340
rect 8392 14356 8444 14408
rect 8668 14399 8720 14408
rect 8668 14365 8677 14399
rect 8677 14365 8711 14399
rect 8711 14365 8720 14399
rect 8668 14356 8720 14365
rect 2320 14263 2372 14272
rect 2320 14229 2329 14263
rect 2329 14229 2363 14263
rect 2363 14229 2372 14263
rect 6184 14288 6236 14340
rect 7564 14288 7616 14340
rect 8576 14288 8628 14340
rect 9680 14288 9732 14340
rect 3424 14263 3476 14272
rect 2320 14220 2372 14229
rect 3424 14229 3433 14263
rect 3433 14229 3467 14263
rect 3467 14229 3476 14263
rect 3424 14220 3476 14229
rect 4436 14220 4488 14272
rect 6828 14220 6880 14272
rect 8484 14220 8536 14272
rect 9956 14220 10008 14272
rect 11612 14220 11664 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 2688 14016 2740 14068
rect 4804 14016 4856 14068
rect 4988 14016 5040 14068
rect 6092 14016 6144 14068
rect 6368 14016 6420 14068
rect 7472 14016 7524 14068
rect 7748 14016 7800 14068
rect 7932 14016 7984 14068
rect 9588 14059 9640 14068
rect 9588 14025 9597 14059
rect 9597 14025 9631 14059
rect 9631 14025 9640 14059
rect 9864 14059 9916 14068
rect 9588 14016 9640 14025
rect 9864 14025 9873 14059
rect 9873 14025 9907 14059
rect 9907 14025 9916 14059
rect 9864 14016 9916 14025
rect 11152 14016 11204 14068
rect 11520 14016 11572 14068
rect 11612 14016 11664 14068
rect 13268 14059 13320 14068
rect 13268 14025 13277 14059
rect 13277 14025 13311 14059
rect 13311 14025 13320 14059
rect 13268 14016 13320 14025
rect 2412 13948 2464 14000
rect 6828 13948 6880 14000
rect 6920 13948 6972 14000
rect 8852 13948 8904 14000
rect 2228 13880 2280 13932
rect 2504 13880 2556 13932
rect 4344 13923 4396 13932
rect 2320 13812 2372 13864
rect 2412 13812 2464 13864
rect 4344 13889 4353 13923
rect 4353 13889 4387 13923
rect 4387 13889 4396 13923
rect 4344 13880 4396 13889
rect 4804 13880 4856 13932
rect 5908 13880 5960 13932
rect 8760 13880 8812 13932
rect 3056 13812 3108 13864
rect 2872 13744 2924 13796
rect 3424 13812 3476 13864
rect 5540 13812 5592 13864
rect 6552 13812 6604 13864
rect 4436 13787 4488 13796
rect 4436 13753 4445 13787
rect 4445 13753 4479 13787
rect 4479 13753 4488 13787
rect 4436 13744 4488 13753
rect 5632 13744 5684 13796
rect 6092 13744 6144 13796
rect 7932 13744 7984 13796
rect 8300 13744 8352 13796
rect 10232 13880 10284 13932
rect 10416 13923 10468 13932
rect 10416 13889 10425 13923
rect 10425 13889 10459 13923
rect 10459 13889 10468 13923
rect 10416 13880 10468 13889
rect 11336 13880 11388 13932
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 12900 13880 12952 13932
rect 9956 13744 10008 13796
rect 10140 13787 10192 13796
rect 10140 13753 10149 13787
rect 10149 13753 10183 13787
rect 10183 13753 10192 13787
rect 10140 13744 10192 13753
rect 1860 13719 1912 13728
rect 1860 13685 1869 13719
rect 1869 13685 1903 13719
rect 1903 13685 1912 13719
rect 1860 13676 1912 13685
rect 2964 13719 3016 13728
rect 2964 13685 2973 13719
rect 2973 13685 3007 13719
rect 3007 13685 3016 13719
rect 2964 13676 3016 13685
rect 3148 13676 3200 13728
rect 6000 13676 6052 13728
rect 8024 13676 8076 13728
rect 9864 13676 9916 13728
rect 13084 13744 13136 13796
rect 10600 13676 10652 13728
rect 11336 13676 11388 13728
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 12992 13676 13044 13728
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 1860 13472 1912 13524
rect 4344 13472 4396 13524
rect 7472 13515 7524 13524
rect 3056 13404 3108 13456
rect 5724 13404 5776 13456
rect 6092 13404 6144 13456
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 8760 13515 8812 13524
rect 8760 13481 8769 13515
rect 8769 13481 8803 13515
rect 8803 13481 8812 13515
rect 8760 13472 8812 13481
rect 9680 13472 9732 13524
rect 10140 13472 10192 13524
rect 12992 13472 13044 13524
rect 8392 13447 8444 13456
rect 8392 13413 8401 13447
rect 8401 13413 8435 13447
rect 8435 13413 8444 13447
rect 8392 13404 8444 13413
rect 9864 13447 9916 13456
rect 9864 13413 9873 13447
rect 9873 13413 9907 13447
rect 9907 13413 9916 13447
rect 9864 13404 9916 13413
rect 9956 13404 10008 13456
rect 11796 13404 11848 13456
rect 2688 13379 2740 13388
rect 2688 13345 2697 13379
rect 2697 13345 2731 13379
rect 2731 13345 2740 13379
rect 2688 13336 2740 13345
rect 2872 13379 2924 13388
rect 2872 13345 2881 13379
rect 2881 13345 2915 13379
rect 2915 13345 2924 13379
rect 2872 13336 2924 13345
rect 6828 13336 6880 13388
rect 7656 13336 7708 13388
rect 7840 13379 7892 13388
rect 7840 13345 7849 13379
rect 7849 13345 7883 13379
rect 7883 13345 7892 13379
rect 7840 13336 7892 13345
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 3976 13268 4028 13320
rect 4896 13268 4948 13320
rect 5356 13268 5408 13320
rect 6644 13268 6696 13320
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 11336 13311 11388 13320
rect 10416 13268 10468 13277
rect 11336 13277 11345 13311
rect 11345 13277 11379 13311
rect 11379 13277 11388 13311
rect 11336 13268 11388 13277
rect 11428 13268 11480 13320
rect 11980 13268 12032 13320
rect 12348 13268 12400 13320
rect 3240 13200 3292 13252
rect 4436 13200 4488 13252
rect 6000 13200 6052 13252
rect 6736 13200 6788 13252
rect 10232 13200 10284 13252
rect 1768 13132 1820 13184
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2320 13132 2372 13141
rect 5356 13175 5408 13184
rect 5356 13141 5365 13175
rect 5365 13141 5399 13175
rect 5399 13141 5408 13175
rect 5356 13132 5408 13141
rect 11980 13132 12032 13184
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 8668 12928 8720 12980
rect 9772 12928 9824 12980
rect 13912 12971 13964 12980
rect 13912 12937 13921 12971
rect 13921 12937 13955 12971
rect 13955 12937 13964 12971
rect 13912 12928 13964 12937
rect 5356 12792 5408 12844
rect 7472 12792 7524 12844
rect 11796 12860 11848 12912
rect 2320 12724 2372 12776
rect 2872 12724 2924 12776
rect 3148 12724 3200 12776
rect 2228 12699 2280 12708
rect 2228 12665 2237 12699
rect 2237 12665 2271 12699
rect 2271 12665 2280 12699
rect 2228 12656 2280 12665
rect 2412 12588 2464 12640
rect 2780 12588 2832 12640
rect 4436 12656 4488 12708
rect 6644 12699 6696 12708
rect 6644 12665 6653 12699
rect 6653 12665 6687 12699
rect 6687 12665 6696 12699
rect 6644 12656 6696 12665
rect 4068 12588 4120 12640
rect 5724 12588 5776 12640
rect 6828 12588 6880 12640
rect 7932 12656 7984 12708
rect 10968 12724 11020 12776
rect 12072 12724 12124 12776
rect 12164 12724 12216 12776
rect 12900 12767 12952 12776
rect 12900 12733 12909 12767
rect 12909 12733 12943 12767
rect 12943 12733 12952 12767
rect 12900 12724 12952 12733
rect 13728 12724 13780 12776
rect 13912 12724 13964 12776
rect 10232 12699 10284 12708
rect 10232 12665 10241 12699
rect 10241 12665 10275 12699
rect 10275 12665 10284 12699
rect 10232 12656 10284 12665
rect 9864 12588 9916 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 2688 12384 2740 12436
rect 3976 12384 4028 12436
rect 4436 12427 4488 12436
rect 4436 12393 4445 12427
rect 4445 12393 4479 12427
rect 4479 12393 4488 12427
rect 4436 12384 4488 12393
rect 4988 12427 5040 12436
rect 4988 12393 4997 12427
rect 4997 12393 5031 12427
rect 5031 12393 5040 12427
rect 4988 12384 5040 12393
rect 5356 12427 5408 12436
rect 5356 12393 5365 12427
rect 5365 12393 5399 12427
rect 5399 12393 5408 12427
rect 5356 12384 5408 12393
rect 9404 12384 9456 12436
rect 3332 12316 3384 12368
rect 6000 12359 6052 12368
rect 6000 12325 6009 12359
rect 6009 12325 6043 12359
rect 6043 12325 6052 12359
rect 6000 12316 6052 12325
rect 7932 12316 7984 12368
rect 9772 12316 9824 12368
rect 11336 12384 11388 12436
rect 11980 12384 12032 12436
rect 10416 12359 10468 12368
rect 10416 12325 10425 12359
rect 10425 12325 10459 12359
rect 10459 12325 10468 12359
rect 10416 12316 10468 12325
rect 11428 12316 11480 12368
rect 1492 12248 1544 12300
rect 1768 12248 1820 12300
rect 2228 12248 2280 12300
rect 4252 12248 4304 12300
rect 10876 12248 10928 12300
rect 1860 12180 1912 12232
rect 2872 12180 2924 12232
rect 6184 12223 6236 12232
rect 1768 12112 1820 12164
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 6920 12180 6972 12232
rect 7748 12180 7800 12232
rect 9588 12180 9640 12232
rect 10232 12180 10284 12232
rect 12072 12180 12124 12232
rect 6092 12112 6144 12164
rect 2320 12044 2372 12096
rect 7840 12044 7892 12096
rect 9864 12044 9916 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 1584 11840 1636 11892
rect 2044 11840 2096 11892
rect 3332 11840 3384 11892
rect 4436 11883 4488 11892
rect 4436 11849 4445 11883
rect 4445 11849 4479 11883
rect 4479 11849 4488 11883
rect 4436 11840 4488 11849
rect 4988 11840 5040 11892
rect 6000 11883 6052 11892
rect 6000 11849 6009 11883
rect 6009 11849 6043 11883
rect 6043 11849 6052 11883
rect 6000 11840 6052 11849
rect 8484 11840 8536 11892
rect 9496 11883 9548 11892
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 12072 11840 12124 11892
rect 13084 11840 13136 11892
rect 1400 11704 1452 11756
rect 2964 11704 3016 11756
rect 5172 11704 5224 11756
rect 6092 11704 6144 11756
rect 4436 11636 4488 11688
rect 5632 11679 5684 11688
rect 5632 11645 5641 11679
rect 5641 11645 5675 11679
rect 5675 11645 5684 11679
rect 5632 11636 5684 11645
rect 2136 11568 2188 11620
rect 5080 11611 5132 11620
rect 5080 11577 5089 11611
rect 5089 11577 5123 11611
rect 5123 11577 5132 11611
rect 5080 11568 5132 11577
rect 3332 11500 3384 11552
rect 3976 11500 4028 11552
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 7196 11747 7248 11756
rect 7196 11713 7205 11747
rect 7205 11713 7239 11747
rect 7239 11713 7248 11747
rect 7196 11704 7248 11713
rect 8668 11704 8720 11756
rect 8116 11636 8168 11688
rect 12072 11636 12124 11688
rect 13452 11636 13504 11688
rect 7656 11568 7708 11620
rect 7932 11543 7984 11552
rect 7932 11509 7941 11543
rect 7941 11509 7975 11543
rect 7975 11509 7984 11543
rect 7932 11500 7984 11509
rect 8116 11500 8168 11552
rect 9496 11500 9548 11552
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 10876 11500 10928 11552
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 1768 11296 1820 11348
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 2964 11296 3016 11348
rect 4252 11339 4304 11348
rect 4252 11305 4261 11339
rect 4261 11305 4295 11339
rect 4295 11305 4304 11339
rect 4252 11296 4304 11305
rect 5172 11296 5224 11348
rect 9404 11339 9456 11348
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 9772 11339 9824 11348
rect 9772 11305 9781 11339
rect 9781 11305 9815 11339
rect 9815 11305 9824 11339
rect 9772 11296 9824 11305
rect 9864 11296 9916 11348
rect 3148 11271 3200 11280
rect 3148 11237 3157 11271
rect 3157 11237 3191 11271
rect 3191 11237 3200 11271
rect 3148 11228 3200 11237
rect 5724 11271 5776 11280
rect 5724 11237 5733 11271
rect 5733 11237 5767 11271
rect 5767 11237 5776 11271
rect 5724 11228 5776 11237
rect 6920 11228 6972 11280
rect 7932 11228 7984 11280
rect 8392 11228 8444 11280
rect 9588 11228 9640 11280
rect 1952 11160 2004 11212
rect 2504 11203 2556 11212
rect 2504 11169 2513 11203
rect 2513 11169 2547 11203
rect 2547 11169 2556 11203
rect 2504 11160 2556 11169
rect 2872 11203 2924 11212
rect 2872 11169 2881 11203
rect 2881 11169 2915 11203
rect 2915 11169 2924 11203
rect 2872 11160 2924 11169
rect 5264 11160 5316 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 1860 11092 1912 11144
rect 6000 11092 6052 11144
rect 7656 11092 7708 11144
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 9496 11092 9548 11144
rect 11060 11160 11112 11212
rect 11152 11092 11204 11144
rect 2964 11024 3016 11076
rect 7380 11024 7432 11076
rect 7748 11067 7800 11076
rect 7748 11033 7757 11067
rect 7757 11033 7791 11067
rect 7791 11033 7800 11067
rect 7748 11024 7800 11033
rect 10048 11024 10100 11076
rect 3332 10956 3384 11008
rect 6828 10956 6880 11008
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 2504 10752 2556 10804
rect 4068 10752 4120 10804
rect 5724 10752 5776 10804
rect 7932 10752 7984 10804
rect 9956 10752 10008 10804
rect 10784 10752 10836 10804
rect 4896 10684 4948 10736
rect 8300 10684 8352 10736
rect 10692 10684 10744 10736
rect 3976 10616 4028 10668
rect 4436 10659 4488 10668
rect 4436 10625 4445 10659
rect 4445 10625 4479 10659
rect 4479 10625 4488 10659
rect 4436 10616 4488 10625
rect 7840 10616 7892 10668
rect 8668 10616 8720 10668
rect 1584 10548 1636 10600
rect 2228 10591 2280 10600
rect 2228 10557 2237 10591
rect 2237 10557 2271 10591
rect 2271 10557 2280 10591
rect 2228 10548 2280 10557
rect 2872 10548 2924 10600
rect 1952 10480 2004 10532
rect 6828 10591 6880 10600
rect 4252 10523 4304 10532
rect 4252 10489 4261 10523
rect 4261 10489 4295 10523
rect 4295 10489 4304 10523
rect 4252 10480 4304 10489
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 7380 10548 7432 10600
rect 8484 10548 8536 10600
rect 8760 10548 8812 10600
rect 10140 10548 10192 10600
rect 9956 10523 10008 10532
rect 9956 10489 9965 10523
rect 9965 10489 9999 10523
rect 9999 10489 10008 10523
rect 9956 10480 10008 10489
rect 1860 10455 1912 10464
rect 1860 10421 1869 10455
rect 1869 10421 1903 10455
rect 1903 10421 1912 10455
rect 1860 10412 1912 10421
rect 5264 10412 5316 10464
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 7196 10412 7248 10464
rect 8392 10412 8444 10464
rect 9496 10412 9548 10464
rect 11060 10412 11112 10464
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 2228 10208 2280 10260
rect 2596 10251 2648 10260
rect 2596 10217 2605 10251
rect 2605 10217 2639 10251
rect 2639 10217 2648 10251
rect 2596 10208 2648 10217
rect 3976 10208 4028 10260
rect 6000 10251 6052 10260
rect 6000 10217 6009 10251
rect 6009 10217 6043 10251
rect 6043 10217 6052 10251
rect 6000 10208 6052 10217
rect 8208 10208 8260 10260
rect 9772 10208 9824 10260
rect 12256 10208 12308 10260
rect 1584 10140 1636 10192
rect 7656 10140 7708 10192
rect 9312 10140 9364 10192
rect 9956 10140 10008 10192
rect 2964 10072 3016 10124
rect 4344 10072 4396 10124
rect 3056 10004 3108 10056
rect 4896 10004 4948 10056
rect 5172 9911 5224 9920
rect 5172 9877 5181 9911
rect 5181 9877 5215 9911
rect 5215 9877 5224 9911
rect 5172 9868 5224 9877
rect 5908 9868 5960 9920
rect 6092 9868 6144 9920
rect 6828 10072 6880 10124
rect 6644 10004 6696 10056
rect 8116 10072 8168 10124
rect 11244 10115 11296 10124
rect 11244 10081 11253 10115
rect 11253 10081 11287 10115
rect 11287 10081 11296 10115
rect 11244 10072 11296 10081
rect 7196 10004 7248 10056
rect 9588 10004 9640 10056
rect 7472 9979 7524 9988
rect 7472 9945 7481 9979
rect 7481 9945 7515 9979
rect 7515 9945 7524 9979
rect 7472 9936 7524 9945
rect 9680 9936 9732 9988
rect 12624 10004 12676 10056
rect 10140 9936 10192 9988
rect 10324 9979 10376 9988
rect 10324 9945 10333 9979
rect 10333 9945 10367 9979
rect 10367 9945 10376 9979
rect 10324 9936 10376 9945
rect 10048 9868 10100 9920
rect 10784 9868 10836 9920
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 3056 9707 3108 9716
rect 3056 9673 3065 9707
rect 3065 9673 3099 9707
rect 3099 9673 3108 9707
rect 3056 9664 3108 9673
rect 4344 9664 4396 9716
rect 4712 9664 4764 9716
rect 9956 9664 10008 9716
rect 12624 9707 12676 9716
rect 12624 9673 12633 9707
rect 12633 9673 12667 9707
rect 12667 9673 12676 9707
rect 12624 9664 12676 9673
rect 2412 9460 2464 9512
rect 2964 9460 3016 9512
rect 4068 9503 4120 9512
rect 4068 9469 4077 9503
rect 4077 9469 4111 9503
rect 4111 9469 4120 9503
rect 4068 9460 4120 9469
rect 5172 9596 5224 9648
rect 12532 9596 12584 9648
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 1860 9392 1912 9444
rect 2688 9392 2740 9444
rect 4344 9435 4396 9444
rect 4344 9401 4353 9435
rect 4353 9401 4387 9435
rect 4387 9401 4396 9435
rect 4344 9392 4396 9401
rect 5356 9460 5408 9512
rect 5908 9460 5960 9512
rect 6000 9460 6052 9512
rect 7196 9392 7248 9444
rect 8392 9392 8444 9444
rect 10048 9435 10100 9444
rect 10048 9401 10057 9435
rect 10057 9401 10091 9435
rect 10091 9401 10100 9435
rect 10048 9392 10100 9401
rect 10140 9435 10192 9444
rect 10140 9401 10149 9435
rect 10149 9401 10183 9435
rect 10183 9401 10192 9435
rect 10140 9392 10192 9401
rect 10692 9392 10744 9444
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 6644 9367 6696 9376
rect 6644 9333 6653 9367
rect 6653 9333 6687 9367
rect 6687 9333 6696 9367
rect 6644 9324 6696 9333
rect 8116 9367 8168 9376
rect 8116 9333 8125 9367
rect 8125 9333 8159 9367
rect 8159 9333 8168 9367
rect 8116 9324 8168 9333
rect 9864 9324 9916 9376
rect 11244 9367 11296 9376
rect 11244 9333 11253 9367
rect 11253 9333 11287 9367
rect 11287 9333 11296 9367
rect 11244 9324 11296 9333
rect 11520 9324 11572 9376
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 2504 9120 2556 9172
rect 2964 9120 3016 9172
rect 4068 9120 4120 9172
rect 7104 9120 7156 9172
rect 7932 9120 7984 9172
rect 9680 9120 9732 9172
rect 2688 9052 2740 9104
rect 4252 9095 4304 9104
rect 4252 9061 4261 9095
rect 4261 9061 4295 9095
rect 4295 9061 4304 9095
rect 4252 9052 4304 9061
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4436 8959 4488 8968
rect 4160 8916 4212 8925
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 2780 8891 2832 8900
rect 2780 8857 2789 8891
rect 2789 8857 2823 8891
rect 2823 8857 2832 8891
rect 2780 8848 2832 8857
rect 3240 8848 3292 8900
rect 8116 9052 8168 9104
rect 9588 9052 9640 9104
rect 9864 9095 9916 9104
rect 9864 9061 9873 9095
rect 9873 9061 9907 9095
rect 9907 9061 9916 9095
rect 9864 9052 9916 9061
rect 10968 9052 11020 9104
rect 5908 9027 5960 9036
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 6736 8984 6788 9036
rect 7472 9027 7524 9036
rect 7472 8993 7481 9027
rect 7481 8993 7515 9027
rect 7515 8993 7524 9027
rect 7472 8984 7524 8993
rect 10416 9027 10468 9036
rect 10416 8993 10425 9027
rect 10425 8993 10459 9027
rect 10459 8993 10468 9027
rect 10692 9027 10744 9036
rect 10416 8984 10468 8993
rect 10692 8993 10701 9027
rect 10701 8993 10735 9027
rect 10735 8993 10744 9027
rect 10692 8984 10744 8993
rect 12164 8984 12216 9036
rect 6000 8916 6052 8968
rect 8484 8916 8536 8968
rect 10784 8916 10836 8968
rect 12440 8916 12492 8968
rect 5724 8891 5776 8900
rect 5724 8857 5733 8891
rect 5733 8857 5767 8891
rect 5767 8857 5776 8891
rect 5724 8848 5776 8857
rect 4068 8780 4120 8832
rect 4896 8780 4948 8832
rect 5172 8780 5224 8832
rect 5356 8823 5408 8832
rect 5356 8789 5365 8823
rect 5365 8789 5399 8823
rect 5399 8789 5408 8823
rect 5356 8780 5408 8789
rect 7196 8780 7248 8832
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8392 8780 8444 8789
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 4252 8576 4304 8628
rect 5908 8576 5960 8628
rect 7288 8576 7340 8628
rect 8116 8576 8168 8628
rect 9588 8576 9640 8628
rect 10968 8619 11020 8628
rect 10968 8585 10977 8619
rect 10977 8585 11011 8619
rect 11011 8585 11020 8619
rect 10968 8576 11020 8585
rect 5080 8508 5132 8560
rect 5448 8508 5500 8560
rect 5724 8508 5776 8560
rect 7840 8508 7892 8560
rect 1952 8372 2004 8424
rect 2412 8372 2464 8424
rect 3332 8415 3384 8424
rect 3332 8381 3341 8415
rect 3341 8381 3375 8415
rect 3375 8381 3384 8415
rect 3332 8372 3384 8381
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 11244 8508 11296 8560
rect 8484 8483 8536 8492
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 10048 8440 10100 8492
rect 10416 8440 10468 8492
rect 12164 8483 12216 8492
rect 12164 8449 12173 8483
rect 12173 8449 12207 8483
rect 12207 8449 12216 8483
rect 12164 8440 12216 8449
rect 3516 8372 3568 8381
rect 2228 8304 2280 8356
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 7104 8415 7156 8424
rect 7104 8381 7113 8415
rect 7113 8381 7147 8415
rect 7147 8381 7156 8415
rect 7104 8372 7156 8381
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 12348 8372 12400 8424
rect 2688 8279 2740 8288
rect 2688 8245 2697 8279
rect 2697 8245 2731 8279
rect 2731 8245 2740 8279
rect 2688 8236 2740 8245
rect 3976 8236 4028 8288
rect 4252 8236 4304 8288
rect 5172 8236 5224 8288
rect 5448 8236 5500 8288
rect 8116 8304 8168 8356
rect 10048 8347 10100 8356
rect 7932 8236 7984 8288
rect 8392 8236 8444 8288
rect 10048 8313 10057 8347
rect 10057 8313 10091 8347
rect 10091 8313 10100 8347
rect 10048 8304 10100 8313
rect 9772 8279 9824 8288
rect 9772 8245 9781 8279
rect 9781 8245 9815 8279
rect 9815 8245 9824 8279
rect 9772 8236 9824 8245
rect 12256 8236 12308 8288
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 2688 8032 2740 8084
rect 3516 8075 3568 8084
rect 3516 8041 3525 8075
rect 3525 8041 3559 8075
rect 3559 8041 3568 8075
rect 3516 8032 3568 8041
rect 3976 8032 4028 8084
rect 4160 8032 4212 8084
rect 4896 8075 4948 8084
rect 4896 8041 4905 8075
rect 4905 8041 4939 8075
rect 4939 8041 4948 8075
rect 4896 8032 4948 8041
rect 6184 8032 6236 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 2412 7964 2464 8016
rect 5264 7964 5316 8016
rect 9772 7964 9824 8016
rect 10048 8032 10100 8084
rect 12256 8032 12308 8084
rect 2136 7896 2188 7948
rect 4068 7896 4120 7948
rect 6092 7896 6144 7948
rect 6552 7939 6604 7948
rect 6552 7905 6561 7939
rect 6561 7905 6595 7939
rect 6595 7905 6604 7939
rect 6552 7896 6604 7905
rect 7932 7896 7984 7948
rect 9496 7896 9548 7948
rect 5356 7828 5408 7880
rect 6736 7828 6788 7880
rect 10508 7896 10560 7948
rect 11244 7939 11296 7948
rect 11244 7905 11253 7939
rect 11253 7905 11287 7939
rect 11287 7905 11296 7939
rect 11244 7896 11296 7905
rect 1952 7692 2004 7744
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 6000 7692 6052 7744
rect 6184 7735 6236 7744
rect 6184 7701 6193 7735
rect 6193 7701 6227 7735
rect 6227 7701 6236 7735
rect 6184 7692 6236 7701
rect 6368 7803 6420 7812
rect 6368 7769 6377 7803
rect 6377 7769 6411 7803
rect 6411 7769 6420 7803
rect 9772 7803 9824 7812
rect 6368 7760 6420 7769
rect 9772 7769 9781 7803
rect 9781 7769 9815 7803
rect 9815 7769 9824 7803
rect 9772 7760 9824 7769
rect 7104 7692 7156 7744
rect 7196 7692 7248 7744
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 5908 7488 5960 7540
rect 6552 7488 6604 7540
rect 6736 7488 6788 7540
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 11244 7531 11296 7540
rect 11244 7497 11253 7531
rect 11253 7497 11287 7531
rect 11287 7497 11296 7531
rect 11244 7488 11296 7497
rect 6368 7463 6420 7472
rect 6368 7429 6377 7463
rect 6377 7429 6411 7463
rect 6411 7429 6420 7463
rect 6368 7420 6420 7429
rect 2228 7352 2280 7404
rect 2596 7395 2648 7404
rect 2596 7361 2605 7395
rect 2605 7361 2639 7395
rect 2639 7361 2648 7395
rect 2596 7352 2648 7361
rect 4344 7352 4396 7404
rect 6184 7352 6236 7404
rect 7380 7352 7432 7404
rect 7840 7420 7892 7472
rect 9772 7284 9824 7336
rect 2412 7191 2464 7200
rect 2412 7157 2421 7191
rect 2421 7157 2455 7191
rect 2455 7157 2464 7191
rect 2412 7148 2464 7157
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 4252 7148 4304 7200
rect 4896 7216 4948 7268
rect 6184 7216 6236 7268
rect 6644 7216 6696 7268
rect 7104 7216 7156 7268
rect 7288 7216 7340 7268
rect 8116 7216 8168 7268
rect 9312 7216 9364 7268
rect 10140 7216 10192 7268
rect 5448 7191 5500 7200
rect 5448 7157 5457 7191
rect 5457 7157 5491 7191
rect 5491 7157 5500 7191
rect 5448 7148 5500 7157
rect 10508 7148 10560 7200
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 2136 6944 2188 6996
rect 1308 6876 1360 6928
rect 1768 6876 1820 6928
rect 3240 6944 3292 6996
rect 4160 6944 4212 6996
rect 4344 6944 4396 6996
rect 7104 6944 7156 6996
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 9588 6944 9640 6996
rect 10140 6987 10192 6996
rect 10140 6953 10149 6987
rect 10149 6953 10183 6987
rect 10183 6953 10192 6987
rect 10140 6944 10192 6953
rect 10508 6987 10560 6996
rect 10508 6953 10517 6987
rect 10517 6953 10551 6987
rect 10551 6953 10560 6987
rect 10508 6944 10560 6953
rect 3516 6876 3568 6928
rect 5448 6919 5500 6928
rect 5448 6885 5457 6919
rect 5457 6885 5491 6919
rect 5491 6885 5500 6919
rect 5448 6876 5500 6885
rect 6092 6876 6144 6928
rect 2228 6808 2280 6860
rect 4068 6808 4120 6860
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 7748 6851 7800 6860
rect 7748 6817 7757 6851
rect 7757 6817 7791 6851
rect 7791 6817 7800 6851
rect 7748 6808 7800 6817
rect 8300 6808 8352 6860
rect 10140 6808 10192 6860
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 5816 6740 5868 6792
rect 3332 6672 3384 6724
rect 4436 6672 4488 6724
rect 7288 6672 7340 6724
rect 8208 6672 8260 6724
rect 2412 6604 2464 6656
rect 4252 6604 4304 6656
rect 5080 6604 5132 6656
rect 8760 6604 8812 6656
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 2504 6443 2556 6452
rect 2504 6409 2513 6443
rect 2513 6409 2547 6443
rect 2547 6409 2556 6443
rect 2504 6400 2556 6409
rect 3240 6400 3292 6452
rect 3424 6400 3476 6452
rect 4068 6400 4120 6452
rect 5448 6400 5500 6452
rect 5632 6400 5684 6452
rect 10968 6400 11020 6452
rect 13728 6400 13780 6452
rect 2780 6332 2832 6384
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 3424 6264 3476 6316
rect 4712 6332 4764 6384
rect 6920 6332 6972 6384
rect 10048 6332 10100 6384
rect 1768 6196 1820 6248
rect 2504 6196 2556 6248
rect 3148 6171 3200 6180
rect 3148 6137 3157 6171
rect 3157 6137 3191 6171
rect 3191 6137 3200 6171
rect 4712 6239 4764 6248
rect 4712 6205 4721 6239
rect 4721 6205 4755 6239
rect 4755 6205 4764 6239
rect 4712 6196 4764 6205
rect 8392 6196 8444 6248
rect 8760 6196 8812 6248
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 9496 6264 9548 6316
rect 8208 6171 8260 6180
rect 3148 6128 3200 6137
rect 8208 6137 8217 6171
rect 8217 6137 8251 6171
rect 8251 6137 8260 6171
rect 8208 6128 8260 6137
rect 8852 6171 8904 6180
rect 8852 6137 8861 6171
rect 8861 6137 8895 6171
rect 8895 6137 8904 6171
rect 8852 6128 8904 6137
rect 9956 6128 10008 6180
rect 3240 6060 3292 6112
rect 4528 6060 4580 6112
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 6644 6103 6696 6112
rect 6644 6069 6653 6103
rect 6653 6069 6687 6103
rect 6687 6069 6696 6103
rect 6644 6060 6696 6069
rect 7748 6060 7800 6112
rect 7932 6060 7984 6112
rect 8944 6060 8996 6112
rect 10140 6103 10192 6112
rect 10140 6069 10149 6103
rect 10149 6069 10183 6103
rect 10183 6069 10192 6103
rect 10140 6060 10192 6069
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 1860 5856 1912 5908
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 3516 5856 3568 5908
rect 6092 5856 6144 5908
rect 7564 5856 7616 5908
rect 10140 5899 10192 5908
rect 10140 5865 10149 5899
rect 10149 5865 10183 5899
rect 10183 5865 10192 5899
rect 10140 5856 10192 5865
rect 2228 5788 2280 5840
rect 2504 5763 2556 5772
rect 2504 5729 2513 5763
rect 2513 5729 2547 5763
rect 2547 5729 2556 5763
rect 2504 5720 2556 5729
rect 2780 5652 2832 5704
rect 8944 5788 8996 5840
rect 3976 5720 4028 5772
rect 4252 5720 4304 5772
rect 6092 5763 6144 5772
rect 4436 5652 4488 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 2872 5584 2924 5636
rect 4988 5584 5040 5636
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 3424 5516 3476 5525
rect 6092 5729 6101 5763
rect 6101 5729 6135 5763
rect 6135 5729 6144 5763
rect 6092 5720 6144 5729
rect 6276 5720 6328 5772
rect 7196 5720 7248 5772
rect 8668 5720 8720 5772
rect 9404 5720 9456 5772
rect 9956 5763 10008 5772
rect 9956 5729 9965 5763
rect 9965 5729 9999 5763
rect 9999 5729 10008 5763
rect 9956 5720 10008 5729
rect 7932 5652 7984 5704
rect 7748 5584 7800 5636
rect 8208 5584 8260 5636
rect 8484 5584 8536 5636
rect 9128 5627 9180 5636
rect 9128 5593 9137 5627
rect 9137 5593 9171 5627
rect 9171 5593 9180 5627
rect 9128 5584 9180 5593
rect 10140 5584 10192 5636
rect 5356 5516 5408 5568
rect 7104 5516 7156 5568
rect 7269 5559 7321 5568
rect 7269 5525 7278 5559
rect 7278 5525 7312 5559
rect 7312 5525 7321 5559
rect 7269 5516 7321 5525
rect 9312 5516 9364 5568
rect 10232 5516 10284 5568
rect 10324 5516 10376 5568
rect 12072 5516 12124 5568
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 1860 5312 1912 5364
rect 3976 5312 4028 5364
rect 4252 5355 4304 5364
rect 4252 5321 4261 5355
rect 4261 5321 4295 5355
rect 4295 5321 4304 5355
rect 4252 5312 4304 5321
rect 6276 5355 6328 5364
rect 6276 5321 6285 5355
rect 6285 5321 6319 5355
rect 6319 5321 6328 5355
rect 6276 5312 6328 5321
rect 9312 5312 9364 5364
rect 9772 5355 9824 5364
rect 9772 5321 9781 5355
rect 9781 5321 9815 5355
rect 9815 5321 9824 5355
rect 9772 5312 9824 5321
rect 9956 5312 10008 5364
rect 2780 5287 2832 5296
rect 2780 5253 2789 5287
rect 2789 5253 2823 5287
rect 2823 5253 2832 5287
rect 2780 5244 2832 5253
rect 6644 5287 6696 5296
rect 3332 5176 3384 5228
rect 1860 5151 1912 5160
rect 1860 5117 1869 5151
rect 1869 5117 1903 5151
rect 1903 5117 1912 5151
rect 1860 5108 1912 5117
rect 2504 5108 2556 5160
rect 2412 5083 2464 5092
rect 2412 5049 2421 5083
rect 2421 5049 2455 5083
rect 2455 5049 2464 5083
rect 2412 5040 2464 5049
rect 3332 5083 3384 5092
rect 3332 5049 3341 5083
rect 3341 5049 3375 5083
rect 3375 5049 3384 5083
rect 3332 5040 3384 5049
rect 6644 5253 6653 5287
rect 6653 5253 6687 5287
rect 6687 5253 6696 5287
rect 6644 5244 6696 5253
rect 8484 5287 8536 5296
rect 8484 5253 8493 5287
rect 8493 5253 8527 5287
rect 8527 5253 8536 5287
rect 8484 5244 8536 5253
rect 10140 5244 10192 5296
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 6644 5108 6696 5160
rect 7288 5176 7340 5228
rect 9404 5176 9456 5228
rect 7104 5151 7156 5160
rect 7104 5117 7113 5151
rect 7113 5117 7147 5151
rect 7147 5117 7156 5151
rect 7104 5108 7156 5117
rect 7472 5108 7524 5160
rect 8392 5151 8444 5160
rect 8392 5117 8401 5151
rect 8401 5117 8435 5151
rect 8435 5117 8444 5151
rect 8392 5108 8444 5117
rect 8668 5151 8720 5160
rect 8668 5117 8677 5151
rect 8677 5117 8711 5151
rect 8711 5117 8720 5151
rect 8668 5108 8720 5117
rect 8760 5108 8812 5160
rect 9956 5151 10008 5160
rect 9956 5117 9965 5151
rect 9965 5117 9999 5151
rect 9999 5117 10008 5151
rect 9956 5108 10008 5117
rect 10232 5151 10284 5160
rect 10232 5117 10241 5151
rect 10241 5117 10275 5151
rect 10275 5117 10284 5151
rect 10232 5108 10284 5117
rect 2964 4972 3016 5024
rect 7656 5040 7708 5092
rect 11060 5040 11112 5092
rect 4344 4972 4396 5024
rect 4620 4972 4672 5024
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 6000 4972 6052 5024
rect 7932 5015 7984 5024
rect 7932 4981 7941 5015
rect 7941 4981 7975 5015
rect 7975 4981 7984 5015
rect 7932 4972 7984 4981
rect 8484 4972 8536 5024
rect 9312 4972 9364 5024
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 2504 4768 2556 4820
rect 4712 4811 4764 4820
rect 4712 4777 4721 4811
rect 4721 4777 4755 4811
rect 4755 4777 4764 4811
rect 4712 4768 4764 4777
rect 2596 4743 2648 4752
rect 2596 4709 2605 4743
rect 2605 4709 2639 4743
rect 2639 4709 2648 4743
rect 2596 4700 2648 4709
rect 3148 4700 3200 4752
rect 5724 4768 5776 4820
rect 6092 4811 6144 4820
rect 6092 4777 6101 4811
rect 6101 4777 6135 4811
rect 6135 4777 6144 4811
rect 6092 4768 6144 4777
rect 7748 4811 7800 4820
rect 5080 4700 5132 4752
rect 1676 4632 1728 4684
rect 5724 4632 5776 4684
rect 6828 4743 6880 4752
rect 6828 4709 6837 4743
rect 6837 4709 6871 4743
rect 6871 4709 6880 4743
rect 6828 4700 6880 4709
rect 7380 4743 7432 4752
rect 7380 4709 7389 4743
rect 7389 4709 7423 4743
rect 7423 4709 7432 4743
rect 7380 4700 7432 4709
rect 7748 4777 7757 4811
rect 7757 4777 7791 4811
rect 7791 4777 7800 4811
rect 7748 4768 7800 4777
rect 8024 4700 8076 4752
rect 8392 4700 8444 4752
rect 9404 4743 9456 4752
rect 9404 4709 9413 4743
rect 9413 4709 9447 4743
rect 9447 4709 9456 4743
rect 9404 4700 9456 4709
rect 10048 4632 10100 4684
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 11244 4675 11296 4684
rect 11244 4641 11253 4675
rect 11253 4641 11287 4675
rect 11287 4641 11296 4675
rect 11244 4632 11296 4641
rect 2044 4564 2096 4616
rect 3240 4564 3292 4616
rect 5356 4564 5408 4616
rect 8116 4564 8168 4616
rect 4804 4496 4856 4548
rect 7564 4496 7616 4548
rect 1768 4428 1820 4480
rect 3332 4428 3384 4480
rect 3976 4428 4028 4480
rect 5816 4471 5868 4480
rect 5816 4437 5825 4471
rect 5825 4437 5859 4471
rect 5859 4437 5868 4471
rect 5816 4428 5868 4437
rect 6644 4428 6696 4480
rect 8392 4471 8444 4480
rect 8392 4437 8401 4471
rect 8401 4437 8435 4471
rect 8435 4437 8444 4471
rect 8392 4428 8444 4437
rect 9956 4428 10008 4480
rect 10784 4428 10836 4480
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 5816 4224 5868 4276
rect 6828 4224 6880 4276
rect 8024 4224 8076 4276
rect 8668 4267 8720 4276
rect 8668 4233 8677 4267
rect 8677 4233 8711 4267
rect 8711 4233 8720 4267
rect 8668 4224 8720 4233
rect 10048 4224 10100 4276
rect 11336 4224 11388 4276
rect 7564 4156 7616 4208
rect 7932 4156 7984 4208
rect 8852 4156 8904 4208
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 4620 4088 4672 4140
rect 7012 4088 7064 4140
rect 7104 4088 7156 4140
rect 8760 4063 8812 4072
rect 8760 4029 8769 4063
rect 8769 4029 8803 4063
rect 8803 4029 8812 4063
rect 8760 4020 8812 4029
rect 12164 4156 12216 4208
rect 10416 4020 10468 4072
rect 11152 4020 11204 4072
rect 11244 4020 11296 4072
rect 11428 4020 11480 4072
rect 2688 3952 2740 4004
rect 2596 3927 2648 3936
rect 2596 3893 2605 3927
rect 2605 3893 2639 3927
rect 2639 3893 2648 3927
rect 2596 3884 2648 3893
rect 2780 3884 2832 3936
rect 2964 3995 3016 4004
rect 2964 3961 2973 3995
rect 2973 3961 3007 3995
rect 3007 3961 3016 3995
rect 2964 3952 3016 3961
rect 5080 3884 5132 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 6828 3884 6880 3936
rect 8116 3952 8168 4004
rect 10692 3952 10744 4004
rect 12072 3952 12124 4004
rect 11980 3884 12032 3936
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 2504 3723 2556 3732
rect 2504 3689 2513 3723
rect 2513 3689 2547 3723
rect 2547 3689 2556 3723
rect 2504 3680 2556 3689
rect 4436 3680 4488 3732
rect 4896 3680 4948 3732
rect 5724 3723 5776 3732
rect 5724 3689 5733 3723
rect 5733 3689 5767 3723
rect 5767 3689 5776 3723
rect 5724 3680 5776 3689
rect 7564 3723 7616 3732
rect 7564 3689 7573 3723
rect 7573 3689 7607 3723
rect 7607 3689 7616 3723
rect 7564 3680 7616 3689
rect 9864 3723 9916 3732
rect 2044 3655 2096 3664
rect 2044 3621 2053 3655
rect 2053 3621 2087 3655
rect 2087 3621 2096 3655
rect 2044 3612 2096 3621
rect 5080 3612 5132 3664
rect 5356 3612 5408 3664
rect 6276 3612 6328 3664
rect 1768 3544 1820 3596
rect 5264 3544 5316 3596
rect 2412 3476 2464 3528
rect 3516 3476 3568 3528
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 7932 3655 7984 3664
rect 7932 3621 7941 3655
rect 7941 3621 7975 3655
rect 7975 3621 7984 3655
rect 7932 3612 7984 3621
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 15752 3680 15804 3732
rect 11980 3612 12032 3664
rect 2780 3408 2832 3460
rect 5908 3408 5960 3460
rect 7104 3408 7156 3460
rect 7748 3408 7800 3460
rect 8300 3476 8352 3528
rect 10324 3544 10376 3596
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 12072 3544 12124 3596
rect 12164 3544 12216 3596
rect 13268 3587 13320 3596
rect 13268 3553 13277 3587
rect 13277 3553 13311 3587
rect 13311 3553 13320 3587
rect 13268 3544 13320 3553
rect 2596 3340 2648 3392
rect 3424 3383 3476 3392
rect 3424 3349 3433 3383
rect 3433 3349 3467 3383
rect 3467 3349 3476 3383
rect 3424 3340 3476 3349
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 6644 3340 6696 3392
rect 7012 3340 7064 3392
rect 7380 3340 7432 3392
rect 15200 3408 15252 3460
rect 9312 3340 9364 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 2964 3136 3016 3188
rect 3516 3179 3568 3188
rect 3516 3145 3525 3179
rect 3525 3145 3559 3179
rect 3559 3145 3568 3179
rect 3516 3136 3568 3145
rect 1676 3068 1728 3120
rect 4896 3136 4948 3188
rect 6276 3179 6328 3188
rect 6276 3145 6285 3179
rect 6285 3145 6319 3179
rect 6319 3145 6328 3179
rect 6276 3136 6328 3145
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 5264 3043 5316 3052
rect 5264 3009 5273 3043
rect 5273 3009 5307 3043
rect 5307 3009 5316 3043
rect 5264 3000 5316 3009
rect 5908 3043 5960 3052
rect 5908 3009 5917 3043
rect 5917 3009 5951 3043
rect 5951 3009 5960 3043
rect 5908 3000 5960 3009
rect 2504 2864 2556 2916
rect 2780 2864 2832 2916
rect 4344 2864 4396 2916
rect 5356 2907 5408 2916
rect 5356 2873 5365 2907
rect 5365 2873 5399 2907
rect 5399 2873 5408 2907
rect 5356 2864 5408 2873
rect 6644 3136 6696 3188
rect 7932 3179 7984 3188
rect 7932 3145 7941 3179
rect 7941 3145 7975 3179
rect 7975 3145 7984 3179
rect 7932 3136 7984 3145
rect 10324 3136 10376 3188
rect 10600 3179 10652 3188
rect 10600 3145 10609 3179
rect 10609 3145 10643 3179
rect 10643 3145 10652 3179
rect 10600 3136 10652 3145
rect 11152 3136 11204 3188
rect 12164 3179 12216 3188
rect 12164 3145 12173 3179
rect 12173 3145 12207 3179
rect 12207 3145 12216 3179
rect 12164 3136 12216 3145
rect 12256 3136 12308 3188
rect 7380 3068 7432 3120
rect 7656 3068 7708 3120
rect 7564 3000 7616 3052
rect 10692 3068 10744 3120
rect 12440 3068 12492 3120
rect 10876 3000 10928 3052
rect 10600 2932 10652 2984
rect 11152 2975 11204 2984
rect 11152 2941 11161 2975
rect 11161 2941 11195 2975
rect 11195 2941 11204 2975
rect 11152 2932 11204 2941
rect 11520 2932 11572 2984
rect 13820 2932 13872 2984
rect 8300 2864 8352 2916
rect 3240 2796 3292 2848
rect 4252 2839 4304 2848
rect 4252 2805 4261 2839
rect 4261 2805 4295 2839
rect 4295 2805 4304 2839
rect 4252 2796 4304 2805
rect 5080 2839 5132 2848
rect 5080 2805 5089 2839
rect 5089 2805 5123 2839
rect 5123 2805 5132 2839
rect 5080 2796 5132 2805
rect 5540 2796 5592 2848
rect 6644 2796 6696 2848
rect 7104 2796 7156 2848
rect 11980 2796 12032 2848
rect 13268 2839 13320 2848
rect 13268 2805 13277 2839
rect 13277 2805 13311 2839
rect 13311 2805 13320 2839
rect 13268 2796 13320 2805
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 2780 2592 2832 2644
rect 2596 2567 2648 2576
rect 2596 2533 2605 2567
rect 2605 2533 2639 2567
rect 2639 2533 2648 2567
rect 2596 2524 2648 2533
rect 3332 2592 3384 2644
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 3240 2524 3292 2576
rect 5080 2524 5132 2576
rect 5356 2567 5408 2576
rect 5356 2533 5365 2567
rect 5365 2533 5399 2567
rect 5399 2533 5408 2567
rect 5356 2524 5408 2533
rect 7012 2524 7064 2576
rect 7104 2567 7156 2576
rect 7104 2533 7113 2567
rect 7113 2533 7147 2567
rect 7147 2533 7156 2567
rect 7104 2524 7156 2533
rect 4528 2456 4580 2508
rect 5540 2456 5592 2508
rect 8576 2456 8628 2508
rect 9864 2499 9916 2508
rect 9864 2465 9873 2499
rect 9873 2465 9907 2499
rect 9907 2465 9916 2499
rect 9864 2456 9916 2465
rect 10968 2456 11020 2508
rect 12532 2456 12584 2508
rect 13268 2456 13320 2508
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 6000 2320 6052 2372
rect 9864 2320 9916 2372
rect 13360 2320 13412 2372
rect 1768 2252 1820 2304
rect 7104 2252 7156 2304
rect 8300 2295 8352 2304
rect 8300 2261 8309 2295
rect 8309 2261 8343 2295
rect 8343 2261 8352 2295
rect 8300 2252 8352 2261
rect 8668 2295 8720 2304
rect 8668 2261 8677 2295
rect 8677 2261 8711 2295
rect 8711 2261 8720 2295
rect 8668 2252 8720 2261
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 1768 2048 1820 2100
rect 7748 2048 7800 2100
rect 8300 2048 8352 2100
rect 1492 1980 1544 2032
rect 5540 1980 5592 2032
rect 5080 1912 5132 1964
rect 10232 1912 10284 1964
rect 4068 1776 4120 1828
rect 5264 1708 5316 1760
rect 8668 1164 8720 1216
rect 13728 1164 13780 1216
rect 296 76 348 128
rect 1032 76 1084 128
rect 1492 76 1544 128
rect 2044 76 2096 128
rect 4252 76 4304 128
rect 12072 76 12124 128
rect 848 8 900 60
rect 5172 8 5224 60
<< metal2 >>
rect 386 39704 442 40000
rect 386 39652 388 39704
rect 440 39652 442 39704
rect 386 39520 442 39652
rect 1214 39658 1270 40000
rect 1214 39630 1348 39658
rect 1214 39520 1270 39630
rect 1030 31920 1086 31929
rect 1030 31855 1086 31864
rect 1044 30394 1072 31855
rect 1032 30388 1084 30394
rect 1032 30330 1084 30336
rect 1122 26888 1178 26897
rect 1122 26823 1178 26832
rect 1136 23322 1164 26823
rect 1320 25838 1348 39630
rect 1492 39636 1544 39642
rect 1492 39578 1544 39584
rect 2134 39636 2190 40000
rect 2134 39584 2136 39636
rect 2188 39584 2190 39636
rect 1504 28626 1532 39578
rect 2134 39520 2190 39584
rect 3054 39636 3110 40000
rect 3054 39584 3056 39636
rect 3108 39584 3110 39636
rect 3054 39520 3110 39584
rect 3882 39636 3938 40000
rect 4802 39658 4858 40000
rect 3882 39584 3884 39636
rect 3936 39584 3938 39636
rect 3882 39520 3938 39584
rect 4356 39630 4858 39658
rect 5540 39704 5592 39710
rect 5540 39646 5592 39652
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3148 30048 3200 30054
rect 3148 29990 3200 29996
rect 1492 28620 1544 28626
rect 1492 28562 1544 28568
rect 1308 25832 1360 25838
rect 1308 25774 1360 25780
rect 1124 23316 1176 23322
rect 1124 23258 1176 23264
rect 1306 22264 1362 22273
rect 1306 22199 1362 22208
rect 1320 22166 1348 22199
rect 1308 22160 1360 22166
rect 1308 22102 1360 22108
rect 1306 16960 1362 16969
rect 1306 16895 1362 16904
rect 1320 16114 1348 16895
rect 1308 16108 1360 16114
rect 1308 16050 1360 16056
rect 1504 13814 1532 28562
rect 2964 27396 3016 27402
rect 2964 27338 3016 27344
rect 2412 26784 2464 26790
rect 2412 26726 2464 26732
rect 2424 26586 2452 26726
rect 2412 26580 2464 26586
rect 2412 26522 2464 26528
rect 2320 25832 2372 25838
rect 2320 25774 2372 25780
rect 2228 25288 2280 25294
rect 2228 25230 2280 25236
rect 1952 24744 2004 24750
rect 1952 24686 2004 24692
rect 1964 23866 1992 24686
rect 2240 24410 2268 25230
rect 2332 24857 2360 25774
rect 2596 25696 2648 25702
rect 2596 25638 2648 25644
rect 2608 25498 2636 25638
rect 2596 25492 2648 25498
rect 2596 25434 2648 25440
rect 2318 24848 2374 24857
rect 2318 24783 2374 24792
rect 2608 24614 2636 25434
rect 2976 24818 3004 27338
rect 3160 27010 3188 29990
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3974 28520 4030 28529
rect 3974 28455 4030 28464
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3988 28150 4016 28455
rect 3976 28144 4028 28150
rect 3976 28086 4028 28092
rect 3332 27940 3384 27946
rect 3332 27882 3384 27888
rect 3240 27532 3292 27538
rect 3240 27474 3292 27480
rect 3252 27130 3280 27474
rect 3240 27124 3292 27130
rect 3240 27066 3292 27072
rect 3160 26982 3280 27010
rect 3148 26512 3200 26518
rect 3148 26454 3200 26460
rect 3160 25974 3188 26454
rect 3148 25968 3200 25974
rect 3148 25910 3200 25916
rect 3160 25226 3188 25910
rect 3148 25220 3200 25226
rect 3148 25162 3200 25168
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2596 24608 2648 24614
rect 2596 24550 2648 24556
rect 2228 24404 2280 24410
rect 2228 24346 2280 24352
rect 2688 24268 2740 24274
rect 2688 24210 2740 24216
rect 1952 23860 2004 23866
rect 1952 23802 2004 23808
rect 1964 23662 1992 23802
rect 2700 23662 2728 24210
rect 3148 24200 3200 24206
rect 3148 24142 3200 24148
rect 1952 23656 2004 23662
rect 1952 23598 2004 23604
rect 2136 23656 2188 23662
rect 2136 23598 2188 23604
rect 2688 23656 2740 23662
rect 2688 23598 2740 23604
rect 1584 23588 1636 23594
rect 1584 23530 1636 23536
rect 1596 20058 1624 23530
rect 2044 23180 2096 23186
rect 2044 23122 2096 23128
rect 1768 22976 1820 22982
rect 1768 22918 1820 22924
rect 1676 22432 1728 22438
rect 1676 22374 1728 22380
rect 1688 22030 1716 22374
rect 1676 22024 1728 22030
rect 1676 21966 1728 21972
rect 1780 21894 1808 22918
rect 2056 22778 2084 23122
rect 2148 23050 2176 23598
rect 2700 23474 2728 23598
rect 3160 23526 3188 24142
rect 2608 23446 2728 23474
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 2608 23118 2636 23446
rect 3056 23180 3108 23186
rect 3056 23122 3108 23128
rect 2596 23112 2648 23118
rect 2596 23054 2648 23060
rect 2136 23044 2188 23050
rect 2136 22986 2188 22992
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2688 22976 2740 22982
rect 2688 22918 2740 22924
rect 2044 22772 2096 22778
rect 2044 22714 2096 22720
rect 2228 22432 2280 22438
rect 2228 22374 2280 22380
rect 2240 22166 2268 22374
rect 2228 22160 2280 22166
rect 2228 22102 2280 22108
rect 2596 22160 2648 22166
rect 2596 22102 2648 22108
rect 1768 21888 1820 21894
rect 1768 21830 1820 21836
rect 1780 21486 1808 21830
rect 2240 21690 2268 22102
rect 2228 21684 2280 21690
rect 2228 21626 2280 21632
rect 1676 21480 1728 21486
rect 1676 21422 1728 21428
rect 1768 21480 1820 21486
rect 1768 21422 1820 21428
rect 1688 21146 1716 21422
rect 1676 21140 1728 21146
rect 1676 21082 1728 21088
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1596 19446 1624 19994
rect 1584 19440 1636 19446
rect 1584 19382 1636 19388
rect 1688 18970 1716 21082
rect 1780 20466 1808 21422
rect 2608 21146 2636 22102
rect 2596 21140 2648 21146
rect 2596 21082 2648 21088
rect 2596 20936 2648 20942
rect 2596 20878 2648 20884
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 1780 19514 1808 20402
rect 1860 20392 1912 20398
rect 1860 20334 1912 20340
rect 1872 19718 1900 20334
rect 2608 20330 2636 20878
rect 2596 20324 2648 20330
rect 2596 20266 2648 20272
rect 2608 20058 2636 20266
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2412 19780 2464 19786
rect 2412 19722 2464 19728
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1768 19508 1820 19514
rect 1768 19450 1820 19456
rect 1676 18964 1728 18970
rect 1596 18924 1676 18952
rect 1596 15094 1624 18924
rect 1676 18906 1728 18912
rect 1768 18352 1820 18358
rect 1768 18294 1820 18300
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 16658 1716 16934
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1688 15706 1716 16594
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1584 15088 1636 15094
rect 1584 15030 1636 15036
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1596 14414 1624 14894
rect 1780 14482 1808 18294
rect 1872 16998 1900 19654
rect 2228 18896 2280 18902
rect 1950 18864 2006 18873
rect 2228 18838 2280 18844
rect 1950 18799 2006 18808
rect 1964 18766 1992 18799
rect 1952 18760 2004 18766
rect 1952 18702 2004 18708
rect 1964 18222 1992 18702
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 1952 18080 2004 18086
rect 2056 18068 2084 18566
rect 2240 18086 2268 18838
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2004 18040 2084 18068
rect 2228 18080 2280 18086
rect 1952 18022 2004 18028
rect 2228 18022 2280 18028
rect 1964 17542 1992 18022
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17134 1992 17478
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1504 13786 1716 13814
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1030 11792 1086 11801
rect 1412 11762 1440 13262
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1030 11727 1086 11736
rect 1400 11756 1452 11762
rect 294 128 350 480
rect 294 76 296 128
rect 348 76 350 128
rect 294 0 350 76
rect 846 60 902 480
rect 1044 134 1072 11727
rect 1400 11698 1452 11704
rect 1306 7032 1362 7041
rect 1306 6967 1362 6976
rect 1320 6934 1348 6967
rect 1308 6928 1360 6934
rect 1308 6870 1360 6876
rect 1504 2038 1532 12242
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1596 10606 1624 11834
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1596 10198 1624 10542
rect 1584 10192 1636 10198
rect 1582 10160 1584 10169
rect 1636 10160 1638 10169
rect 1582 10095 1638 10104
rect 1688 4690 1716 13786
rect 1780 13190 1808 14418
rect 1872 13814 1900 16934
rect 1964 15162 1992 17070
rect 2056 16250 2084 17614
rect 2136 17060 2188 17066
rect 2136 17002 2188 17008
rect 2148 16726 2176 17002
rect 2136 16720 2188 16726
rect 2136 16662 2188 16668
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2056 15638 2084 16186
rect 2148 15978 2176 16662
rect 2136 15972 2188 15978
rect 2136 15914 2188 15920
rect 2044 15632 2096 15638
rect 2044 15574 2096 15580
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 2240 13938 2268 18022
rect 2332 17678 2360 18770
rect 2424 18426 2452 19722
rect 2596 19304 2648 19310
rect 2700 19292 2728 22918
rect 2792 22778 2820 22986
rect 3068 22778 3096 23122
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 3056 22772 3108 22778
rect 3056 22714 3108 22720
rect 3056 21888 3108 21894
rect 3160 21876 3188 23462
rect 3108 21848 3188 21876
rect 3056 21830 3108 21836
rect 2872 21412 2924 21418
rect 2872 21354 2924 21360
rect 2884 21078 2912 21354
rect 2872 21072 2924 21078
rect 2872 21014 2924 21020
rect 2884 20602 2912 21014
rect 2872 20596 2924 20602
rect 2872 20538 2924 20544
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 2976 19961 3004 20334
rect 2962 19952 3018 19961
rect 2962 19887 3018 19896
rect 2976 19854 3004 19887
rect 2964 19848 3016 19854
rect 2964 19790 3016 19796
rect 2648 19264 2728 19292
rect 2780 19304 2832 19310
rect 2596 19246 2648 19252
rect 2780 19246 2832 19252
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2320 17536 2372 17542
rect 2320 17478 2372 17484
rect 2332 16046 2360 17478
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2332 15434 2360 15982
rect 2424 15570 2452 18362
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2320 15428 2372 15434
rect 2320 15370 2372 15376
rect 2424 15094 2452 15506
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2424 14634 2452 15030
rect 2424 14606 2544 14634
rect 2412 14476 2464 14482
rect 2412 14418 2464 14424
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2332 13870 2360 14214
rect 2424 14006 2452 14418
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 2516 13938 2544 14606
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2320 13864 2372 13870
rect 1872 13786 2084 13814
rect 2320 13806 2372 13812
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2502 13832 2558 13841
rect 1860 13728 1912 13734
rect 1860 13670 1912 13676
rect 1872 13530 1900 13670
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1780 12306 1808 13126
rect 1768 12300 1820 12306
rect 1768 12242 1820 12248
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1768 12164 1820 12170
rect 1768 12106 1820 12112
rect 1780 11354 1808 12106
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1872 11150 1900 12174
rect 2056 11898 2084 13786
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2332 12782 2360 13126
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 2240 12306 2268 12650
rect 2424 12646 2452 13806
rect 2608 13814 2636 19246
rect 2792 18834 2820 19246
rect 3068 18902 3096 21830
rect 3148 21480 3200 21486
rect 3148 21422 3200 21428
rect 3160 21146 3188 21422
rect 3148 21140 3200 21146
rect 3148 21082 3200 21088
rect 3252 19854 3280 26982
rect 3344 26790 3372 27882
rect 4356 27538 4384 39630
rect 4802 39520 4858 39630
rect 5080 39636 5132 39642
rect 5080 39578 5132 39584
rect 4620 34604 4672 34610
rect 4620 34546 4672 34552
rect 4436 28552 4488 28558
rect 4436 28494 4488 28500
rect 4448 28218 4476 28494
rect 4632 28218 4660 34546
rect 5092 28966 5120 39578
rect 5264 34400 5316 34406
rect 5264 34342 5316 34348
rect 5080 28960 5132 28966
rect 5080 28902 5132 28908
rect 4988 28620 5040 28626
rect 4988 28562 5040 28568
rect 5000 28218 5028 28562
rect 4436 28212 4488 28218
rect 4436 28154 4488 28160
rect 4620 28212 4672 28218
rect 4620 28154 4672 28160
rect 4988 28212 5040 28218
rect 4988 28154 5040 28160
rect 4632 27946 4660 28154
rect 4620 27940 4672 27946
rect 4620 27882 4672 27888
rect 4988 27940 5040 27946
rect 4988 27882 5040 27888
rect 5000 27674 5028 27882
rect 4988 27668 5040 27674
rect 4988 27610 5040 27616
rect 4344 27532 4396 27538
rect 4344 27474 4396 27480
rect 3516 27328 3568 27334
rect 3516 27270 3568 27276
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 3528 26994 3556 27270
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 3332 26784 3384 26790
rect 3332 26726 3384 26732
rect 3344 23474 3372 26726
rect 3528 26586 3556 26930
rect 3608 26852 3660 26858
rect 3608 26794 3660 26800
rect 3516 26580 3568 26586
rect 3516 26522 3568 26528
rect 3516 26240 3568 26246
rect 3620 26228 3648 26794
rect 3568 26200 3648 26228
rect 3516 26182 3568 26188
rect 3528 25838 3556 26182
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3424 25832 3476 25838
rect 3424 25774 3476 25780
rect 3516 25832 3568 25838
rect 3516 25774 3568 25780
rect 3436 25158 3464 25774
rect 4080 25276 4108 27270
rect 4356 27130 4384 27474
rect 5000 27470 5028 27610
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 4344 27124 4396 27130
rect 4344 27066 4396 27072
rect 4160 26444 4212 26450
rect 4160 26386 4212 26392
rect 4172 26042 4200 26386
rect 4160 26036 4212 26042
rect 4160 25978 4212 25984
rect 4252 25832 4304 25838
rect 4252 25774 4304 25780
rect 4264 25430 4292 25774
rect 4252 25424 4304 25430
rect 4252 25366 4304 25372
rect 4160 25288 4212 25294
rect 4080 25248 4160 25276
rect 4160 25230 4212 25236
rect 3424 25152 3476 25158
rect 3424 25094 3476 25100
rect 3516 25152 3568 25158
rect 3516 25094 3568 25100
rect 3436 23730 3464 25094
rect 3528 24954 3556 25094
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3516 24948 3568 24954
rect 3516 24890 3568 24896
rect 4252 24880 4304 24886
rect 4252 24822 4304 24828
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3896 24052 3924 24686
rect 3976 24608 4028 24614
rect 4160 24608 4212 24614
rect 4028 24568 4160 24596
rect 3976 24550 4028 24556
rect 3976 24064 4028 24070
rect 3896 24024 3976 24052
rect 3976 24006 4028 24012
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3344 23446 3556 23474
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 3424 19236 3476 19242
rect 3424 19178 3476 19184
rect 3056 18896 3108 18902
rect 3056 18838 3108 18844
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2976 18290 3004 18702
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2688 17808 2740 17814
rect 2688 17750 2740 17756
rect 2700 16794 2728 17750
rect 2792 17066 2820 18022
rect 2976 17882 3004 18226
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 3436 17746 3464 19178
rect 3424 17740 3476 17746
rect 3424 17682 3476 17688
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 3160 16454 3188 17070
rect 3436 16794 3464 17682
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3068 16046 3096 16390
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2976 15162 3004 15506
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2976 14958 3004 15098
rect 3068 15026 3096 15982
rect 3160 15638 3188 16390
rect 3240 16176 3292 16182
rect 3240 16118 3292 16124
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2700 14074 2728 14418
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2792 13841 2820 14894
rect 3252 14482 3280 16118
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3056 13864 3108 13870
rect 2778 13832 2834 13841
rect 2608 13786 2728 13814
rect 2502 13767 2558 13776
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 2136 11620 2188 11626
rect 2332 11608 2360 12038
rect 2188 11580 2360 11608
rect 2136 11562 2188 11568
rect 2332 11354 2360 11580
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2516 11218 2544 13767
rect 2700 13394 2728 13786
rect 3056 13806 3108 13812
rect 2778 13767 2834 13776
rect 2872 13796 2924 13802
rect 2872 13738 2924 13744
rect 2884 13394 2912 13738
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2700 12442 2728 13330
rect 2884 12782 2912 13330
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 1872 10470 1900 11086
rect 1964 10538 1992 11154
rect 2516 10810 2544 11154
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 1952 10532 2004 10538
rect 1952 10474 2004 10480
rect 1860 10464 1912 10470
rect 1860 10406 1912 10412
rect 1964 9489 1992 10474
rect 2240 10266 2268 10542
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2412 9512 2464 9518
rect 1950 9480 2006 9489
rect 1860 9444 1912 9450
rect 2516 9500 2544 10746
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2464 9472 2544 9500
rect 2412 9454 2464 9460
rect 1950 9415 2006 9424
rect 1860 9386 1912 9392
rect 1768 6928 1820 6934
rect 1768 6870 1820 6876
rect 1780 6254 1808 6870
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1872 5914 1900 9386
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 7750 1992 8366
rect 2148 7954 2176 9318
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2240 8362 2268 8910
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1964 6322 1992 7686
rect 2148 7002 2176 7890
rect 2240 7410 2268 8298
rect 2424 8022 2452 8366
rect 2412 8016 2464 8022
rect 2412 7958 2464 7964
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2424 7206 2452 7958
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1872 5370 1900 5850
rect 2240 5846 2268 6802
rect 2424 6662 2452 7142
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2516 6458 2544 9114
rect 2608 7410 2636 10202
rect 2700 9450 2728 12378
rect 2792 10452 2820 12582
rect 2884 12238 2912 12718
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2884 11218 2912 12174
rect 2976 11762 3004 13670
rect 3068 13462 3096 13806
rect 3160 13734 3188 14282
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3436 13870 3464 14214
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2976 11354 3004 11698
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2884 10606 2912 11154
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2792 10424 2912 10452
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2700 8294 2728 9046
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2700 8090 2728 8230
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2792 6798 2820 8842
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2516 6254 2544 6394
rect 2792 6390 2820 6734
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2504 6248 2556 6254
rect 2884 6236 2912 10424
rect 2976 10130 3004 11018
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2976 9518 3004 10066
rect 3068 10062 3096 13398
rect 3240 13252 3292 13258
rect 3160 13212 3240 13240
rect 3160 12782 3188 13212
rect 3240 13194 3292 13200
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3160 11286 3188 12718
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 3344 11898 3372 12310
rect 3332 11892 3384 11898
rect 3332 11834 3384 11840
rect 3344 11558 3372 11834
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3344 11014 3372 11494
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3238 10160 3294 10169
rect 3238 10095 3294 10104
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3068 9722 3096 9998
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 2976 9178 3004 9454
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3252 8906 3280 10095
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 2504 6190 2556 6196
rect 2792 6208 2912 6236
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2228 5840 2280 5846
rect 2228 5782 2280 5788
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1872 5166 1900 5306
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1688 4146 1716 4626
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1688 3126 1716 4082
rect 1780 3602 1808 4422
rect 2056 3670 2084 4558
rect 2044 3664 2096 3670
rect 2044 3606 2096 3612
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 2056 3505 2084 3606
rect 2042 3496 2098 3505
rect 2042 3431 2098 3440
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 2332 3058 2360 5850
rect 2516 5778 2544 6190
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2516 5166 2544 5714
rect 2792 5710 2820 6208
rect 3160 6186 3188 7686
rect 3252 7002 3280 8842
rect 3344 8430 3372 10950
rect 3528 8956 3556 23446
rect 3988 23118 4016 23598
rect 4080 23254 4108 24568
rect 4160 24550 4212 24556
rect 4264 24342 4292 24822
rect 4356 24818 4384 27066
rect 4896 26852 4948 26858
rect 4896 26794 4948 26800
rect 4436 26376 4488 26382
rect 4436 26318 4488 26324
rect 4448 25294 4476 26318
rect 4712 26240 4764 26246
rect 4712 26182 4764 26188
rect 4724 25770 4752 26182
rect 4908 25906 4936 26794
rect 4988 26784 5040 26790
rect 4988 26726 5040 26732
rect 5000 26518 5028 26726
rect 4988 26512 5040 26518
rect 4988 26454 5040 26460
rect 5000 26246 5028 26454
rect 4988 26240 5040 26246
rect 4988 26182 5040 26188
rect 4896 25900 4948 25906
rect 4896 25842 4948 25848
rect 4620 25764 4672 25770
rect 4620 25706 4672 25712
rect 4712 25764 4764 25770
rect 4712 25706 4764 25712
rect 4632 25498 4660 25706
rect 4620 25492 4672 25498
rect 4620 25434 4672 25440
rect 4436 25288 4488 25294
rect 4436 25230 4488 25236
rect 4344 24812 4396 24818
rect 4344 24754 4396 24760
rect 4344 24608 4396 24614
rect 4344 24550 4396 24556
rect 4252 24336 4304 24342
rect 4252 24278 4304 24284
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 4172 23730 4200 24006
rect 4264 23866 4292 24278
rect 4356 24206 4384 24550
rect 4344 24200 4396 24206
rect 4344 24142 4396 24148
rect 4252 23860 4304 23866
rect 4252 23802 4304 23808
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 4068 23248 4120 23254
rect 4068 23190 4120 23196
rect 3976 23112 4028 23118
rect 3976 23054 4028 23060
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 4448 22778 4476 25230
rect 4620 25220 4672 25226
rect 4724 25208 4752 25706
rect 4672 25180 4752 25208
rect 4620 25162 4672 25168
rect 4528 24676 4580 24682
rect 4528 24618 4580 24624
rect 4540 24138 4568 24618
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 4712 24404 4764 24410
rect 4712 24346 4764 24352
rect 4528 24132 4580 24138
rect 4528 24074 4580 24080
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4632 23322 4660 24006
rect 4620 23316 4672 23322
rect 4620 23258 4672 23264
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 4080 22642 4108 22714
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 4252 22636 4304 22642
rect 4252 22578 4304 22584
rect 4160 22500 4212 22506
rect 4160 22442 4212 22448
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3988 20330 4016 21286
rect 4172 21146 4200 22442
rect 4264 22030 4292 22578
rect 4344 22092 4396 22098
rect 4344 22034 4396 22040
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 4160 21140 4212 21146
rect 4160 21082 4212 21088
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3976 20324 4028 20330
rect 3976 20266 4028 20272
rect 4080 19990 4108 20878
rect 4172 20534 4200 20946
rect 4160 20528 4212 20534
rect 4160 20470 4212 20476
rect 4264 20466 4292 21966
rect 4356 21690 4384 22034
rect 4344 21684 4396 21690
rect 4344 21626 4396 21632
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4632 21078 4660 21286
rect 4620 21072 4672 21078
rect 4620 21014 4672 21020
rect 4632 20602 4660 21014
rect 4724 21010 4752 24346
rect 4816 23322 4844 24550
rect 4908 24342 4936 25842
rect 5000 25702 5028 26182
rect 4988 25696 5040 25702
rect 4988 25638 5040 25644
rect 4988 25424 5040 25430
rect 4988 25366 5040 25372
rect 5000 24954 5028 25366
rect 4988 24948 5040 24954
rect 4988 24890 5040 24896
rect 4988 24812 5040 24818
rect 4988 24754 5040 24760
rect 4896 24336 4948 24342
rect 4896 24278 4948 24284
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4160 20324 4212 20330
rect 4160 20266 4212 20272
rect 4068 19984 4120 19990
rect 4068 19926 4120 19932
rect 4172 19786 4200 20266
rect 3976 19780 4028 19786
rect 3976 19722 4028 19728
rect 4160 19780 4212 19786
rect 4160 19722 4212 19728
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3988 19378 4016 19722
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3988 19249 4016 19314
rect 3884 19236 3936 19242
rect 3884 19178 3936 19184
rect 3896 18748 3924 19178
rect 4080 19145 4108 19654
rect 4160 19168 4212 19174
rect 4066 19136 4122 19145
rect 4160 19110 4212 19116
rect 4434 19136 4490 19145
rect 4066 19071 4122 19080
rect 3976 18760 4028 18766
rect 3896 18720 3976 18748
rect 3976 18702 4028 18708
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3988 17241 4016 18702
rect 4172 18426 4200 19110
rect 4434 19071 4490 19080
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 3974 17232 4030 17241
rect 3974 17167 4030 17176
rect 4356 17066 4384 17818
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3896 16726 3924 16934
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 4252 16720 4304 16726
rect 4252 16662 4304 16668
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15638 3924 15846
rect 3988 15706 4016 16526
rect 4264 16250 4292 16662
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 3884 15632 3936 15638
rect 3884 15574 3936 15580
rect 4080 15434 4108 15642
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 4264 13512 4292 15914
rect 4448 14822 4476 19071
rect 4528 18896 4580 18902
rect 4528 18838 4580 18844
rect 4540 18086 4568 18838
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 4540 17882 4568 18022
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4632 17814 4660 20538
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4908 19514 4936 19994
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4816 18766 4844 19246
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4804 18760 4856 18766
rect 4856 18720 4936 18748
rect 4804 18702 4856 18708
rect 4724 18290 4752 18702
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4712 18284 4764 18290
rect 4712 18226 4764 18232
rect 4816 18154 4844 18362
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 4620 17808 4672 17814
rect 4620 17750 4672 17756
rect 4724 17542 4752 18090
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 4816 16794 4844 17070
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4816 15638 4844 16526
rect 4908 16114 4936 18720
rect 5000 16572 5028 24754
rect 5092 23186 5120 28902
rect 5172 27600 5224 27606
rect 5172 27542 5224 27548
rect 5184 26858 5212 27542
rect 5172 26852 5224 26858
rect 5172 26794 5224 26800
rect 5172 26036 5224 26042
rect 5172 25978 5224 25984
rect 5080 23180 5132 23186
rect 5080 23122 5132 23128
rect 5092 22574 5120 23122
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5184 22114 5212 25978
rect 5276 24818 5304 34342
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 5368 27946 5396 28358
rect 5552 28150 5580 39646
rect 5722 39636 5778 40000
rect 6184 39772 6236 39778
rect 6184 39714 6236 39720
rect 5722 39584 5724 39636
rect 5776 39584 5778 39636
rect 5722 39520 5778 39584
rect 5816 39500 5868 39506
rect 5816 39442 5868 39448
rect 5632 33312 5684 33318
rect 5632 33254 5684 33260
rect 5540 28144 5592 28150
rect 5540 28086 5592 28092
rect 5356 27940 5408 27946
rect 5356 27882 5408 27888
rect 5368 26586 5396 27882
rect 5540 27872 5592 27878
rect 5540 27814 5592 27820
rect 5356 26580 5408 26586
rect 5356 26522 5408 26528
rect 5552 26450 5580 27814
rect 5540 26444 5592 26450
rect 5540 26386 5592 26392
rect 5644 26042 5672 33254
rect 5724 28144 5776 28150
rect 5724 28086 5776 28092
rect 5736 27062 5764 28086
rect 5724 27056 5776 27062
rect 5724 26998 5776 27004
rect 5632 26036 5684 26042
rect 5632 25978 5684 25984
rect 5448 25424 5500 25430
rect 5448 25366 5500 25372
rect 5460 24954 5488 25366
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 5448 24948 5500 24954
rect 5448 24890 5500 24896
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5264 24132 5316 24138
rect 5264 24074 5316 24080
rect 5276 23594 5304 24074
rect 5552 24070 5580 25230
rect 5724 24200 5776 24206
rect 5724 24142 5776 24148
rect 5540 24064 5592 24070
rect 5540 24006 5592 24012
rect 5632 23724 5684 23730
rect 5632 23666 5684 23672
rect 5644 23594 5672 23666
rect 5264 23588 5316 23594
rect 5264 23530 5316 23536
rect 5632 23588 5684 23594
rect 5632 23530 5684 23536
rect 5276 23322 5304 23530
rect 5264 23316 5316 23322
rect 5264 23258 5316 23264
rect 5540 23248 5592 23254
rect 5540 23190 5592 23196
rect 5552 22710 5580 23190
rect 5540 22704 5592 22710
rect 5540 22646 5592 22652
rect 5552 22438 5580 22646
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 5552 22234 5580 22374
rect 5644 22234 5672 23530
rect 5736 23526 5764 24142
rect 5724 23520 5776 23526
rect 5724 23462 5776 23468
rect 5736 22642 5764 23462
rect 5828 22982 5856 39442
rect 6092 29776 6144 29782
rect 6092 29718 6144 29724
rect 6000 29640 6052 29646
rect 6000 29582 6052 29588
rect 5908 29300 5960 29306
rect 5908 29242 5960 29248
rect 5816 22976 5868 22982
rect 5816 22918 5868 22924
rect 5920 22778 5948 29242
rect 6012 28762 6040 29582
rect 6104 28966 6132 29718
rect 6196 29238 6224 39714
rect 6550 39704 6606 40000
rect 6550 39652 6552 39704
rect 6604 39652 6606 39704
rect 6550 39520 6606 39652
rect 7470 39636 7526 40000
rect 8390 39658 8446 40000
rect 9218 39658 9274 40000
rect 10138 39658 10194 40000
rect 11058 39658 11114 40000
rect 11886 39658 11942 40000
rect 12806 39658 12862 40000
rect 13726 39658 13782 40000
rect 7470 39584 7472 39636
rect 7524 39584 7526 39636
rect 7470 39520 7526 39584
rect 8024 39636 8076 39642
rect 8024 39578 8076 39584
rect 8128 39630 8446 39658
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 7102 37224 7158 37233
rect 7102 37159 7158 37168
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 7116 29850 7144 37159
rect 7656 35148 7708 35154
rect 7656 35090 7708 35096
rect 7668 34406 7696 35090
rect 7656 34400 7708 34406
rect 7656 34342 7708 34348
rect 7104 29844 7156 29850
rect 7104 29786 7156 29792
rect 7840 29708 7892 29714
rect 7840 29650 7892 29656
rect 7196 29640 7248 29646
rect 7196 29582 7248 29588
rect 6276 29504 6328 29510
rect 6276 29446 6328 29452
rect 6288 29306 6316 29446
rect 6276 29300 6328 29306
rect 6276 29242 6328 29248
rect 6184 29232 6236 29238
rect 6184 29174 6236 29180
rect 6288 29102 6316 29242
rect 7104 29232 7156 29238
rect 7104 29174 7156 29180
rect 6276 29096 6328 29102
rect 6276 29038 6328 29044
rect 6920 29028 6972 29034
rect 6920 28970 6972 28976
rect 6092 28960 6144 28966
rect 6092 28902 6144 28908
rect 6644 28960 6696 28966
rect 6644 28902 6696 28908
rect 6000 28756 6052 28762
rect 6000 28698 6052 28704
rect 6104 28694 6132 28902
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6092 28688 6144 28694
rect 6092 28630 6144 28636
rect 6000 28552 6052 28558
rect 6000 28494 6052 28500
rect 6012 27674 6040 28494
rect 6104 27878 6132 28630
rect 6092 27872 6144 27878
rect 6092 27814 6144 27820
rect 6000 27668 6052 27674
rect 6000 27610 6052 27616
rect 6104 27130 6132 27814
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6656 27538 6684 28902
rect 6932 28762 6960 28970
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 7012 28552 7064 28558
rect 7012 28494 7064 28500
rect 6920 28008 6972 28014
rect 6920 27950 6972 27956
rect 6736 27872 6788 27878
rect 6736 27814 6788 27820
rect 6644 27532 6696 27538
rect 6644 27474 6696 27480
rect 6184 27396 6236 27402
rect 6184 27338 6236 27344
rect 6092 27124 6144 27130
rect 6092 27066 6144 27072
rect 6196 26994 6224 27338
rect 6748 26994 6776 27814
rect 6932 27334 6960 27950
rect 7024 27946 7052 28494
rect 7012 27940 7064 27946
rect 7012 27882 7064 27888
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 6184 26988 6236 26994
rect 6184 26930 6236 26936
rect 6736 26988 6788 26994
rect 6736 26930 6788 26936
rect 6920 26784 6972 26790
rect 6920 26726 6972 26732
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6644 26580 6696 26586
rect 6644 26522 6696 26528
rect 6000 26376 6052 26382
rect 6000 26318 6052 26324
rect 6012 25702 6040 26318
rect 6656 26042 6684 26522
rect 6736 26444 6788 26450
rect 6736 26386 6788 26392
rect 6644 26036 6696 26042
rect 6644 25978 6696 25984
rect 6656 25702 6684 25978
rect 6748 25906 6776 26386
rect 6736 25900 6788 25906
rect 6736 25842 6788 25848
rect 6000 25696 6052 25702
rect 6000 25638 6052 25644
rect 6644 25696 6696 25702
rect 6644 25638 6696 25644
rect 6012 25498 6040 25638
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6000 25492 6052 25498
rect 6000 25434 6052 25440
rect 6736 24812 6788 24818
rect 6788 24772 6868 24800
rect 6736 24754 6788 24760
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6092 24336 6144 24342
rect 6092 24278 6144 24284
rect 6104 23866 6132 24278
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 6000 23588 6052 23594
rect 6000 23530 6052 23536
rect 6012 23050 6040 23530
rect 6104 23322 6132 23802
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6092 23316 6144 23322
rect 6092 23258 6144 23264
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 6000 23044 6052 23050
rect 6000 22986 6052 22992
rect 5908 22772 5960 22778
rect 5908 22714 5960 22720
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 6092 22568 6144 22574
rect 6092 22510 6144 22516
rect 5908 22500 5960 22506
rect 5908 22442 5960 22448
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5632 22228 5684 22234
rect 5632 22170 5684 22176
rect 5184 22086 5488 22114
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5080 21888 5132 21894
rect 5080 21830 5132 21836
rect 5092 21486 5120 21830
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 5184 21078 5212 21966
rect 5172 21072 5224 21078
rect 5172 21014 5224 21020
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 5368 20602 5396 20742
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 5368 19990 5396 20538
rect 5264 19984 5316 19990
rect 5264 19926 5316 19932
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 5276 19718 5304 19926
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5276 19514 5304 19654
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5262 18864 5318 18873
rect 5262 18799 5318 18808
rect 5000 16544 5120 16572
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4620 15632 4672 15638
rect 4620 15574 4672 15580
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4344 14544 4396 14550
rect 4448 14521 4476 14758
rect 4632 14618 4660 15574
rect 4908 15502 4936 16050
rect 5000 15978 5028 16186
rect 4988 15972 5040 15978
rect 4988 15914 5040 15920
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 4988 14544 5040 14550
rect 4344 14486 4396 14492
rect 4434 14512 4490 14521
rect 4356 13938 4384 14486
rect 4988 14486 5040 14492
rect 4434 14447 4490 14456
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4436 14272 4488 14278
rect 4436 14214 4488 14220
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4448 13802 4476 14214
rect 4618 14104 4674 14113
rect 4618 14039 4674 14048
rect 4436 13796 4488 13802
rect 4436 13738 4488 13744
rect 4344 13524 4396 13530
rect 4264 13484 4344 13512
rect 4344 13466 4396 13472
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 3988 12442 4016 13262
rect 4356 12696 4384 13466
rect 4448 13258 4476 13738
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 4436 12708 4488 12714
rect 4356 12668 4436 12696
rect 4436 12650 4488 12656
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 3988 10674 4016 11494
rect 4080 10810 4108 12582
rect 4448 12442 4476 12650
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4264 11354 4292 12242
rect 4448 11898 4476 12378
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4436 11688 4488 11694
rect 4434 11656 4436 11665
rect 4488 11656 4490 11665
rect 4434 11591 4490 11600
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 4080 10520 4108 10746
rect 4448 10674 4476 11591
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4252 10532 4304 10538
rect 4080 10492 4252 10520
rect 4252 10474 4304 10480
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3436 8928 3556 8956
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 3252 6118 3280 6394
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2792 5302 2820 5646
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2412 5092 2464 5098
rect 2412 5034 2464 5040
rect 2424 3534 2452 5034
rect 2516 4826 2544 5102
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2596 4752 2648 4758
rect 2596 4694 2648 4700
rect 2608 3942 2636 4694
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2516 2922 2544 3674
rect 2608 3398 2636 3878
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 2608 2582 2636 3334
rect 2596 2576 2648 2582
rect 2596 2518 2648 2524
rect 2700 2417 2728 3946
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2792 3466 2820 3878
rect 2780 3460 2832 3466
rect 2780 3402 2832 3408
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2792 2650 2820 2858
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2686 2408 2742 2417
rect 2686 2343 2742 2352
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 1780 2106 1808 2246
rect 1768 2100 1820 2106
rect 1768 2042 1820 2048
rect 1492 2032 1544 2038
rect 1492 1974 1544 1980
rect 1032 128 1084 134
rect 1032 70 1084 76
rect 1398 96 1454 480
rect 1504 134 1532 1974
rect 846 8 848 60
rect 900 8 902 60
rect 846 0 902 8
rect 1492 128 1544 134
rect 1492 70 1544 76
rect 2042 128 2098 480
rect 2042 76 2044 128
rect 2096 76 2098 128
rect 1398 0 1454 40
rect 2042 0 2098 76
rect 2594 82 2650 480
rect 2884 82 2912 5578
rect 3344 5250 3372 6666
rect 3436 6458 3464 8928
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3988 8378 4016 10202
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4356 9722 4384 10066
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4080 9178 4108 9454
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4080 8838 4108 9114
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3528 8090 3556 8366
rect 3988 8350 4108 8378
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 8090 4016 8230
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4080 7954 4108 8350
rect 4172 8090 4200 8910
rect 4264 8634 4292 9046
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4264 8294 4292 8570
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3528 6934 3556 7142
rect 3516 6928 3568 6934
rect 3516 6870 3568 6876
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3436 5574 3464 6258
rect 3528 5914 3556 6870
rect 4080 6866 4108 7890
rect 4172 7002 4200 8026
rect 4356 7410 4384 9386
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4264 6662 4292 7142
rect 4356 7002 4384 7346
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4448 6730 4476 8910
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3252 5234 3372 5250
rect 3252 5228 3384 5234
rect 3252 5222 3332 5228
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2976 4010 3004 4966
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2976 3194 3004 3946
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2594 54 2912 82
rect 3160 82 3188 4694
rect 3252 4622 3280 5222
rect 3332 5170 3384 5176
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3344 4486 3372 5034
rect 3332 4480 3384 4486
rect 3332 4422 3384 4428
rect 3436 4154 3464 5510
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3988 5370 4016 5714
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3344 4146 3464 4154
rect 3332 4140 3464 4146
rect 3384 4126 3464 4140
rect 3332 4082 3384 4088
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 3252 2582 3280 2790
rect 3344 2650 3372 4082
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 3436 1601 3464 3334
rect 3528 3194 3556 3470
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3988 3097 4016 4422
rect 3974 3088 4030 3097
rect 3974 3023 4030 3032
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 4080 1834 4108 6394
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4264 5370 4292 5714
rect 4448 5710 4476 6666
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4344 5024 4396 5030
rect 4344 4966 4396 4972
rect 4356 2922 4384 4966
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4448 3534 4476 3674
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4068 1828 4120 1834
rect 4068 1770 4120 1776
rect 3422 1592 3478 1601
rect 3422 1527 3478 1536
rect 3238 82 3294 480
rect 3160 54 3294 82
rect 2594 0 2650 54
rect 3238 0 3294 54
rect 3790 82 3846 480
rect 4080 82 4108 1770
rect 4264 134 4292 2790
rect 3790 54 4108 82
rect 4252 128 4304 134
rect 4252 70 4304 76
rect 4356 82 4384 2858
rect 4540 2514 4568 6054
rect 4632 5030 4660 14039
rect 4724 9722 4752 14350
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4816 13938 4844 14010
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4908 13326 4936 14350
rect 5000 14074 5028 14486
rect 5092 14249 5120 16544
rect 5276 15706 5304 18799
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5276 14958 5304 15642
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5078 14240 5134 14249
rect 5078 14175 5134 14184
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 5000 12442 5028 14010
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5368 13190 5396 13262
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5368 12442 5396 12786
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5000 11898 5028 12378
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5000 11608 5028 11834
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5080 11620 5132 11626
rect 5000 11580 5080 11608
rect 5080 11562 5132 11568
rect 5184 11354 5212 11698
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 4986 11112 5042 11121
rect 4986 11047 5042 11056
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 4908 10062 4936 10678
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4908 8838 4936 9998
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4908 7274 4936 8026
rect 4896 7268 4948 7274
rect 4896 7210 4948 7216
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4724 6254 4752 6326
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4724 4826 4752 5646
rect 5000 5642 5028 11047
rect 5276 10470 5304 11154
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5184 9654 5212 9862
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 5080 8560 5132 8566
rect 5080 8502 5132 8508
rect 5092 8106 5120 8502
rect 5184 8294 5212 8774
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5092 8078 5212 8106
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 4988 5636 5040 5642
rect 4988 5578 5040 5584
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4712 4820 4764 4826
rect 4632 4780 4712 4808
rect 4632 4146 4660 4780
rect 4712 4762 4764 4768
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4434 82 4490 480
rect 4356 54 4490 82
rect 4816 82 4844 4490
rect 4908 3738 4936 4966
rect 5092 4758 5120 6598
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 5092 3942 5120 4694
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5092 3670 5120 3878
rect 5080 3664 5132 3670
rect 4894 3632 4950 3641
rect 5080 3606 5132 3612
rect 4894 3567 4950 3576
rect 4908 3194 4936 3567
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5092 2854 5120 3606
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5092 2582 5120 2790
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 5092 1970 5120 2518
rect 5080 1964 5132 1970
rect 5080 1906 5132 1912
rect 4986 82 5042 480
rect 4816 54 5042 82
rect 5184 66 5212 8078
rect 5276 8022 5304 10406
rect 5356 9512 5408 9518
rect 5460 9489 5488 22086
rect 5552 21418 5580 22170
rect 5920 21690 5948 22442
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5908 21480 5960 21486
rect 5908 21422 5960 21428
rect 5540 21412 5592 21418
rect 5540 21354 5592 21360
rect 5920 21146 5948 21422
rect 6000 21412 6052 21418
rect 6000 21354 6052 21360
rect 5908 21140 5960 21146
rect 5908 21082 5960 21088
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5828 20330 5856 20946
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 5816 20324 5868 20330
rect 5816 20266 5868 20272
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5552 18358 5580 20198
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5644 19174 5672 19790
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5644 18970 5672 19110
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 5540 18352 5592 18358
rect 5540 18294 5592 18300
rect 5630 17776 5686 17785
rect 5630 17711 5686 17720
rect 5644 17678 5672 17711
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5736 17338 5764 19110
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5552 16726 5580 17002
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5736 16726 5764 16934
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 5552 15910 5580 16662
rect 5736 16250 5764 16662
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5736 14822 5764 14894
rect 5724 14816 5776 14822
rect 5724 14758 5776 14764
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5356 9454 5408 9460
rect 5446 9480 5502 9489
rect 5368 8838 5396 9454
rect 5446 9415 5502 9424
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5368 8362 5396 8774
rect 5460 8566 5488 9415
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5368 7886 5396 8298
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5460 7732 5488 8230
rect 5368 7704 5488 7732
rect 5368 5574 5396 7704
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 6934 5488 7142
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5460 6458 5488 6870
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5368 5166 5396 5510
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5368 4622 5396 5102
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5368 4185 5396 4558
rect 5354 4176 5410 4185
rect 5354 4111 5410 4120
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3670 5396 3878
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5276 3058 5304 3538
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5368 2922 5396 3334
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5368 2582 5396 2858
rect 5552 2854 5580 13806
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5644 11694 5672 13738
rect 5724 13456 5776 13462
rect 5724 13398 5776 13404
rect 5736 12646 5764 13398
rect 5724 12640 5776 12646
rect 5724 12582 5776 12588
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5736 11286 5764 12582
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5736 10810 5764 11222
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5630 9344 5686 9353
rect 5630 9279 5686 9288
rect 5644 6458 5672 9279
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5736 8566 5764 8842
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5828 6882 5856 17070
rect 5920 16114 5948 20334
rect 6012 20058 6040 21354
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 6012 17338 6040 17750
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 6012 16250 6040 16526
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6104 16130 6132 22510
rect 6656 22438 6684 23054
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6656 22234 6684 22374
rect 6644 22228 6696 22234
rect 6644 22170 6696 22176
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6196 21010 6224 21286
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6368 19984 6420 19990
rect 6368 19926 6420 19932
rect 6380 19378 6408 19926
rect 6656 19514 6684 20538
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 6656 19310 6684 19450
rect 6184 19304 6236 19310
rect 6184 19246 6236 19252
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6196 18834 6224 19246
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6196 18426 6224 18770
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6748 18358 6776 18770
rect 6736 18352 6788 18358
rect 6736 18294 6788 18300
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6196 17678 6224 18158
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6196 16590 6224 17614
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6656 16250 6684 17206
rect 6748 17202 6776 18294
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6840 17134 6868 24772
rect 6932 24614 6960 26726
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 7024 23322 7052 27882
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 7024 22642 7052 23258
rect 7012 22636 7064 22642
rect 7012 22578 7064 22584
rect 7116 22234 7144 29174
rect 7208 29034 7236 29582
rect 7852 29306 7880 29650
rect 7840 29300 7892 29306
rect 7840 29242 7892 29248
rect 7288 29164 7340 29170
rect 7288 29106 7340 29112
rect 7196 29028 7248 29034
rect 7196 28970 7248 28976
rect 7208 25906 7236 28970
rect 7300 28762 7328 29106
rect 7656 28960 7708 28966
rect 7656 28902 7708 28908
rect 7288 28756 7340 28762
rect 7288 28698 7340 28704
rect 7668 28694 7696 28902
rect 7656 28688 7708 28694
rect 7656 28630 7708 28636
rect 7668 28218 7696 28630
rect 7656 28212 7708 28218
rect 7656 28154 7708 28160
rect 7380 27464 7432 27470
rect 7380 27406 7432 27412
rect 7392 26246 7420 27406
rect 7564 27328 7616 27334
rect 7564 27270 7616 27276
rect 7380 26240 7432 26246
rect 7380 26182 7432 26188
rect 7196 25900 7248 25906
rect 7196 25842 7248 25848
rect 7208 24138 7236 25842
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 7300 24750 7328 25094
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7300 24410 7328 24686
rect 7576 24410 7604 27270
rect 7656 25356 7708 25362
rect 7656 25298 7708 25304
rect 7668 25158 7696 25298
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7852 24614 7880 25230
rect 7840 24608 7892 24614
rect 7840 24550 7892 24556
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 7288 24404 7340 24410
rect 7288 24346 7340 24352
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7196 24132 7248 24138
rect 7196 24074 7248 24080
rect 7300 23474 7328 24346
rect 7472 24268 7524 24274
rect 7472 24210 7524 24216
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7392 23594 7420 24142
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7208 23446 7328 23474
rect 7104 22228 7156 22234
rect 7104 22170 7156 22176
rect 7208 21962 7236 23446
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 7196 21956 7248 21962
rect 7196 21898 7248 21904
rect 7208 21486 7236 21898
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 6920 21344 6972 21350
rect 6920 21286 6972 21292
rect 6932 21078 6960 21286
rect 6920 21072 6972 21078
rect 6920 21014 6972 21020
rect 7208 21010 7236 21422
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6932 20534 6960 20742
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 7196 19440 7248 19446
rect 7196 19382 7248 19388
rect 6828 17128 6880 17134
rect 6826 17096 6828 17105
rect 6880 17096 6882 17105
rect 6826 17031 6882 17040
rect 7208 16658 7236 19382
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 6012 16102 6132 16130
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5920 13938 5948 14894
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 6012 13734 6040 16102
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6288 15026 6316 15506
rect 6748 15162 6776 16526
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6840 16046 6868 16390
rect 7208 16250 7236 16594
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6276 15020 6328 15026
rect 6196 14980 6276 15008
rect 6196 14550 6224 14980
rect 6276 14962 6328 14968
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6184 14544 6236 14550
rect 6104 14504 6184 14532
rect 6104 14074 6132 14504
rect 6184 14486 6236 14492
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6104 13462 6132 13738
rect 6092 13456 6144 13462
rect 6092 13398 6144 13404
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 6012 12374 6040 13194
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 6012 11898 6040 12310
rect 6196 12238 6224 14282
rect 6380 14074 6408 14418
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6564 13870 6592 14418
rect 6840 14278 6868 15982
rect 6932 15434 6960 15982
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 7300 14498 7328 22714
rect 7392 22642 7420 23530
rect 7484 23322 7512 24210
rect 7852 23798 7880 24550
rect 7944 24274 7972 24550
rect 7932 24268 7984 24274
rect 7932 24210 7984 24216
rect 7944 23866 7972 24210
rect 7932 23860 7984 23866
rect 7932 23802 7984 23808
rect 7840 23792 7892 23798
rect 7840 23734 7892 23740
rect 7932 23588 7984 23594
rect 7852 23548 7932 23576
rect 7748 23520 7800 23526
rect 7668 23480 7748 23508
rect 7472 23316 7524 23322
rect 7472 23258 7524 23264
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7484 22166 7512 23258
rect 7472 22160 7524 22166
rect 7472 22102 7524 22108
rect 7380 21616 7432 21622
rect 7380 21558 7432 21564
rect 7392 17746 7420 21558
rect 7484 21146 7512 22102
rect 7668 21690 7696 23480
rect 7748 23462 7800 23468
rect 7852 23254 7880 23548
rect 7932 23530 7984 23536
rect 8036 23497 8064 39578
rect 8128 35290 8156 39630
rect 8390 39520 8446 39630
rect 8864 39630 9274 39658
rect 8116 35284 8168 35290
rect 8116 35226 8168 35232
rect 8300 34536 8352 34542
rect 8300 34478 8352 34484
rect 8116 34060 8168 34066
rect 8116 34002 8168 34008
rect 8128 33318 8156 34002
rect 8116 33312 8168 33318
rect 8116 33254 8168 33260
rect 8312 29510 8340 34478
rect 8864 34202 8892 39630
rect 9218 39520 9274 39630
rect 9784 39630 10194 39658
rect 9404 39568 9456 39574
rect 9404 39510 9456 39516
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 9312 34536 9364 34542
rect 9312 34478 9364 34484
rect 8852 34196 8904 34202
rect 8852 34138 8904 34144
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8300 29504 8352 29510
rect 8300 29446 8352 29452
rect 8484 29504 8536 29510
rect 8484 29446 8536 29452
rect 8496 29034 8524 29446
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8484 29028 8536 29034
rect 8484 28970 8536 28976
rect 8576 29028 8628 29034
rect 8576 28970 8628 28976
rect 8208 28416 8260 28422
rect 8208 28358 8260 28364
rect 8116 27600 8168 27606
rect 8116 27542 8168 27548
rect 8128 26994 8156 27542
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 8128 26518 8156 26930
rect 8116 26512 8168 26518
rect 8116 26454 8168 26460
rect 8128 25702 8156 26454
rect 8116 25696 8168 25702
rect 8116 25638 8168 25644
rect 8128 23594 8156 25638
rect 8116 23588 8168 23594
rect 8116 23530 8168 23536
rect 8022 23488 8078 23497
rect 7944 23446 8022 23474
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7748 23112 7800 23118
rect 7748 23054 7800 23060
rect 7760 21894 7788 23054
rect 7852 22710 7880 23190
rect 7840 22704 7892 22710
rect 7840 22646 7892 22652
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7484 20602 7512 21082
rect 7668 21010 7696 21626
rect 7944 21026 7972 23446
rect 8022 23423 8078 23432
rect 8220 22216 8248 28358
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 8312 27674 8340 27814
rect 8300 27668 8352 27674
rect 8300 27610 8352 27616
rect 8496 27402 8524 28970
rect 8484 27396 8536 27402
rect 8484 27338 8536 27344
rect 8588 26586 8616 28970
rect 9324 28422 9352 34478
rect 9416 28608 9444 39510
rect 9784 34746 9812 39630
rect 10138 39520 10194 39630
rect 10704 39630 11114 39658
rect 10704 34746 10732 39630
rect 11058 39520 11114 39630
rect 11532 39630 11942 39658
rect 9772 34740 9824 34746
rect 9772 34682 9824 34688
rect 10692 34740 10744 34746
rect 10692 34682 10744 34688
rect 10508 34400 10560 34406
rect 10508 34342 10560 34348
rect 10048 30048 10100 30054
rect 10048 29990 10100 29996
rect 9588 28620 9640 28626
rect 9416 28580 9588 28608
rect 9588 28562 9640 28568
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8760 27940 8812 27946
rect 8760 27882 8812 27888
rect 9404 27940 9456 27946
rect 9404 27882 9456 27888
rect 8772 27470 8800 27882
rect 8760 27464 8812 27470
rect 8760 27406 8812 27412
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9416 26858 9444 27882
rect 9600 27878 9628 28562
rect 9680 28416 9732 28422
rect 9680 28358 9732 28364
rect 9588 27872 9640 27878
rect 9588 27814 9640 27820
rect 9692 27674 9720 28358
rect 10060 28218 10088 29990
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 10048 28212 10100 28218
rect 10048 28154 10100 28160
rect 10060 28082 10088 28154
rect 10428 28150 10456 28358
rect 10416 28144 10468 28150
rect 10416 28086 10468 28092
rect 10048 28076 10100 28082
rect 10048 28018 10100 28024
rect 10428 27946 10456 28086
rect 9864 27940 9916 27946
rect 9864 27882 9916 27888
rect 10416 27940 10468 27946
rect 10416 27882 10468 27888
rect 9680 27668 9732 27674
rect 9680 27610 9732 27616
rect 9404 26852 9456 26858
rect 9404 26794 9456 26800
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 8576 26580 8628 26586
rect 8576 26522 8628 26528
rect 8484 26240 8536 26246
rect 8484 26182 8536 26188
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 8312 24750 8340 25094
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 8312 23186 8340 24686
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 7656 21004 7708 21010
rect 7656 20946 7708 20952
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7852 20998 7972 21026
rect 8128 22188 8248 22216
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7484 18358 7512 19382
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 7380 17740 7432 17746
rect 7432 17700 7512 17728
rect 7380 17682 7432 17688
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 16794 7420 17478
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7484 16726 7512 17700
rect 7576 17678 7604 19110
rect 7668 18873 7696 20946
rect 7760 19854 7788 20946
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 7852 19378 7880 20998
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 7944 19922 7972 20878
rect 8024 20392 8076 20398
rect 8128 20380 8156 22188
rect 8404 22098 8432 25298
rect 8496 24614 8524 26182
rect 8668 25764 8720 25770
rect 8668 25706 8720 25712
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8484 24064 8536 24070
rect 8484 24006 8536 24012
rect 8496 23730 8524 24006
rect 8680 23866 8708 25706
rect 8668 23860 8720 23866
rect 8668 23802 8720 23808
rect 8484 23724 8536 23730
rect 8484 23666 8536 23672
rect 8496 23474 8524 23666
rect 8496 23446 8616 23474
rect 8588 23118 8616 23446
rect 8576 23112 8628 23118
rect 8576 23054 8628 23060
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 8392 22092 8444 22098
rect 8392 22034 8444 22040
rect 8220 21350 8248 22034
rect 8588 21894 8616 22510
rect 8680 22506 8708 23802
rect 8772 22642 8800 26726
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 8852 25900 8904 25906
rect 9324 25888 9352 26318
rect 9416 26246 9444 26794
rect 9692 26586 9720 27610
rect 9876 27606 9904 27882
rect 9864 27600 9916 27606
rect 9864 27542 9916 27548
rect 9876 27130 9904 27542
rect 10520 27538 10548 34342
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10612 28082 10640 29106
rect 10600 28076 10652 28082
rect 10600 28018 10652 28024
rect 10508 27532 10560 27538
rect 10508 27474 10560 27480
rect 9956 27396 10008 27402
rect 9956 27338 10008 27344
rect 9864 27124 9916 27130
rect 9864 27066 9916 27072
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 9404 26240 9456 26246
rect 9404 26182 9456 26188
rect 9324 25860 9444 25888
rect 8852 25842 8904 25848
rect 8864 25158 8892 25842
rect 8852 25152 8904 25158
rect 8852 25094 8904 25100
rect 8864 23050 8892 25094
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 9416 23526 9444 25860
rect 9864 25764 9916 25770
rect 9968 25752 9996 27338
rect 10416 27056 10468 27062
rect 10416 26998 10468 27004
rect 9916 25724 9996 25752
rect 9864 25706 9916 25712
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9600 24342 9628 24550
rect 9588 24336 9640 24342
rect 9588 24278 9640 24284
rect 9404 23520 9456 23526
rect 9404 23462 9456 23468
rect 9600 23508 9628 24278
rect 9876 24206 9904 25706
rect 10048 25152 10100 25158
rect 10048 25094 10100 25100
rect 10060 24818 10088 25094
rect 10048 24812 10100 24818
rect 9968 24772 10048 24800
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 9784 23866 9812 24142
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9680 23520 9732 23526
rect 9600 23480 9680 23508
rect 9600 23322 9628 23480
rect 9680 23462 9732 23468
rect 9784 23474 9812 23802
rect 9784 23446 9904 23474
rect 9588 23316 9640 23322
rect 9588 23258 9640 23264
rect 9404 23180 9456 23186
rect 9404 23122 9456 23128
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 8852 23044 8904 23050
rect 8852 22986 8904 22992
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8668 22500 8720 22506
rect 8668 22442 8720 22448
rect 8864 22438 8892 22510
rect 8852 22432 8904 22438
rect 8852 22374 8904 22380
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8496 21350 8524 21830
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8076 20352 8156 20380
rect 8024 20334 8076 20340
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 8128 20058 8156 20198
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 7932 19916 7984 19922
rect 7932 19858 7984 19864
rect 7944 19514 7972 19858
rect 8024 19712 8076 19718
rect 8024 19654 8076 19660
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 8036 19310 8064 19654
rect 8128 19378 8156 19994
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 7654 18864 7710 18873
rect 7654 18799 7710 18808
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7852 17134 7880 17682
rect 8036 17202 8064 19246
rect 8128 18970 8156 19314
rect 8116 18964 8168 18970
rect 8116 18906 8168 18912
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8128 17814 8156 18226
rect 8220 18086 8248 21286
rect 8300 20324 8352 20330
rect 8300 20266 8352 20272
rect 8312 19990 8340 20266
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8392 18352 8444 18358
rect 8392 18294 8444 18300
rect 8404 18154 8432 18294
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8496 17882 8524 18770
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8116 17808 8168 17814
rect 8116 17750 8168 17756
rect 8392 17808 8444 17814
rect 8392 17750 8444 17756
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7576 16998 7604 17070
rect 8404 16998 8432 17750
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7576 15570 7604 15982
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7392 14618 7420 15370
rect 7484 15162 7512 15370
rect 7576 15162 7604 15506
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6840 14006 6868 14214
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6552 13864 6604 13870
rect 6932 13841 6960 13942
rect 6552 13806 6604 13812
rect 6918 13832 6974 13841
rect 6918 13767 6974 13776
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6656 12714 6684 13262
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6644 12708 6696 12714
rect 6644 12650 6696 12656
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6092 12164 6144 12170
rect 6092 12106 6144 12112
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6104 11762 6132 12106
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6012 10266 6040 11086
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 5920 9518 5948 9862
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5920 9042 5948 9454
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5920 8634 5948 8978
rect 6012 8974 6040 9454
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5920 7546 5948 8570
rect 6012 7750 6040 8910
rect 6104 7954 6132 9862
rect 6196 8090 6224 10406
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6656 9382 6684 9998
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5736 6854 5856 6882
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5736 4826 5764 6854
rect 5816 6792 5868 6798
rect 5868 6752 5948 6780
rect 5816 6734 5868 6740
rect 5920 6118 5948 6752
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5736 3738 5764 4626
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5828 4282 5856 4422
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5920 3466 5948 6054
rect 6012 5030 6040 7686
rect 6104 6934 6132 7890
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6196 7410 6224 7686
rect 6380 7478 6408 7754
rect 6564 7546 6592 7890
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6656 7274 6684 9318
rect 6748 9042 6776 13194
rect 6840 12646 6868 13330
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 11132 6868 12582
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6932 11762 6960 12174
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6932 11286 6960 11698
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 6840 11104 6960 11132
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10606 6868 10950
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6840 10130 6868 10542
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6748 7546 6776 7822
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6184 7268 6236 7274
rect 6184 7210 6236 7216
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 6104 5914 6132 6870
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6104 4826 6132 5714
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6196 4154 6224 7210
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6932 6390 6960 11104
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6288 5370 6316 5714
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6656 5302 6684 6054
rect 7024 5352 7052 14486
rect 7300 14470 7420 14498
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7208 11665 7236 11698
rect 7194 11656 7250 11665
rect 7194 11591 7250 11600
rect 7392 11257 7420 14470
rect 7484 14074 7512 15098
rect 7576 14482 7604 15098
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7484 12850 7512 13466
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7378 11248 7434 11257
rect 7378 11183 7434 11192
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7392 10606 7420 11018
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7208 10062 7236 10406
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 9450 7236 9998
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7116 8430 7144 9114
rect 7208 8838 7236 9386
rect 7484 9042 7512 9930
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7208 7750 7236 8774
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7300 8430 7328 8570
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7484 8090 7512 8978
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7116 7274 7144 7686
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7116 7002 7144 7210
rect 7104 6996 7156 7002
rect 7104 6938 7156 6944
rect 7208 5778 7236 7686
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7300 6730 7328 7210
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7269 5568 7321 5574
rect 7321 5516 7328 5556
rect 7269 5510 7328 5516
rect 6932 5324 7052 5352
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6656 4486 6684 5102
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6840 4282 6868 4694
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6104 4126 6224 4154
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 5920 3058 5948 3402
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5356 2576 5408 2582
rect 5356 2518 5408 2524
rect 5722 2544 5778 2553
rect 5540 2508 5592 2514
rect 5722 2479 5778 2488
rect 5540 2450 5592 2456
rect 5552 2038 5580 2450
rect 5736 2446 5764 2479
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 5262 1864 5318 1873
rect 5262 1799 5318 1808
rect 5276 1766 5304 1799
rect 5264 1760 5316 1766
rect 5264 1702 5316 1708
rect 5630 82 5686 480
rect 6012 82 6040 2314
rect 3790 0 3846 54
rect 4434 0 4490 54
rect 4986 0 5042 54
rect 5172 60 5224 66
rect 5172 2 5224 8
rect 5630 54 6040 82
rect 6104 82 6132 4126
rect 6840 3942 6868 4218
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 6288 3194 6316 3606
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6656 3194 6684 3334
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6182 82 6238 480
rect 6104 54 6238 82
rect 6656 82 6684 2790
rect 6734 82 6790 480
rect 6656 54 6790 82
rect 6932 82 6960 5324
rect 7116 5166 7144 5510
rect 7300 5234 7328 5510
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7392 4758 7420 7346
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7484 5166 7512 6802
rect 7576 5914 7604 14282
rect 7668 13394 7696 16186
rect 8220 15910 8248 16594
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7760 14958 7788 15438
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 7944 14482 7972 14826
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 7944 14074 7972 14418
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 7760 13569 7788 14010
rect 7932 13796 7984 13802
rect 7932 13738 7984 13744
rect 7746 13560 7802 13569
rect 7746 13495 7802 13504
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7668 11150 7696 11562
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7760 11082 7788 12174
rect 7852 12102 7880 13330
rect 7944 12714 7972 13738
rect 8024 13728 8076 13734
rect 8024 13670 8076 13676
rect 7932 12708 7984 12714
rect 7932 12650 7984 12656
rect 7944 12374 7972 12650
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7944 11558 7972 12310
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7944 11286 7972 11494
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7852 10674 7880 11086
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7668 5794 7696 10134
rect 7944 9178 7972 10746
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7852 7478 7880 8502
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7944 7954 7972 8230
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7944 7546 7972 7890
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7760 6118 7788 6802
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7576 5766 7696 5794
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7024 3398 7052 4082
rect 7116 3466 7144 4082
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7392 3398 7420 4694
rect 7576 4554 7604 5766
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7576 3738 7604 4150
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7024 2582 7052 3334
rect 7392 3126 7420 3334
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7576 3058 7604 3674
rect 7668 3126 7696 5034
rect 7760 4826 7788 5578
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7116 2582 7144 2790
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7116 2310 7144 2518
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7760 2106 7788 3402
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 7378 82 7434 480
rect 6932 54 7434 82
rect 7852 82 7880 7414
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7944 5710 7972 6054
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7944 5030 7972 5646
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7944 4214 7972 4966
rect 8036 4758 8064 13670
rect 8128 11694 8156 15370
rect 8220 15094 8248 15846
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8208 15088 8260 15094
rect 8208 15030 8260 15036
rect 8312 14822 8340 15302
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8312 13802 8340 14758
rect 8404 14521 8432 16934
rect 8390 14512 8446 14521
rect 8390 14447 8446 14456
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8300 13796 8352 13802
rect 8300 13738 8352 13744
rect 8404 13462 8432 14350
rect 8588 14346 8616 21490
rect 8864 21486 8892 22374
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8680 21078 8708 21422
rect 8864 21146 8892 21422
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 8668 21072 8720 21078
rect 8668 21014 8720 21020
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 8772 20058 8800 20198
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 9324 19922 9352 21830
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8772 18834 8800 19178
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8680 16522 8708 17070
rect 8668 16516 8720 16522
rect 8668 16458 8720 16464
rect 8772 15450 8800 18634
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8864 18290 8892 18566
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 9324 18154 9352 19110
rect 9416 18834 9444 23122
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9312 18148 9364 18154
rect 9312 18090 9364 18096
rect 9404 18080 9456 18086
rect 9404 18022 9456 18028
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8680 15422 8800 15450
rect 8680 14550 8708 15422
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8772 15026 8800 15302
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8574 14240 8630 14249
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8496 11898 8524 14214
rect 8574 14175 8630 14184
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8128 11558 8156 11630
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 10130 8156 11494
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8220 9586 8248 10202
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8128 9110 8156 9318
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8128 8634 8156 9046
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8128 7274 8156 8298
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8312 6866 8340 10678
rect 8404 10470 8432 11222
rect 8496 10606 8524 11834
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 9450 8432 10406
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 8294 8432 8774
rect 8496 8498 8524 8910
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8220 6186 8248 6666
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8220 5642 8248 6122
rect 8208 5636 8260 5642
rect 8404 5624 8432 6190
rect 8484 5636 8536 5642
rect 8404 5596 8484 5624
rect 8208 5578 8260 5584
rect 8484 5578 8536 5584
rect 8496 5302 8524 5578
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8404 4758 8432 5102
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8036 4282 8064 4694
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 7932 4208 7984 4214
rect 7932 4150 7984 4156
rect 8036 3913 8064 4218
rect 8128 4010 8156 4558
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8404 4049 8432 4422
rect 8390 4040 8446 4049
rect 8116 4004 8168 4010
rect 8390 3975 8446 3984
rect 8116 3946 8168 3952
rect 8022 3904 8078 3913
rect 8022 3839 8078 3848
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 7944 3194 7972 3606
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 7932 3188 7984 3194
rect 7932 3130 7984 3136
rect 8312 2922 8340 3470
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 8312 2106 8340 2246
rect 8300 2100 8352 2106
rect 8300 2042 8352 2048
rect 7930 82 7986 480
rect 7852 54 7986 82
rect 8496 82 8524 4966
rect 8588 2514 8616 14175
rect 8680 12986 8708 14350
rect 8864 14006 8892 16934
rect 9232 16504 9260 17138
rect 9324 17134 9352 17478
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9312 16516 9364 16522
rect 9232 16476 9312 16504
rect 9312 16458 9364 16464
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 9220 16108 9272 16114
rect 9324 16096 9352 16458
rect 9272 16068 9352 16096
rect 9220 16050 9272 16056
rect 9232 15638 9260 16050
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8956 14550 8984 14758
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8772 13530 8800 13874
rect 9416 13814 9444 18022
rect 9508 17814 9536 21830
rect 9692 21690 9720 22034
rect 9784 21894 9812 23122
rect 9876 22030 9904 23446
rect 9968 22234 9996 24772
rect 10048 24754 10100 24760
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 10060 23186 10088 23598
rect 10048 23180 10100 23186
rect 10048 23122 10100 23128
rect 10060 22438 10088 23122
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 10060 21962 10088 22374
rect 10428 22114 10456 26998
rect 10612 26994 10640 28018
rect 11244 27532 11296 27538
rect 11244 27474 11296 27480
rect 11256 27130 11284 27474
rect 11244 27124 11296 27130
rect 11244 27066 11296 27072
rect 10600 26988 10652 26994
rect 10600 26930 10652 26936
rect 10692 26240 10744 26246
rect 10692 26182 10744 26188
rect 10704 24682 10732 26182
rect 10968 25356 11020 25362
rect 10968 25298 11020 25304
rect 10980 24954 11008 25298
rect 10968 24948 11020 24954
rect 10968 24890 11020 24896
rect 10692 24676 10744 24682
rect 10692 24618 10744 24624
rect 10704 22642 10732 24618
rect 11532 24410 11560 39630
rect 11886 39520 11942 39630
rect 12544 39630 12862 39658
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 12544 34610 12572 39630
rect 12806 39520 12862 39630
rect 13464 39630 13782 39658
rect 14554 39658 14610 40000
rect 13464 34678 13492 39630
rect 13726 39520 13782 39630
rect 13820 39636 13872 39642
rect 13820 39578 13872 39584
rect 14554 39630 14688 39658
rect 13452 34672 13504 34678
rect 13452 34614 13504 34620
rect 12532 34604 12584 34610
rect 12532 34546 12584 34552
rect 11980 34536 12032 34542
rect 11980 34478 12032 34484
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11992 28529 12020 34478
rect 12714 30016 12770 30025
rect 12714 29951 12770 29960
rect 11978 28520 12034 28529
rect 11978 28455 12034 28464
rect 12072 27872 12124 27878
rect 12072 27814 12124 27820
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11978 24848 12034 24857
rect 11978 24783 12034 24792
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11520 24404 11572 24410
rect 11520 24346 11572 24352
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 11256 23662 11284 24210
rect 11520 24064 11572 24070
rect 11520 24006 11572 24012
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 11334 23488 11390 23497
rect 10980 23322 11008 23462
rect 11334 23423 11390 23432
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 10980 22710 11008 23258
rect 11348 23186 11376 23423
rect 11336 23180 11388 23186
rect 11336 23122 11388 23128
rect 10968 22704 11020 22710
rect 10968 22646 11020 22652
rect 10692 22636 10744 22642
rect 10692 22578 10744 22584
rect 10508 22500 10560 22506
rect 10508 22442 10560 22448
rect 10520 22234 10548 22442
rect 11348 22438 11376 23122
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 10508 22228 10560 22234
rect 10508 22170 10560 22176
rect 10428 22086 10548 22114
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9680 21684 9732 21690
rect 9600 21644 9680 21672
rect 9600 17882 9628 21644
rect 9680 21626 9732 21632
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9876 20602 9904 21014
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 9784 20058 9812 20334
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9692 19514 9720 19858
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9784 19174 9812 19858
rect 9968 19718 9996 20878
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10428 20466 10456 20742
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10048 19984 10100 19990
rect 10048 19926 10100 19932
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9784 18834 9812 19110
rect 9772 18828 9824 18834
rect 9692 18788 9772 18816
rect 9692 18086 9720 18788
rect 9772 18770 9824 18776
rect 9772 18216 9824 18222
rect 9772 18158 9824 18164
rect 9784 18086 9812 18158
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9692 17898 9720 18022
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9692 17870 9812 17898
rect 9496 17808 9548 17814
rect 9496 17750 9548 17756
rect 9588 17740 9640 17746
rect 9692 17728 9720 17870
rect 9640 17700 9720 17728
rect 9588 17682 9640 17688
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9600 16114 9628 16390
rect 9692 16114 9720 16594
rect 9784 16504 9812 17870
rect 9876 17814 9904 18090
rect 9864 17808 9916 17814
rect 9968 17785 9996 19450
rect 10060 19378 10088 19926
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 10428 18698 10456 20402
rect 10520 19428 10548 22086
rect 10692 22092 10744 22098
rect 10692 22034 10744 22040
rect 10704 21554 10732 22034
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10612 20330 10640 20878
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 10612 19786 10640 20266
rect 10796 19961 10824 20742
rect 11072 20262 11100 20946
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10782 19952 10838 19961
rect 10782 19887 10838 19896
rect 10600 19780 10652 19786
rect 10600 19722 10652 19728
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10600 19440 10652 19446
rect 10520 19400 10600 19428
rect 10600 19382 10652 19388
rect 10508 19236 10560 19242
rect 10508 19178 10560 19184
rect 10520 18970 10548 19178
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 9864 17750 9916 17756
rect 9954 17776 10010 17785
rect 9876 17338 9904 17750
rect 10428 17746 10456 18634
rect 9954 17711 10010 17720
rect 10416 17740 10468 17746
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9968 17218 9996 17711
rect 10416 17682 10468 17688
rect 10048 17672 10100 17678
rect 10048 17614 10100 17620
rect 10060 17338 10088 17614
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 9968 17190 10088 17218
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9968 16658 9996 17070
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9864 16516 9916 16522
rect 9784 16476 9864 16504
rect 9864 16458 9916 16464
rect 9968 16250 9996 16594
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9508 15638 9536 15914
rect 9600 15706 9628 16050
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9496 15632 9548 15638
rect 9496 15574 9548 15580
rect 9692 15434 9720 16050
rect 9968 15638 9996 16186
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9876 15162 9904 15574
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9784 14618 9812 14894
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9588 14544 9640 14550
rect 9588 14486 9640 14492
rect 9600 14074 9628 14486
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9324 13786 9444 13814
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 9324 12345 9352 13786
rect 9494 13696 9550 13705
rect 9494 13631 9550 13640
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9310 12336 9366 12345
rect 9310 12271 9366 12280
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8680 10674 8708 11698
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8668 10668 8720 10674
rect 8668 10610 8720 10616
rect 8772 10606 8800 10950
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 9324 10198 9352 12271
rect 9416 11354 9444 12378
rect 9508 11898 9536 13631
rect 9692 13530 9720 14282
rect 9968 14278 9996 15438
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9876 13734 9904 14010
rect 10060 13841 10088 17190
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10244 13938 10272 15914
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 14550 10456 15438
rect 10416 14544 10468 14550
rect 10336 14504 10416 14532
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10046 13832 10102 13841
rect 9956 13796 10008 13802
rect 10230 13832 10286 13841
rect 10046 13767 10102 13776
rect 10140 13796 10192 13802
rect 9956 13738 10008 13744
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9968 13462 9996 13738
rect 10060 13705 10088 13767
rect 10230 13767 10286 13776
rect 10140 13738 10192 13744
rect 10046 13696 10102 13705
rect 10046 13631 10102 13640
rect 10152 13530 10180 13738
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9784 12986 9812 13262
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9784 12374 9812 12922
rect 9876 12646 9904 13398
rect 10244 13258 10272 13767
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10232 12708 10284 12714
rect 10336 12696 10364 14504
rect 10416 14486 10468 14492
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10428 13326 10456 13874
rect 10612 13814 10640 19382
rect 10796 19310 10824 19654
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10704 17202 10732 18226
rect 10796 18204 10824 19246
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10888 18426 10916 18702
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10980 18222 11008 18838
rect 10876 18216 10928 18222
rect 10796 18176 10876 18204
rect 10876 18158 10928 18164
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10888 17610 10916 18158
rect 10876 17604 10928 17610
rect 10876 17546 10928 17552
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10796 17241 10824 17478
rect 10782 17232 10838 17241
rect 10692 17196 10744 17202
rect 10782 17167 10838 17176
rect 10692 17138 10744 17144
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10888 16697 10916 17070
rect 10968 16720 11020 16726
rect 10874 16688 10930 16697
rect 10968 16662 11020 16668
rect 10874 16623 10930 16632
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10520 13786 10640 13814
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10284 12668 10364 12696
rect 10232 12650 10284 12656
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 10244 12238 10272 12650
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9508 11150 9536 11494
rect 9600 11286 9628 12174
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9876 11354 9904 12038
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9508 10470 9536 11086
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 9508 8514 9536 10406
rect 9784 10266 9812 11290
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9968 10810 9996 11154
rect 10060 11082 10088 11494
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 9956 10532 10008 10538
rect 9956 10474 10008 10480
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9968 10198 9996 10474
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9600 9110 9628 9998
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9692 9178 9720 9930
rect 9968 9722 9996 10134
rect 10152 9994 10180 10542
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 10060 9450 10088 9862
rect 10152 9450 10180 9930
rect 10336 9586 10364 9930
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9876 9110 9904 9318
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9600 8634 9628 9046
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9508 8486 9628 8514
rect 10060 8498 10088 9386
rect 10428 9042 10456 12310
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10428 8498 10456 8978
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8772 6254 8800 6598
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8680 5166 8708 5714
rect 8772 5166 8800 6190
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8680 4282 8708 5102
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8864 4214 8892 6122
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8956 5846 8984 6054
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 9140 5642 9168 6190
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 9324 5574 9352 7210
rect 9508 7002 9536 7890
rect 9600 7002 9628 8486
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9784 8022 9812 8230
rect 10060 8090 10088 8298
rect 10048 8084 10100 8090
rect 10520 8072 10548 13786
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10048 8026 10100 8032
rect 10428 8044 10548 8072
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9784 7342 9812 7754
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9324 5370 9352 5510
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9324 5030 9352 5306
rect 9416 5234 9444 5714
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9416 4758 9444 5170
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 8852 4208 8904 4214
rect 8852 4150 8904 4156
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8680 1222 8708 2246
rect 8668 1216 8720 1222
rect 8668 1158 8720 1164
rect 8574 82 8630 480
rect 8496 54 8630 82
rect 8772 82 8800 4014
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 9324 1601 9352 3334
rect 9508 2961 9536 6258
rect 9784 5370 9812 7278
rect 10140 7268 10192 7274
rect 10140 7210 10192 7216
rect 10152 7002 10180 7210
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10048 6384 10100 6390
rect 10048 6326 10100 6332
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9968 5778 9996 6122
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9968 5370 9996 5714
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9968 4486 9996 5102
rect 10060 4690 10088 6326
rect 10152 6118 10180 6802
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10152 5914 10180 6054
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 10152 5302 10180 5578
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9862 4176 9918 4185
rect 9968 4154 9996 4422
rect 10060 4282 10088 4626
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9968 4126 10088 4154
rect 9862 4111 9918 4120
rect 9876 3738 9904 4111
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9494 2952 9550 2961
rect 9494 2887 9550 2896
rect 10060 2650 10088 4126
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9876 2378 9904 2450
rect 9864 2372 9916 2378
rect 9864 2314 9916 2320
rect 9310 1592 9366 1601
rect 9310 1527 9366 1536
rect 9126 82 9182 480
rect 8772 54 9182 82
rect 5630 0 5686 54
rect 6182 0 6238 54
rect 6734 0 6790 54
rect 7378 0 7434 54
rect 7930 0 7986 54
rect 8574 0 8630 54
rect 9126 0 9182 54
rect 9770 82 9826 480
rect 10152 82 10180 5238
rect 10244 5166 10272 5510
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10244 4185 10272 4626
rect 10230 4176 10286 4185
rect 10230 4111 10286 4120
rect 10336 3602 10364 5510
rect 10428 4078 10456 8044
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10520 7206 10548 7890
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10520 7002 10548 7142
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10336 3194 10364 3538
rect 10612 3194 10640 13670
rect 10704 10742 10732 15914
rect 10888 12306 10916 16526
rect 10980 16250 11008 16662
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10980 14550 11008 16186
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 11072 13841 11100 20198
rect 11428 19984 11480 19990
rect 11428 19926 11480 19932
rect 11440 19242 11468 19926
rect 11532 19310 11560 24006
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11428 19236 11480 19242
rect 11428 19178 11480 19184
rect 11624 19156 11652 19722
rect 11716 19514 11744 19790
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11532 19128 11652 19156
rect 11428 18896 11480 18902
rect 11428 18838 11480 18844
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11348 17814 11376 18566
rect 11440 18358 11468 18838
rect 11532 18698 11560 19128
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11520 18692 11572 18698
rect 11520 18634 11572 18640
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11440 17814 11468 18294
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 11428 17808 11480 17814
rect 11428 17750 11480 17756
rect 11348 17338 11376 17750
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11440 17202 11468 17750
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11518 17096 11574 17105
rect 11518 17031 11574 17040
rect 11532 16726 11560 17031
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11520 16720 11572 16726
rect 11520 16662 11572 16668
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11256 15978 11284 16594
rect 11244 15972 11296 15978
rect 11244 15914 11296 15920
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11348 14822 11376 15302
rect 11440 15162 11468 15506
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11532 14482 11560 14894
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11702 14512 11758 14521
rect 11520 14476 11572 14482
rect 11702 14447 11704 14456
rect 11520 14418 11572 14424
rect 11756 14447 11758 14456
rect 11704 14418 11756 14424
rect 11532 14074 11560 14418
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11624 14074 11652 14214
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11058 13832 11114 13841
rect 11058 13767 11114 13776
rect 11164 13569 11192 14010
rect 11716 13938 11744 14418
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11348 13734 11376 13874
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11150 13560 11206 13569
rect 11622 13552 11918 13572
rect 11150 13495 11206 13504
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10782 12200 10838 12209
rect 10782 12135 10838 12144
rect 10796 10810 10824 12135
rect 10888 11558 10916 12242
rect 10980 11801 11008 12718
rect 10966 11792 11022 11801
rect 10966 11727 11022 11736
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10704 9042 10732 9386
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10796 8974 10824 9862
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10704 3641 10732 3946
rect 10690 3632 10746 3641
rect 10690 3567 10746 3576
rect 10796 3505 10824 4422
rect 10782 3496 10838 3505
rect 10782 3431 10838 3440
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10612 2990 10640 3130
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 9770 54 10180 82
rect 10244 82 10272 1906
rect 10322 82 10378 480
rect 10244 54 10378 82
rect 10704 82 10732 3062
rect 10888 3058 10916 11494
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11072 10470 11100 11154
rect 11164 11150 11192 13495
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11348 12442 11376 13262
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11440 12374 11468 13262
rect 11808 12918 11836 13398
rect 11992 13326 12020 24783
rect 12084 18290 12112 27814
rect 12348 27124 12400 27130
rect 12348 27066 12400 27072
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12072 18148 12124 18154
rect 12072 18090 12124 18096
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11992 12442 12020 13126
rect 12084 12782 12112 18090
rect 12176 17134 12204 23462
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 12070 12336 12126 12345
rect 12070 12271 12126 12280
rect 12084 12238 12112 12271
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12084 11898 12112 12174
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10968 9104 11020 9110
rect 10968 9046 11020 9052
rect 10980 8634 11008 9046
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10980 2514 11008 6394
rect 11072 5098 11100 10406
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11256 9489 11284 10066
rect 11242 9480 11298 9489
rect 11242 9415 11298 9424
rect 11256 9382 11284 9415
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 11256 7954 11284 8502
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11256 7546 11284 7890
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11256 4078 11284 4626
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11164 3602 11192 4014
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11164 3194 11192 3538
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 11164 2417 11192 2926
rect 11150 2408 11206 2417
rect 11150 2343 11206 2352
rect 10966 82 11022 480
rect 10704 54 11022 82
rect 11348 82 11376 4218
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11440 3913 11468 4014
rect 11426 3904 11482 3913
rect 11426 3839 11482 3848
rect 11532 2990 11560 9318
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 12084 5574 12112 11630
rect 12176 11121 12204 12718
rect 12162 11112 12218 11121
rect 12162 11047 12218 11056
rect 12268 10266 12296 19246
rect 12360 18222 12388 27066
rect 12728 24070 12756 29951
rect 13832 25498 13860 39578
rect 14554 39520 14610 39630
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14660 34746 14688 39630
rect 15474 39636 15530 40000
rect 15474 39584 15476 39636
rect 15528 39584 15530 39636
rect 15474 39520 15530 39584
rect 14648 34740 14700 34746
rect 14648 34682 14700 34688
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 13820 25492 13872 25498
rect 13820 25434 13872 25440
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12348 18216 12400 18222
rect 12348 18158 12400 18164
rect 12452 15570 12480 22374
rect 12992 20528 13044 20534
rect 12992 20470 13044 20476
rect 13004 20058 13032 20470
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12636 19242 12664 19858
rect 12624 19236 12676 19242
rect 12544 19196 12624 19224
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12176 8498 12204 8978
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12360 8430 12388 13262
rect 12438 10024 12494 10033
rect 12438 9959 12494 9968
rect 12452 8974 12480 9959
rect 12544 9654 12572 19196
rect 12624 19178 12676 19184
rect 13280 18834 13308 22918
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 13268 18828 13320 18834
rect 13268 18770 13320 18776
rect 13280 18426 13308 18770
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 13268 18420 13320 18426
rect 13188 18380 13268 18408
rect 12900 17128 12952 17134
rect 12900 17070 12952 17076
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12636 16250 12664 16594
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12728 14550 12756 14894
rect 12716 14544 12768 14550
rect 12716 14486 12768 14492
rect 12912 13938 12940 17070
rect 13188 16590 13216 18380
rect 13268 18362 13320 18368
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13924 18086 13952 18226
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 13280 17338 13308 17682
rect 13372 17678 13400 18022
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13280 14482 13308 17274
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13464 14822 13492 15506
rect 13452 14816 13504 14822
rect 13452 14758 13504 14764
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13280 14074 13308 14418
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12912 13734 12940 13874
rect 13084 13796 13136 13802
rect 13084 13738 13136 13744
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 12912 12782 12940 13670
rect 13004 13530 13032 13670
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 13096 11898 13124 13738
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13464 11694 13492 14758
rect 13740 14385 13768 17070
rect 13726 14376 13782 14385
rect 13726 14311 13782 14320
rect 13924 12986 13952 18022
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13924 12782 13952 12922
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 9722 12664 9998
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12348 8424 12400 8430
rect 12348 8366 12400 8372
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12268 8090 12296 8230
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 12164 4208 12216 4214
rect 12164 4154 12216 4156
rect 12360 4154 12388 8366
rect 13740 6458 13768 12718
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 12164 4150 12388 4154
rect 12176 4126 12388 4150
rect 12072 4004 12124 4010
rect 12072 3946 12124 3952
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11992 3670 12020 3878
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 12084 3602 12112 3946
rect 12176 3602 12204 4126
rect 14186 4040 14242 4049
rect 14186 3975 14242 3984
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 12176 3194 12204 3538
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12268 3097 12296 3130
rect 12440 3120 12492 3126
rect 12254 3088 12310 3097
rect 12440 3062 12492 3068
rect 12254 3023 12310 3032
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 11992 2553 12020 2790
rect 11978 2544 12034 2553
rect 11978 2479 12034 2488
rect 11518 82 11574 480
rect 11348 54 11574 82
rect 9770 0 9826 54
rect 10322 0 10378 54
rect 10966 0 11022 54
rect 11518 0 11574 54
rect 12070 128 12126 480
rect 12070 76 12072 128
rect 12124 76 12126 128
rect 12070 0 12126 76
rect 12452 82 12480 3062
rect 13280 2854 13308 3538
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13280 2514 13308 2790
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 12544 2009 12572 2450
rect 13360 2372 13412 2378
rect 13360 2314 13412 2320
rect 12530 2000 12586 2009
rect 12530 1935 12586 1944
rect 12714 82 12770 480
rect 12452 54 12770 82
rect 12714 0 12770 54
rect 13266 82 13322 480
rect 13372 82 13400 2314
rect 13832 1873 13860 2926
rect 13818 1864 13874 1873
rect 13818 1799 13874 1808
rect 13728 1216 13780 1222
rect 13728 1158 13780 1164
rect 13266 54 13400 82
rect 13740 82 13768 1158
rect 13910 82 13966 480
rect 13740 54 13966 82
rect 14200 82 14228 3975
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14462 82 14518 480
rect 14200 54 14518 82
rect 13266 0 13322 54
rect 13910 0 13966 54
rect 14462 0 14518 54
rect 15106 82 15162 480
rect 15212 82 15240 3402
rect 15106 54 15240 82
rect 15658 82 15714 480
rect 15764 82 15792 3674
rect 15658 54 15792 82
rect 15106 0 15162 54
rect 15658 0 15714 54
<< via2 >>
rect 1030 31864 1086 31920
rect 1122 26832 1178 26888
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 1306 22208 1362 22264
rect 1306 16904 1362 16960
rect 2318 24792 2374 24848
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3974 28464 4030 28520
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 1950 18808 2006 18864
rect 1030 11736 1086 11792
rect 1306 6976 1362 7032
rect 1582 10140 1584 10160
rect 1584 10140 1636 10160
rect 1636 10140 1638 10160
rect 1582 10104 1638 10140
rect 2962 19896 3018 19952
rect 2502 13776 2558 13832
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 2778 13776 2834 13832
rect 1950 9424 2006 9480
rect 3238 10104 3294 10160
rect 2042 3440 2098 3496
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 4066 19080 4122 19136
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 4434 19080 4490 19136
rect 3974 17176 4030 17232
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 7102 37168 7158 37224
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 5262 18808 5318 18864
rect 4434 14456 4490 14512
rect 4618 14048 4674 14104
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 4434 11636 4436 11656
rect 4436 11636 4488 11656
rect 4488 11636 4490 11656
rect 4434 11600 4490 11636
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 2686 2352 2742 2408
rect 1398 40 1454 96
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 3974 3032 4030 3088
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 3422 1536 3478 1592
rect 5078 14184 5134 14240
rect 4986 11056 5042 11112
rect 4894 3576 4950 3632
rect 5630 17720 5686 17776
rect 5446 9424 5502 9480
rect 5354 4120 5410 4176
rect 5630 9288 5686 9344
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6826 17076 6828 17096
rect 6828 17076 6880 17096
rect 6880 17076 6882 17096
rect 6826 17040 6882 17076
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8022 23432 8078 23488
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 7654 18808 7710 18864
rect 6918 13776 6974 13832
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 7194 11600 7250 11656
rect 7378 11192 7434 11248
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 5722 2488 5778 2544
rect 5262 1808 5318 1864
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 7746 13504 7802 13560
rect 8390 14456 8446 14512
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8574 14184 8630 14240
rect 8390 3984 8446 4040
rect 8022 3848 8078 3904
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 12714 29960 12770 30016
rect 11978 28464 12034 28520
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11978 24792 12034 24848
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11334 23432 11390 23488
rect 10782 19896 10838 19952
rect 9954 17720 10010 17776
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 9494 13640 9550 13696
rect 9310 12280 9366 12336
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 10046 13776 10102 13832
rect 10230 13776 10286 13832
rect 10046 13640 10102 13696
rect 10782 17176 10838 17232
rect 10874 16632 10930 16688
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 9862 4120 9918 4176
rect 9494 2896 9550 2952
rect 9310 1536 9366 1592
rect 10230 4120 10286 4176
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11518 17040 11574 17096
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11702 14476 11758 14512
rect 11702 14456 11704 14476
rect 11704 14456 11756 14476
rect 11756 14456 11758 14476
rect 11058 13776 11114 13832
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11150 13504 11206 13560
rect 10782 12144 10838 12200
rect 10966 11736 11022 11792
rect 10690 3576 10746 3632
rect 10782 3440 10838 3496
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 12070 12280 12126 12336
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11242 9424 11298 9480
rect 11150 2352 11206 2408
rect 11426 3848 11482 3904
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 12162 11056 12218 11112
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 12438 9968 12494 10024
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 13726 14320 13782 14376
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 14186 3984 14242 4040
rect 12254 3032 12310 3088
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 11978 2488 12034 2544
rect 12530 1944 12586 2000
rect 13818 1808 13874 1864
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
<< metal3 >>
rect 6277 37568 6597 37569
rect 0 37408 480 37528
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 62 37226 122 37408
rect 7097 37226 7163 37229
rect 62 37224 7163 37226
rect 62 37168 7102 37224
rect 7158 37168 7163 37224
rect 62 37166 7163 37168
rect 7097 37163 7163 37166
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 0 32376 480 32496
rect 62 31922 122 32376
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 1025 31922 1091 31925
rect 62 31920 1091 31922
rect 62 31864 1030 31920
rect 1086 31864 1091 31920
rect 62 31862 1091 31864
rect 1025 31859 1091 31862
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 12709 30018 12775 30021
rect 15520 30018 16000 30048
rect 12709 30016 16000 30018
rect 12709 29960 12714 30016
rect 12770 29960 16000 30016
rect 12709 29958 16000 29960
rect 12709 29955 12775 29958
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 15520 29928 16000 29958
rect 11610 29887 11930 29888
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 3969 28522 4035 28525
rect 5758 28522 5764 28524
rect 3969 28520 5764 28522
rect 3969 28464 3974 28520
rect 4030 28464 5764 28520
rect 3969 28462 5764 28464
rect 3969 28459 4035 28462
rect 5758 28460 5764 28462
rect 5828 28522 5834 28524
rect 11973 28522 12039 28525
rect 5828 28520 12039 28522
rect 5828 28464 11978 28520
rect 12034 28464 12039 28520
rect 5828 28462 12039 28464
rect 5828 28460 5834 28462
rect 11973 28459 12039 28462
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 0 27344 480 27464
rect 62 26890 122 27344
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 1117 26890 1183 26893
rect 62 26888 1183 26890
rect 62 26832 1122 26888
rect 1178 26832 1183 26888
rect 62 26830 1183 26832
rect 1117 26827 1183 26830
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 2313 24850 2379 24853
rect 11973 24850 12039 24853
rect 2313 24848 12039 24850
rect 2313 24792 2318 24848
rect 2374 24792 11978 24848
rect 12034 24792 12039 24848
rect 2313 24790 12039 24792
rect 2313 24787 2379 24790
rect 11973 24787 12039 24790
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 8017 23490 8083 23493
rect 11329 23490 11395 23493
rect 8017 23488 11395 23490
rect 8017 23432 8022 23488
rect 8078 23432 11334 23488
rect 11390 23432 11395 23488
rect 8017 23430 11395 23432
rect 8017 23427 8083 23430
rect 11329 23427 11395 23430
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 0 22448 480 22568
rect 62 22266 122 22448
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 1301 22266 1367 22269
rect 62 22264 1367 22266
rect 62 22208 1306 22264
rect 1362 22208 1367 22264
rect 62 22206 1367 22208
rect 1301 22203 1367 22206
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 2957 19954 3023 19957
rect 10777 19954 10843 19957
rect 2957 19952 10843 19954
rect 2957 19896 2962 19952
rect 3018 19896 10782 19952
rect 10838 19896 10843 19952
rect 2957 19894 10843 19896
rect 2957 19891 3023 19894
rect 10777 19891 10843 19894
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 4061 19138 4127 19141
rect 4429 19138 4495 19141
rect 4061 19136 4495 19138
rect 4061 19080 4066 19136
rect 4122 19080 4434 19136
rect 4490 19080 4495 19136
rect 4061 19078 4495 19080
rect 4061 19075 4127 19078
rect 4429 19075 4495 19078
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 1945 18866 2011 18869
rect 5257 18866 5323 18869
rect 7649 18866 7715 18869
rect 1945 18864 7715 18866
rect 1945 18808 1950 18864
rect 2006 18808 5262 18864
rect 5318 18808 7654 18864
rect 7710 18808 7715 18864
rect 1945 18806 7715 18808
rect 1945 18803 2011 18806
rect 5257 18803 5323 18806
rect 7649 18803 7715 18806
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 5625 17778 5691 17781
rect 9949 17778 10015 17781
rect 5625 17776 10015 17778
rect 5625 17720 5630 17776
rect 5686 17720 9954 17776
rect 10010 17720 10015 17776
rect 5625 17718 10015 17720
rect 5625 17715 5691 17718
rect 9949 17715 10015 17718
rect 0 17416 480 17536
rect 3610 17440 3930 17441
rect 62 16962 122 17416
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 3969 17234 4035 17237
rect 10777 17234 10843 17237
rect 3969 17232 10843 17234
rect 3969 17176 3974 17232
rect 4030 17176 10782 17232
rect 10838 17176 10843 17232
rect 3969 17174 10843 17176
rect 3969 17171 4035 17174
rect 10777 17171 10843 17174
rect 6821 17098 6887 17101
rect 11513 17098 11579 17101
rect 6821 17096 11579 17098
rect 6821 17040 6826 17096
rect 6882 17040 11518 17096
rect 11574 17040 11579 17096
rect 6821 17038 11579 17040
rect 6821 17035 6887 17038
rect 11513 17035 11579 17038
rect 1301 16962 1367 16965
rect 62 16960 1367 16962
rect 62 16904 1306 16960
rect 1362 16904 1367 16960
rect 62 16902 1367 16904
rect 1301 16899 1367 16902
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 5758 16628 5764 16692
rect 5828 16690 5834 16692
rect 10869 16690 10935 16693
rect 5828 16688 10935 16690
rect 5828 16632 10874 16688
rect 10930 16632 10935 16688
rect 5828 16630 10935 16632
rect 5828 16628 5834 16630
rect 10869 16627 10935 16630
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 4429 14514 4495 14517
rect 8385 14514 8451 14517
rect 11697 14514 11763 14517
rect 4429 14512 11763 14514
rect 4429 14456 4434 14512
rect 4490 14456 8390 14512
rect 8446 14456 11702 14512
rect 11758 14456 11763 14512
rect 4429 14454 11763 14456
rect 4429 14451 4495 14454
rect 8385 14451 8451 14454
rect 11697 14451 11763 14454
rect 13721 14378 13787 14381
rect 8572 14376 13787 14378
rect 8572 14320 13726 14376
rect 13782 14320 13787 14376
rect 8572 14318 13787 14320
rect 8572 14245 8632 14318
rect 13721 14315 13787 14318
rect 5073 14242 5139 14245
rect 8569 14242 8635 14245
rect 5073 14240 8635 14242
rect 5073 14184 5078 14240
rect 5134 14184 8574 14240
rect 8630 14184 8635 14240
rect 5073 14182 8635 14184
rect 5073 14179 5139 14182
rect 8569 14179 8635 14182
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 4613 14106 4679 14109
rect 5758 14106 5764 14108
rect 4613 14104 5764 14106
rect 4613 14048 4618 14104
rect 4674 14048 5764 14104
rect 4613 14046 5764 14048
rect 4613 14043 4679 14046
rect 5758 14044 5764 14046
rect 5828 14044 5834 14108
rect 2497 13834 2563 13837
rect 2773 13834 2839 13837
rect 2497 13832 2839 13834
rect 2497 13776 2502 13832
rect 2558 13776 2778 13832
rect 2834 13776 2839 13832
rect 2497 13774 2839 13776
rect 2497 13771 2563 13774
rect 2773 13771 2839 13774
rect 6913 13834 6979 13837
rect 10041 13834 10107 13837
rect 6913 13832 10107 13834
rect 6913 13776 6918 13832
rect 6974 13776 10046 13832
rect 10102 13776 10107 13832
rect 6913 13774 10107 13776
rect 6913 13771 6979 13774
rect 10041 13771 10107 13774
rect 10225 13834 10291 13837
rect 11053 13834 11119 13837
rect 10225 13832 11119 13834
rect 10225 13776 10230 13832
rect 10286 13776 11058 13832
rect 11114 13776 11119 13832
rect 10225 13774 11119 13776
rect 10225 13771 10291 13774
rect 11053 13771 11119 13774
rect 9489 13698 9555 13701
rect 10041 13698 10107 13701
rect 9362 13696 10107 13698
rect 9362 13640 9494 13696
rect 9550 13640 10046 13696
rect 10102 13640 10107 13696
rect 9362 13638 10107 13640
rect 9489 13635 9555 13638
rect 10041 13635 10107 13638
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 7741 13562 7807 13565
rect 11145 13562 11211 13565
rect 7741 13560 11211 13562
rect 7741 13504 7746 13560
rect 7802 13504 11150 13560
rect 11206 13504 11211 13560
rect 7741 13502 11211 13504
rect 7741 13499 7807 13502
rect 11145 13499 11211 13502
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 6277 12544 6597 12545
rect 0 12384 480 12504
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 62 12202 122 12384
rect 9305 12338 9371 12341
rect 12065 12338 12131 12341
rect 9305 12336 12131 12338
rect 9305 12280 9310 12336
rect 9366 12280 12070 12336
rect 12126 12280 12131 12336
rect 9305 12278 12131 12280
rect 9305 12275 9371 12278
rect 12065 12275 12131 12278
rect 10777 12202 10843 12205
rect 62 12200 10843 12202
rect 62 12144 10782 12200
rect 10838 12144 10843 12200
rect 62 12142 10843 12144
rect 10777 12139 10843 12142
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 1025 11794 1091 11797
rect 10961 11794 11027 11797
rect 1025 11792 11027 11794
rect 1025 11736 1030 11792
rect 1086 11736 10966 11792
rect 11022 11736 11027 11792
rect 1025 11734 11027 11736
rect 1025 11731 1091 11734
rect 10961 11731 11027 11734
rect 4429 11658 4495 11661
rect 7189 11658 7255 11661
rect 4429 11656 7255 11658
rect 4429 11600 4434 11656
rect 4490 11600 7194 11656
rect 7250 11600 7255 11656
rect 4429 11598 7255 11600
rect 4429 11595 4495 11598
rect 7189 11595 7255 11598
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 6126 11188 6132 11252
rect 6196 11250 6202 11252
rect 7373 11250 7439 11253
rect 6196 11248 7439 11250
rect 6196 11192 7378 11248
rect 7434 11192 7439 11248
rect 6196 11190 7439 11192
rect 6196 11188 6202 11190
rect 7373 11187 7439 11190
rect 4981 11114 5047 11117
rect 12157 11114 12223 11117
rect 4981 11112 12223 11114
rect 4981 11056 4986 11112
rect 5042 11056 12162 11112
rect 12218 11056 12223 11112
rect 4981 11054 12223 11056
rect 4981 11051 5047 11054
rect 12157 11051 12223 11054
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 1577 10162 1643 10165
rect 3233 10162 3299 10165
rect 1577 10160 3299 10162
rect 1577 10104 1582 10160
rect 1638 10104 3238 10160
rect 3294 10104 3299 10160
rect 1577 10102 3299 10104
rect 1577 10099 1643 10102
rect 3233 10099 3299 10102
rect 12433 10026 12499 10029
rect 15520 10026 16000 10056
rect 12433 10024 16000 10026
rect 12433 9968 12438 10024
rect 12494 9968 16000 10024
rect 12433 9966 16000 9968
rect 12433 9963 12499 9966
rect 15520 9936 16000 9966
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 1945 9482 2011 9485
rect 5441 9482 5507 9485
rect 11237 9482 11303 9485
rect 1945 9480 4170 9482
rect 1945 9424 1950 9480
rect 2006 9424 4170 9480
rect 1945 9422 4170 9424
rect 1945 9419 2011 9422
rect 4110 9346 4170 9422
rect 5441 9480 11303 9482
rect 5441 9424 5446 9480
rect 5502 9424 11242 9480
rect 11298 9424 11303 9480
rect 5441 9422 11303 9424
rect 5441 9419 5507 9422
rect 11237 9419 11303 9422
rect 5625 9346 5691 9349
rect 4110 9344 5691 9346
rect 4110 9288 5630 9344
rect 5686 9288 5691 9344
rect 4110 9286 5691 9288
rect 5625 9283 5691 9286
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 0 7352 480 7472
rect 62 7034 122 7352
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 1301 7034 1367 7037
rect 62 7032 1367 7034
rect 62 6976 1306 7032
rect 1362 6976 1367 7032
rect 62 6974 1367 6976
rect 1301 6971 1367 6974
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 5349 4178 5415 4181
rect 9857 4178 9923 4181
rect 10225 4178 10291 4181
rect 5349 4176 10291 4178
rect 5349 4120 5354 4176
rect 5410 4120 9862 4176
rect 9918 4120 10230 4176
rect 10286 4120 10291 4176
rect 5349 4118 10291 4120
rect 5349 4115 5415 4118
rect 9857 4115 9923 4118
rect 10225 4115 10291 4118
rect 8385 4042 8451 4045
rect 14181 4042 14247 4045
rect 8385 4040 14247 4042
rect 8385 3984 8390 4040
rect 8446 3984 14186 4040
rect 14242 3984 14247 4040
rect 8385 3982 14247 3984
rect 8385 3979 8451 3982
rect 14181 3979 14247 3982
rect 8017 3906 8083 3909
rect 11421 3906 11487 3909
rect 8017 3904 11487 3906
rect 8017 3848 8022 3904
rect 8078 3848 11426 3904
rect 11482 3848 11487 3904
rect 8017 3846 11487 3848
rect 8017 3843 8083 3846
rect 11421 3843 11487 3846
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 4889 3634 4955 3637
rect 10685 3634 10751 3637
rect 4889 3632 10751 3634
rect 4889 3576 4894 3632
rect 4950 3576 10690 3632
rect 10746 3576 10751 3632
rect 4889 3574 10751 3576
rect 4889 3571 4955 3574
rect 10685 3571 10751 3574
rect 2037 3498 2103 3501
rect 10777 3498 10843 3501
rect 2037 3496 10843 3498
rect 2037 3440 2042 3496
rect 2098 3440 10782 3496
rect 10838 3440 10843 3496
rect 2037 3438 10843 3440
rect 2037 3435 2103 3438
rect 10777 3435 10843 3438
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 3969 3090 4035 3093
rect 12249 3090 12315 3093
rect 3969 3088 12315 3090
rect 3969 3032 3974 3088
rect 4030 3032 12254 3088
rect 12310 3032 12315 3088
rect 3969 3030 12315 3032
rect 3969 3027 4035 3030
rect 12249 3027 12315 3030
rect 9489 2954 9555 2957
rect 62 2952 9555 2954
rect 62 2896 9494 2952
rect 9550 2896 9555 2952
rect 62 2894 9555 2896
rect 62 2576 122 2894
rect 9489 2891 9555 2894
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 0 2456 480 2576
rect 5717 2546 5783 2549
rect 11973 2546 12039 2549
rect 5717 2544 12039 2546
rect 5717 2488 5722 2544
rect 5778 2488 11978 2544
rect 12034 2488 12039 2544
rect 5717 2486 12039 2488
rect 5717 2483 5783 2486
rect 11973 2483 12039 2486
rect 2681 2410 2747 2413
rect 11145 2410 11211 2413
rect 2681 2408 11211 2410
rect 2681 2352 2686 2408
rect 2742 2352 11150 2408
rect 11206 2352 11211 2408
rect 2681 2350 11211 2352
rect 2681 2347 2747 2350
rect 11145 2347 11211 2350
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 6126 1940 6132 2004
rect 6196 2002 6202 2004
rect 12525 2002 12591 2005
rect 6196 2000 12591 2002
rect 6196 1944 12530 2000
rect 12586 1944 12591 2000
rect 6196 1942 12591 1944
rect 6196 1940 6202 1942
rect 12525 1939 12591 1942
rect 5257 1866 5323 1869
rect 13813 1866 13879 1869
rect 5257 1864 13879 1866
rect 5257 1808 5262 1864
rect 5318 1808 13818 1864
rect 13874 1808 13879 1864
rect 5257 1806 13879 1808
rect 5257 1803 5323 1806
rect 13813 1803 13879 1806
rect 3417 1594 3483 1597
rect 9305 1594 9371 1597
rect 3417 1592 9371 1594
rect 3417 1536 3422 1592
rect 3478 1536 9310 1592
rect 9366 1536 9371 1592
rect 3417 1534 9371 1536
rect 3417 1531 3483 1534
rect 9305 1531 9371 1534
rect 1393 98 1459 101
rect 6126 98 6132 100
rect 1393 96 6132 98
rect 1393 40 1398 96
rect 1454 40 6132 96
rect 1393 38 6132 40
rect 1393 35 1459 38
rect 6126 36 6132 38
rect 6196 36 6202 100
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 5764 28460 5828 28524
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 5764 16628 5828 16692
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 5764 14044 5828 14108
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 6132 11188 6196 11252
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
rect 6132 1940 6196 2004
rect 6132 36 6196 100
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 5763 28524 5829 28525
rect 5763 28460 5764 28524
rect 5828 28460 5829 28524
rect 5763 28459 5829 28460
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 5766 16693 5826 28459
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 5763 16692 5829 16693
rect 5763 16628 5764 16692
rect 5828 16628 5829 16692
rect 5763 16627 5829 16628
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 5766 14109 5826 16627
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 5763 14108 5829 14109
rect 5763 14044 5764 14108
rect 5828 14044 5829 14108
rect 5763 14043 5829 14044
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6131 11252 6197 11253
rect 6131 11188 6132 11252
rect 6196 11188 6197 11252
rect 6131 11187 6197 11188
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6134 2005 6194 11187
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
rect 6131 2004 6197 2005
rect 6131 1940 6132 2004
rect 6196 1940 6197 2004
rect 6131 1939 6197 1940
rect 6134 101 6194 1939
rect 6131 100 6197 101
rect 6131 36 6132 100
rect 6196 36 6197 100
rect 6131 35 6197 36
use scs8hd_decap_4  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_9
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_24
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _186_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_130 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_28
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_47
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_43
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_76
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_72
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _183_
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _152_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_buf_2  _188_
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_84
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_88 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 590 592
use scs8hd_buf_2  _185_
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_103 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_100
timestamp 1586364061
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_104
timestamp 1586364061
transform 1 0 10672 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_111 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _184_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_130
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_126
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_128
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_137
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_132 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_144
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_141
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_145
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 1050 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_22
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_26
timestamp 1586364061
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_47
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_51
timestamp 1586364061
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_81
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_85
timestamp 1586364061
transform 1 0 8924 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _180_
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_2  _181_
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_101
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_113
timestamp 1586364061
transform 1 0 11500 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_124
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_143
timestamp 1586364061
transform 1 0 14260 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_10
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_14
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_31
timestamp 1586364061
transform 1 0 3956 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_47
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _187_
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_92
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_100
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_104
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11868 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_111
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_115
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_119
timestamp 1586364061
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_126
timestamp 1586364061
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_130
timestamp 1586364061
transform 1 0 13064 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 4232 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_36
timestamp 1586364061
transform 1 0 4416 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_40
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_52
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_69
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_2  _182_
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_73
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _087_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__C
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_89
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_113
timestamp 1586364061
transform 1 0 11500 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_137
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3220 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_19
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_32
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__D
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_49
timestamp 1586364061
transform 1 0 5612 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_or3_4  _099_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_or3_4  _153_
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_8
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_12
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_19
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_16
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _076_
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_29
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_33
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6072 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_53
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_46
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_50
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_54
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_58
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_61
timestamp 1586364061
transform 1 0 6716 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_57
timestamp 1586364061
transform 1 0 6348 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_or4_4  _135_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_8  _126_
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_74
timestamp 1586364061
transform 1 0 7912 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_78
timestamp 1586364061
transform 1 0 8280 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_81
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_78
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_82
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_or3_4  _066_
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 866 592
use scs8hd_or3_4  _154_
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_85
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_102
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_106
timestamp 1586364061
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_114
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_126
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_6_138
timestamp 1586364061
transform 1 0 13800 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_conb_1  _173_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_35
timestamp 1586364061
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_39
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_2  FILLER_8_43
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_54
timestamp 1586364061
transform 1 0 6072 0 -1 7072
box -38 -48 222 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__C
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_64
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__066__C
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_96
timestamp 1586364061
transform 1 0 9936 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 10120 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_100
timestamp 1586364061
transform 1 0 10304 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_104
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_116
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_128
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 590 592
use scs8hd_conb_1  _172_
timestamp 1586364061
transform 1 0 1564 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_8
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_12
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 2576 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_54
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_58
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use scs8hd_inv_8  _081_
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_105
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_109
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_120
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_143
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_8
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_48
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_52
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 222 592
use scs8hd_or3_4  _082_
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 406 592
use scs8hd_inv_8  _146_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_4  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 406 592
use scs8hd_or3_4  _068_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_buf_1  _101_
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_106
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_113
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_125
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_18
timestamp 1586364061
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_22
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_37
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 314 592
use scs8hd_or2_4  _100_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _084_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_88
timestamp 1586364061
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_109
timestamp 1586364061
transform 1 0 11132 0 1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_117
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_126
timestamp 1586364061
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_130
timestamp 1586364061
transform 1 0 13064 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_20
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_24
timestamp 1586364061
transform 1 0 3312 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 406 592
use scs8hd_or3_4  _110_
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_48
timestamp 1586364061
transform 1 0 5520 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_58
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 590 592
use scs8hd_conb_1  _171_
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_106
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_113
timestamp 1586364061
transform 1 0 11500 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_124
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_12_136
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_9
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 1840 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 2300 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_19
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_23
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 590 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_28
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__C
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_54
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_50
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_or3_4  _118_
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_or2_4  _102_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 682 592
use scs8hd_nor3_4  _144_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__C
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_69
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use scs8hd_conb_1  _170_
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_73
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_72
timestamp 1586364061
transform 1 0 7728 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_76
timestamp 1586364061
transform 1 0 8096 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_4  FILLER_13_88
timestamp 1586364061
transform 1 0 9200 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_90
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_92
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_105
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_109
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_120
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_113
timestamp 1586364061
transform 1 0 11500 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_124
timestamp 1586364061
transform 1 0 12512 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_136
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_13_139
timestamp 1586364061
transform 1 0 13892 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_145
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_20
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_24
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_28
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_41
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _083_
timestamp 1586364061
transform 1 0 5612 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 5060 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_45
timestamp 1586364061
transform 1 0 5244 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_52
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_nor3_4  _143_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_56
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_79
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 314 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_97
timestamp 1586364061
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_116
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 590 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_39
timestamp 1586364061
transform 1 0 4692 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_4  FILLER_16_43
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_47
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__C
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_57
timestamp 1586364061
transform 1 0 6348 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_61
timestamp 1586364061
transform 1 0 6716 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_102
timestamp 1586364061
transform 1 0 10488 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_113
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_137
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_14
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_18
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_33
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_37
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_50
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_54
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_58
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 130 592
use scs8hd_inv_8  _148_
timestamp 1586364061
transform 1 0 8372 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_75
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _163_
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_88
timestamp 1586364061
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_92
timestamp 1586364061
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_105
timestamp 1586364061
transform 1 0 10764 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_109
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_120
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_17
timestamp 1586364061
transform 1 0 2668 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_21
timestamp 1586364061
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_25
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_43
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_47
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_60
timestamp 1586364061
transform 1 0 6624 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_64
timestamp 1586364061
transform 1 0 6992 0 -1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_18_70
timestamp 1586364061
transform 1 0 7544 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 590 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_124
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_136
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_144
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_conb_1  _174_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_13
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 1472 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_17
timestamp 1586364061
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_32
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_43
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_47
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 406 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_68
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_60
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_77
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_81
timestamp 1586364061
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_87
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_85
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_100
timestamp 1586364061
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_104
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_111
timestamp 1586364061
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_115
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_119
timestamp 1586364061
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_119
timestamp 1586364061
transform 1 0 12052 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_126
timestamp 1586364061
transform 1 0 12696 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_130
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_137
timestamp 1586364061
transform 1 0 13708 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_131
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_141
timestamp 1586364061
transform 1 0 14076 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_145
timestamp 1586364061
transform 1 0 14444 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_143
timestamp 1586364061
transform 1 0 14260 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_1  _063_
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_21_9
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_13
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 130 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_16
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_26
timestamp 1586364061
transform 1 0 3496 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 3680 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_30
timestamp 1586364061
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_43
timestamp 1586364061
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_47
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_buf_1  _162_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_65
timestamp 1586364061
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_69
timestamp 1586364061
transform 1 0 7452 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 8280 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_89
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_106
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_21_116
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 590 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_126
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_130
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_137
timestamp 1586364061
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_141
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_145
timestamp 1586364061
transform 1 0 14444 0 1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_or3_4  _167_
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_49
timestamp 1586364061
transform 1 0 5612 0 -1 14688
box -38 -48 774 592
use scs8hd_or3_4  _062_
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_4  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_83
timestamp 1586364061
transform 1 0 8740 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_119
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_130
timestamp 1586364061
transform 1 0 13064 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_142
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 1472 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_24
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_28
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_32
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_36
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_65
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_69
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_90
timestamp 1586364061
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_105
timestamp 1586364061
transform 1 0 10764 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_109
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _175_
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_10
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_8  _147_
timestamp 1586364061
transform 1 0 5704 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 406 592
use scs8hd_or3_4  _157_
timestamp 1586364061
transform 1 0 7268 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_59
timestamp 1586364061
transform 1 0 6532 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  FILLER_24_64
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8280 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_76
timestamp 1586364061
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_88
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_8  _160_
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_8  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_left_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_130
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_142
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_6
timestamp 1586364061
transform 1 0 1656 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_10
timestamp 1586364061
transform 1 0 2024 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_14
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_35
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_49
timestamp 1586364061
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_or3_4  _149_
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_79
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _168_
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_102
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_127
timestamp 1586364061
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use scs8hd_decap_6  FILLER_25_139
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_145
timestamp 1586364061
transform 1 0 14444 0 1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 1050 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_12
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_17
timestamp 1586364061
transform 1 0 2668 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_22
timestamp 1586364061
transform 1 0 3128 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_26
timestamp 1586364061
transform 1 0 3496 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4784 0 1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_31
timestamp 1586364061
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_35
timestamp 1586364061
transform 1 0 4324 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_45
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_55
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 406 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 866 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__C
timestamp 1586364061
transform 1 0 6808 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_58
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_64
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 8280 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_75
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_79
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_83
timestamp 1586364061
transform 1 0 8740 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_76
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_80
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use scs8hd_or3_4  _161_
timestamp 1586364061
transform 1 0 8832 0 1 16864
box -38 -48 866 592
use scs8hd_or3_4  _164_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_86
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_91
timestamp 1586364061
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_93
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 11224 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_104
timestamp 1586364061
transform 1 0 10672 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_108
timestamp 1586364061
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_113
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_26_124
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_112
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_116
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 590 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_136
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_126
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_130
timestamp 1586364061
transform 1 0 13064 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_137
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_144
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_141
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_145
timestamp 1586364061
transform 1 0 14444 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_18
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_22
timestamp 1586364061
transform 1 0 3128 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_26
timestamp 1586364061
transform 1 0 3496 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_43
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_47
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_60
timestamp 1586364061
transform 1 0 6624 0 -1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_77
timestamp 1586364061
transform 1 0 8188 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_81
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_8  FILLER_28_119
timestamp 1586364061
transform 1 0 12052 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_130
timestamp 1586364061
transform 1 0 13064 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_142
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 406 592
use scs8hd_buf_1  _071_
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 2300 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_11
timestamp 1586364061
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_30
timestamp 1586364061
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_47
timestamp 1586364061
transform 1 0 5428 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_69
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_73
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_88
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_92
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_105
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_109
timestamp 1586364061
transform 1 0 11132 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_113
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_117
timestamp 1586364061
transform 1 0 11868 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_126
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_130
timestamp 1586364061
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_137
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_141
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_145
timestamp 1586364061
transform 1 0 14444 0 1 17952
box -38 -48 130 592
use scs8hd_buf_1  _073_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_10
timestamp 1586364061
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_6  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 6164 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_45
timestamp 1586364061
transform 1 0 5244 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_53
timestamp 1586364061
transform 1 0 5980 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_30_72
timestamp 1586364061
transform 1 0 7728 0 -1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_119
timestamp 1586364061
transform 1 0 12052 0 -1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_130
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_30_142
timestamp 1586364061
transform 1 0 14168 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 866 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 1656 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_8
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_21
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_25
timestamp 1586364061
transform 1 0 3404 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_38
timestamp 1586364061
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use scs8hd_buf_1  _151_
timestamp 1586364061
transform 1 0 5704 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_42
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_46
timestamp 1586364061
transform 1 0 5336 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7176 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_69
timestamp 1586364061
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_73
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_88
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_92
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_105
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_109
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_113
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_117
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_126
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_130
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_134
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 1840 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_10
timestamp 1586364061
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_36
timestamp 1586364061
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6072 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_32_46
timestamp 1586364061
transform 1 0 5336 0 -1 20128
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_65
timestamp 1586364061
transform 1 0 7084 0 -1 20128
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_32_70
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 314 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_106
timestamp 1586364061
transform 1 0 10856 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_32_119
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 774 592
use scs8hd_buf_1  _119_
timestamp 1586364061
transform 1 0 12788 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_130
timestamp 1586364061
transform 1 0 13064 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_142
timestamp 1586364061
transform 1 0 14168 0 -1 20128
box -38 -48 406 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 2024 0 -1 21216
box -38 -48 1050 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 1564 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_17
timestamp 1586364061
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_21
timestamp 1586364061
transform 1 0 3036 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_25
timestamp 1586364061
transform 1 0 3404 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_21
timestamp 1586364061
transform 1 0 3036 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_25
timestamp 1586364061
transform 1 0 3404 0 -1 21216
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3680 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_37
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_41
timestamp 1586364061
transform 1 0 4876 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_30
timestamp 1586364061
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_47
timestamp 1586364061
transform 1 0 5428 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_43
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_47
timestamp 1586364061
transform 1 0 5428 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 5244 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use scs8hd_buf_1  _150_
timestamp 1586364061
transform 1 0 5704 0 1 20128
box -38 -48 314 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 5796 0 -1 21216
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_60
timestamp 1586364061
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_57
timestamp 1586364061
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_64
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_68
timestamp 1586364061
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 7176 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7084 0 1 20128
box -38 -48 314 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 8096 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7544 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_72
timestamp 1586364061
transform 1 0 7728 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_77
timestamp 1586364061
transform 1 0 8188 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_81
timestamp 1586364061
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_87
timestamp 1586364061
transform 1 0 9108 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_91
timestamp 1586364061
transform 1 0 9476 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_85
timestamp 1586364061
transform 1 0 8924 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_91
timestamp 1586364061
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 11224 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_104
timestamp 1586364061
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_108
timestamp 1586364061
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_102
timestamp 1586364061
transform 1 0 10488 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_106
timestamp 1586364061
transform 1 0 10856 0 -1 21216
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_112
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_120
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_113
timestamp 1586364061
transform 1 0 11500 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_125
timestamp 1586364061
transform 1 0 12604 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_137
timestamp 1586364061
transform 1 0 13708 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_145
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 130 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 866 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_12
timestamp 1586364061
transform 1 0 2208 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 2944 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_16
timestamp 1586364061
transform 1 0 2576 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 4140 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_31
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4968 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_53
timestamp 1586364061
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_57
timestamp 1586364061
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_71
timestamp 1586364061
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_conb_1  _178_
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 10672 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_99
timestamp 1586364061
transform 1 0 10212 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_103
timestamp 1586364061
transform 1 0 10580 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_35_143
timestamp 1586364061
transform 1 0 14260 0 1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 1840 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_6
timestamp 1586364061
transform 1 0 1656 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_10
timestamp 1586364061
transform 1 0 2024 0 -1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_36_23
timestamp 1586364061
transform 1 0 3220 0 -1 22304
box -38 -48 774 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 4140 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_36
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_55
timestamp 1586364061
transform 1 0 6164 0 -1 22304
box -38 -48 774 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 6900 0 -1 22304
box -38 -48 866 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7912 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_72
timestamp 1586364061
transform 1 0 7728 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_76
timestamp 1586364061
transform 1 0 8096 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_83
timestamp 1586364061
transform 1 0 8740 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 8924 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_87
timestamp 1586364061
transform 1 0 9108 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_91
timestamp 1586364061
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_96
timestamp 1586364061
transform 1 0 9936 0 -1 22304
box -38 -48 222 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 10672 0 -1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 10120 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_100
timestamp 1586364061
transform 1 0 10304 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_36_107
timestamp 1586364061
transform 1 0 10948 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_119
timestamp 1586364061
transform 1 0 12052 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_131
timestamp 1586364061
transform 1 0 13156 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_36_143
timestamp 1586364061
transform 1 0 14260 0 -1 22304
box -38 -48 314 592
use scs8hd_conb_1  _176_
timestamp 1586364061
transform 1 0 2208 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_7
timestamp 1586364061
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_11
timestamp 1586364061
transform 1 0 2116 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 2944 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_19
timestamp 1586364061
transform 1 0 2852 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_22
timestamp 1586364061
transform 1 0 3128 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3956 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_40
timestamp 1586364061
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use scs8hd_conb_1  _177_
timestamp 1586364061
transform 1 0 5704 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 5428 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_37_44
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 314 592
use scs8hd_fill_1  FILLER_37_49
timestamp 1586364061
transform 1 0 5612 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 8372 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_88
timestamp 1586364061
transform 1 0 9200 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_105
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_109
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_112
timestamp 1586364061
transform 1 0 11408 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_120
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use scs8hd_decap_3  FILLER_37_143
timestamp 1586364061
transform 1 0 14260 0 1 22304
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 2024 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_6
timestamp 1586364061
transform 1 0 1656 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_12
timestamp 1586364061
transform 1 0 2208 0 -1 23392
box -38 -48 222 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 2944 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 2392 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_16
timestamp 1586364061
transform 1 0 2576 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_23
timestamp 1586364061
transform 1 0 3220 0 -1 23392
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4232 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_29
timestamp 1586364061
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_37
timestamp 1586364061
transform 1 0 4508 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_41
timestamp 1586364061
transform 1 0 4876 0 -1 23392
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 23392
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_46
timestamp 1586364061
transform 1 0 5336 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 7452 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_58
timestamp 1586364061
transform 1 0 6440 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_38_64
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7728 0 -1 23392
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_38_71
timestamp 1586364061
transform 1 0 7636 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_83
timestamp 1586364061
transform 1 0 8740 0 -1 23392
box -38 -48 774 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_91
timestamp 1586364061
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_106
timestamp 1586364061
transform 1 0 10856 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_113
timestamp 1586364061
transform 1 0 11500 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_125
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_38_137
timestamp 1586364061
transform 1 0 13708 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_4  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_9
timestamp 1586364061
transform 1 0 1932 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2024 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 866 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 2208 0 -1 24480
box -38 -48 866 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_19
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_23
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_21
timestamp 1586364061
transform 1 0 3036 0 -1 24480
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_36
timestamp 1586364061
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_40
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_41
timestamp 1586364061
transform 1 0 4876 0 -1 24480
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_53
timestamp 1586364061
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_51
timestamp 1586364061
transform 1 0 5796 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_61
timestamp 1586364061
transform 1 0 6716 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_65
timestamp 1586364061
transform 1 0 7084 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_68
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 7176 0 -1 24480
box -38 -48 222 592
use scs8hd_nor2_4  _137_
timestamp 1586364061
transform 1 0 7452 0 -1 24480
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7728 0 1 23392
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_83
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_78
timestamp 1586364061
transform 1 0 8280 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_82
timestamp 1586364061
transform 1 0 8648 0 -1 24480
box -38 -48 774 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 9476 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 9292 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_87
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_90
timestamp 1586364061
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 11224 0 -1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_100
timestamp 1586364061
transform 1 0 10304 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_104
timestamp 1586364061
transform 1 0 10672 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_102
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 11868 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_111
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_115
timestamp 1586364061
transform 1 0 11684 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_119
timestamp 1586364061
transform 1 0 12052 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_114
timestamp 1586364061
transform 1 0 11592 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_126
timestamp 1586364061
transform 1 0 12696 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_138
timestamp 1586364061
transform 1 0 13800 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_39_143
timestamp 1586364061
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 2208 0 1 24480
box -38 -48 866 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2024 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 1656 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_8
timestamp 1586364061
transform 1 0 1840 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_21
timestamp 1586364061
transform 1 0 3036 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_25
timestamp 1586364061
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 3772 0 1 24480
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_41_40
timestamp 1586364061
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5520 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_44
timestamp 1586364061
transform 1 0 5152 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_55
timestamp 1586364061
transform 1 0 6164 0 1 24480
box -38 -48 406 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 8372 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 8188 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_71
timestamp 1586364061
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_75
timestamp 1586364061
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_41_88
timestamp 1586364061
transform 1 0 9200 0 1 24480
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 10948 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_105
timestamp 1586364061
transform 1 0 10764 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_109
timestamp 1586364061
transform 1 0 11132 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_121
timestamp 1586364061
transform 1 0 12236 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 25568
box -38 -48 1050 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_8  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_11
timestamp 1586364061
transform 1 0 2116 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_23
timestamp 1586364061
transform 1 0 3220 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_42_41
timestamp 1586364061
transform 1 0 4876 0 -1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_45
timestamp 1586364061
transform 1 0 5244 0 -1 25568
box -38 -48 406 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 7176 0 -1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_58
timestamp 1586364061
transform 1 0 6440 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_64
timestamp 1586364061
transform 1 0 6992 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 8372 0 -1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 406 592
use scs8hd_fill_2  FILLER_42_81
timestamp 1586364061
transform 1 0 8556 0 -1 25568
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_6  FILLER_42_85
timestamp 1586364061
transform 1 0 8924 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_42_91
timestamp 1586364061
transform 1 0 9476 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_3  FILLER_42_93
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 314 592
use scs8hd_buf_2  _189_
timestamp 1586364061
transform 1 0 10120 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_102
timestamp 1586364061
transform 1 0 10488 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_114
timestamp 1586364061
transform 1 0 11592 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_126
timestamp 1586364061
transform 1 0 12696 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_42_138
timestamp 1586364061
transform 1 0 13800 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1748 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_86
timestamp 1586364061
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_3
timestamp 1586364061
transform 1 0 1380 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_10
timestamp 1586364061
transform 1 0 2024 0 1 25568
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2760 0 1 25568
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_14
timestamp 1586364061
transform 1 0 2392 0 1 25568
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4508 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_29
timestamp 1586364061
transform 1 0 3772 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_34
timestamp 1586364061
transform 1 0 4232 0 1 25568
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5520 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_46
timestamp 1586364061
transform 1 0 5336 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_50
timestamp 1586364061
transform 1 0 5704 0 1 25568
box -38 -48 222 592
use scs8hd_decap_4  FILLER_43_54
timestamp 1586364061
transform 1 0 6072 0 1 25568
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_43_58
timestamp 1586364061
transform 1 0 6440 0 1 25568
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 25568
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 25568
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8280 0 1 25568
box -38 -48 222 592
use scs8hd_fill_2  FILLER_43_71
timestamp 1586364061
transform 1 0 7636 0 1 25568
box -38 -48 222 592
use scs8hd_decap_3  FILLER_43_75
timestamp 1586364061
transform 1 0 8004 0 1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_43_89
timestamp 1586364061
transform 1 0 9292 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_43_101
timestamp 1586364061
transform 1 0 10396 0 1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_43_113
timestamp 1586364061
transform 1 0 11500 0 1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_43_121
timestamp 1586364061
transform 1 0 12236 0 1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_43_123
timestamp 1586364061
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_43_135
timestamp 1586364061
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use scs8hd_decap_3  PHY_87
timestamp 1586364061
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  FILLER_43_143
timestamp 1586364061
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use scs8hd_decap_3  PHY_88
timestamp 1586364061
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_44_3
timestamp 1586364061
transform 1 0 1380 0 -1 26656
box -38 -48 774 592
use scs8hd_fill_1  FILLER_44_11
timestamp 1586364061
transform 1 0 2116 0 -1 26656
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_23
timestamp 1586364061
transform 1 0 3220 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_27
timestamp 1586364061
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 26656
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_35
timestamp 1586364061
transform 1 0 4324 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_4  FILLER_44_39
timestamp 1586364061
transform 1 0 4692 0 -1 26656
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5336 0 -1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5060 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_44_45
timestamp 1586364061
transform 1 0 5244 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7360 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6992 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6624 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_3  FILLER_44_57
timestamp 1586364061
transform 1 0 6348 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_2  FILLER_44_62
timestamp 1586364061
transform 1 0 6808 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_44_66
timestamp 1586364061
transform 1 0 7176 0 -1 26656
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7544 0 -1 26656
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_44_81
timestamp 1586364061
transform 1 0 8556 0 -1 26656
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 -1 26656
box -38 -48 222 592
use scs8hd_fill_1  FILLER_44_91
timestamp 1586364061
transform 1 0 9476 0 -1 26656
box -38 -48 130 592
use scs8hd_fill_2  FILLER_44_93
timestamp 1586364061
transform 1 0 9660 0 -1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_44_97
timestamp 1586364061
transform 1 0 10028 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_109
timestamp 1586364061
transform 1 0 11132 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_121
timestamp 1586364061
transform 1 0 12236 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_44_133
timestamp 1586364061
transform 1 0 13340 0 -1 26656
box -38 -48 1142 592
use scs8hd_decap_3  PHY_89
timestamp 1586364061
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use scs8hd_fill_1  FILLER_44_145
timestamp 1586364061
transform 1 0 14444 0 -1 26656
box -38 -48 130 592
use scs8hd_decap_3  PHY_90
timestamp 1586364061
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use scs8hd_decap_8  FILLER_45_3
timestamp 1586364061
transform 1 0 1380 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  FILLER_45_11
timestamp 1586364061
transform 1 0 2116 0 1 26656
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 26656
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3404 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_17
timestamp 1586364061
transform 1 0 2668 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_21
timestamp 1586364061
transform 1 0 3036 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_34
timestamp 1586364061
transform 1 0 4232 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_38
timestamp 1586364061
transform 1 0 4600 0 1 26656
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_53
timestamp 1586364061
transform 1 0 5980 0 1 26656
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7360 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6992 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_57
timestamp 1586364061
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_62
timestamp 1586364061
transform 1 0 6808 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_66
timestamp 1586364061
transform 1 0 7176 0 1 26656
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7544 0 1 26656
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_81
timestamp 1586364061
transform 1 0 8556 0 1 26656
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9292 0 1 26656
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9108 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_85
timestamp 1586364061
transform 1 0 8924 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 26656
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 26656
box -38 -48 222 592
use scs8hd_fill_2  FILLER_45_98
timestamp 1586364061
transform 1 0 10120 0 1 26656
box -38 -48 222 592
use scs8hd_decap_8  FILLER_45_102
timestamp 1586364061
transform 1 0 10488 0 1 26656
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use scs8hd_decap_8  FILLER_45_112
timestamp 1586364061
transform 1 0 11408 0 1 26656
box -38 -48 774 592
use scs8hd_fill_2  FILLER_45_120
timestamp 1586364061
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use scs8hd_decap_12  FILLER_45_123
timestamp 1586364061
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_45_135
timestamp 1586364061
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use scs8hd_decap_3  PHY_91
timestamp 1586364061
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  FILLER_45_143
timestamp 1586364061
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use scs8hd_decap_3  PHY_92
timestamp 1586364061
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_94
timestamp 1586364061
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use scs8hd_decap_12  FILLER_46_3
timestamp 1586364061
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_47_3
timestamp 1586364061
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_47_15
timestamp 1586364061
transform 1 0 2484 0 1 27744
box -38 -48 590 592
use scs8hd_fill_1  FILLER_46_19
timestamp 1586364061
transform 1 0 2852 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_15
timestamp 1586364061
transform 1 0 2484 0 -1 27744
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_25
timestamp 1586364061
transform 1 0 3404 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_21
timestamp 1586364061
transform 1 0 3036 0 1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_27
timestamp 1586364061
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_46_23
timestamp 1586364061
transform 1 0 3220 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3588 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3128 0 1 27744
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 27744
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 1 27744
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_6  FILLER_46_35
timestamp 1586364061
transform 1 0 4324 0 -1 27744
box -38 -48 590 592
use scs8hd_decap_4  FILLER_47_29
timestamp 1586364061
transform 1 0 3772 0 1 27744
box -38 -48 406 592
use scs8hd_fill_2  FILLER_47_36
timestamp 1586364061
transform 1 0 4416 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_40
timestamp 1586364061
transform 1 0 4784 0 1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5060 0 -1 27744
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_46_54
timestamp 1586364061
transform 1 0 6072 0 -1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_53
timestamp 1586364061
transform 1 0 5980 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_47_62
timestamp 1586364061
transform 1 0 6808 0 1 27744
box -38 -48 130 592
use scs8hd_fill_2  FILLER_47_57
timestamp 1586364061
transform 1 0 6348 0 1 27744
box -38 -48 222 592
use scs8hd_fill_1  FILLER_46_62
timestamp 1586364061
transform 1 0 6808 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_4  FILLER_46_58
timestamp 1586364061
transform 1 0 6440 0 -1 27744
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use scs8hd_decap_3  FILLER_46_65
timestamp 1586364061
transform 1 0 7084 0 -1 27744
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6900 0 -1 27744
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6900 0 1 27744
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7360 0 -1 27744
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8648 0 1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8464 0 1 27744
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8648 0 -1 27744
box -38 -48 222 592
use scs8hd_decap_3  FILLER_46_79
timestamp 1586364061
transform 1 0 8372 0 -1 27744
box -38 -48 314 592
use scs8hd_fill_2  FILLER_47_74
timestamp 1586364061
transform 1 0 7912 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_78
timestamp 1586364061
transform 1 0 8280 0 1 27744
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 27744
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_84
timestamp 1586364061
transform 1 0 8832 0 -1 27744
box -38 -48 774 592
use scs8hd_fill_2  FILLER_47_91
timestamp 1586364061
transform 1 0 9476 0 1 27744
box -38 -48 222 592
use scs8hd_fill_2  FILLER_47_95
timestamp 1586364061
transform 1 0 9844 0 1 27744
box -38 -48 222 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 -1 27744
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 27744
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 27744
box -38 -48 222 592
use scs8hd_decap_8  FILLER_46_102
timestamp 1586364061
transform 1 0 10488 0 -1 27744
box -38 -48 774 592
use scs8hd_decap_12  FILLER_47_108
timestamp 1586364061
transform 1 0 11040 0 1 27744
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use scs8hd_decap_12  FILLER_46_113
timestamp 1586364061
transform 1 0 11500 0 -1 27744
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_47_120
timestamp 1586364061
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use scs8hd_decap_12  FILLER_47_123
timestamp 1586364061
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_46_125
timestamp 1586364061
transform 1 0 12604 0 -1 27744
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_46_137
timestamp 1586364061
transform 1 0 13708 0 -1 27744
box -38 -48 774 592
use scs8hd_decap_8  FILLER_47_135
timestamp 1586364061
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use scs8hd_decap_3  PHY_93
timestamp 1586364061
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_95
timestamp 1586364061
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use scs8hd_fill_1  FILLER_46_145
timestamp 1586364061
transform 1 0 14444 0 -1 27744
box -38 -48 130 592
use scs8hd_decap_3  FILLER_47_143
timestamp 1586364061
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use scs8hd_decap_3  PHY_96
timestamp 1586364061
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_48_3
timestamp 1586364061
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_15
timestamp 1586364061
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_48_27
timestamp 1586364061
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_48_32
timestamp 1586364061
transform 1 0 4048 0 -1 28832
box -38 -48 774 592
use scs8hd_fill_1  FILLER_48_40
timestamp 1586364061
transform 1 0 4784 0 -1 28832
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5704 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_44
timestamp 1586364061
transform 1 0 5152 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_48
timestamp 1586364061
transform 1 0 5520 0 -1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6900 0 -1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_61
timestamp 1586364061
transform 1 0 6716 0 -1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_48_65
timestamp 1586364061
transform 1 0 7084 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_48_78
timestamp 1586364061
transform 1 0 8280 0 -1 28832
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 28832
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use scs8hd_fill_2  FILLER_48_90
timestamp 1586364061
transform 1 0 9384 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_3  FILLER_48_96
timestamp 1586364061
transform 1 0 9936 0 -1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 -1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_48_101
timestamp 1586364061
transform 1 0 10396 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_113
timestamp 1586364061
transform 1 0 11500 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_48_125
timestamp 1586364061
transform 1 0 12604 0 -1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_48_137
timestamp 1586364061
transform 1 0 13708 0 -1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_97
timestamp 1586364061
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use scs8hd_fill_1  FILLER_48_145
timestamp 1586364061
transform 1 0 14444 0 -1 28832
box -38 -48 130 592
use scs8hd_decap_3  PHY_98
timestamp 1586364061
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use scs8hd_decap_12  FILLER_49_3
timestamp 1586364061
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_15
timestamp 1586364061
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_27
timestamp 1586364061
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 28832
box -38 -48 314 592
use scs8hd_inv_1  mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 28832
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_42
timestamp 1586364061
transform 1 0 4968 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_46
timestamp 1586364061
transform 1 0 5336 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_53
timestamp 1586364061
transform 1 0 5980 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 28832
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_57
timestamp 1586364061
transform 1 0 6348 0 1 28832
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 28832
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 28832
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_71
timestamp 1586364061
transform 1 0 7636 0 1 28832
box -38 -48 222 592
use scs8hd_fill_2  FILLER_49_75
timestamp 1586364061
transform 1 0 8004 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_88
timestamp 1586364061
transform 1 0 9200 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_49_100
timestamp 1586364061
transform 1 0 10304 0 1 28832
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use scs8hd_decap_8  FILLER_49_112
timestamp 1586364061
transform 1 0 11408 0 1 28832
box -38 -48 774 592
use scs8hd_fill_2  FILLER_49_120
timestamp 1586364061
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use scs8hd_decap_12  FILLER_49_123
timestamp 1586364061
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_49_135
timestamp 1586364061
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use scs8hd_decap_3  PHY_99
timestamp 1586364061
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  FILLER_49_143
timestamp 1586364061
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use scs8hd_decap_3  PHY_100
timestamp 1586364061
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_3
timestamp 1586364061
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_15
timestamp 1586364061
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_50_27
timestamp 1586364061
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_50_32
timestamp 1586364061
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 29920
box -38 -48 866 592
use scs8hd_decap_8  FILLER_50_44
timestamp 1586364061
transform 1 0 5152 0 -1 29920
box -38 -48 774 592
use scs8hd_inv_1  mux_right_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7452 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_8  FILLER_50_61
timestamp 1586364061
transform 1 0 6716 0 -1 29920
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 -1 29920
box -38 -48 222 592
use scs8hd_decap_6  FILLER_50_72
timestamp 1586364061
transform 1 0 7728 0 -1 29920
box -38 -48 590 592
use scs8hd_fill_1  FILLER_50_78
timestamp 1586364061
transform 1 0 8280 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_8  FILLER_50_81
timestamp 1586364061
transform 1 0 8556 0 -1 29920
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use scs8hd_decap_3  FILLER_50_89
timestamp 1586364061
transform 1 0 9292 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_12  FILLER_50_93
timestamp 1586364061
transform 1 0 9660 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_105
timestamp 1586364061
transform 1 0 10764 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_117
timestamp 1586364061
transform 1 0 11868 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_50_129
timestamp 1586364061
transform 1 0 12972 0 -1 29920
box -38 -48 1142 592
use scs8hd_decap_3  PHY_101
timestamp 1586364061
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use scs8hd_decap_4  FILLER_50_141
timestamp 1586364061
transform 1 0 14076 0 -1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_50_145
timestamp 1586364061
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use scs8hd_inv_1  mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_102
timestamp 1586364061
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 29920
box -38 -48 222 592
use scs8hd_fill_2  FILLER_51_6
timestamp 1586364061
transform 1 0 1656 0 1 29920
box -38 -48 222 592
use scs8hd_decap_12  FILLER_51_10
timestamp 1586364061
transform 1 0 2024 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_22
timestamp 1586364061
transform 1 0 3128 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_34
timestamp 1586364061
transform 1 0 4232 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_46
timestamp 1586364061
transform 1 0 5336 0 1 29920
box -38 -48 1142 592
use scs8hd_conb_1  _179_
timestamp 1586364061
transform 1 0 7268 0 1 29920
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use scs8hd_decap_3  FILLER_51_58
timestamp 1586364061
transform 1 0 6440 0 1 29920
box -38 -48 314 592
use scs8hd_decap_4  FILLER_51_62
timestamp 1586364061
transform 1 0 6808 0 1 29920
box -38 -48 406 592
use scs8hd_fill_1  FILLER_51_66
timestamp 1586364061
transform 1 0 7176 0 1 29920
box -38 -48 130 592
use scs8hd_decap_12  FILLER_51_70
timestamp 1586364061
transform 1 0 7544 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_82
timestamp 1586364061
transform 1 0 8648 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_94
timestamp 1586364061
transform 1 0 9752 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_51_106
timestamp 1586364061
transform 1 0 10856 0 1 29920
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use scs8hd_decap_4  FILLER_51_118
timestamp 1586364061
transform 1 0 11960 0 1 29920
box -38 -48 406 592
use scs8hd_decap_12  FILLER_51_123
timestamp 1586364061
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_51_135
timestamp 1586364061
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use scs8hd_decap_3  PHY_103
timestamp 1586364061
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  FILLER_51_143
timestamp 1586364061
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use scs8hd_decap_3  PHY_104
timestamp 1586364061
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_106
timestamp 1586364061
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use scs8hd_decap_12  FILLER_52_3
timestamp 1586364061
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_3
timestamp 1586364061
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_15
timestamp 1586364061
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_52_27
timestamp 1586364061
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use scs8hd_decap_12  FILLER_53_15
timestamp 1586364061
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_27
timestamp 1586364061
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_32
timestamp 1586364061
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_39
timestamp 1586364061
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_44
timestamp 1586364061
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_51
timestamp 1586364061
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_56
timestamp 1586364061
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_68
timestamp 1586364061
transform 1 0 7360 0 -1 31008
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_53_59
timestamp 1586364061
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use scs8hd_decap_12  FILLER_53_62
timestamp 1586364061
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_80
timestamp 1586364061
transform 1 0 8464 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_74
timestamp 1586364061
transform 1 0 7912 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_93
timestamp 1586364061
transform 1 0 9660 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_86
timestamp 1586364061
transform 1 0 9016 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_105
timestamp 1586364061
transform 1 0 10764 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_98
timestamp 1586364061
transform 1 0 10120 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_110
timestamp 1586364061
transform 1 0 11224 0 1 31008
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use scs8hd_decap_12  FILLER_52_117
timestamp 1586364061
transform 1 0 11868 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_53_123
timestamp 1586364061
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_52_129
timestamp 1586364061
transform 1 0 12972 0 -1 31008
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_53_135
timestamp 1586364061
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use scs8hd_decap_3  PHY_105
timestamp 1586364061
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_107
timestamp 1586364061
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use scs8hd_decap_4  FILLER_52_141
timestamp 1586364061
transform 1 0 14076 0 -1 31008
box -38 -48 406 592
use scs8hd_fill_1  FILLER_52_145
timestamp 1586364061
transform 1 0 14444 0 -1 31008
box -38 -48 130 592
use scs8hd_decap_3  FILLER_53_143
timestamp 1586364061
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use scs8hd_decap_3  PHY_108
timestamp 1586364061
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_54_3
timestamp 1586364061
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_15
timestamp 1586364061
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_54_27
timestamp 1586364061
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_32
timestamp 1586364061
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_44
timestamp 1586364061
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_56
timestamp 1586364061
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_68
timestamp 1586364061
transform 1 0 7360 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_80
timestamp 1586364061
transform 1 0 8464 0 -1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_54_93
timestamp 1586364061
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_105
timestamp 1586364061
transform 1 0 10764 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_117
timestamp 1586364061
transform 1 0 11868 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_54_129
timestamp 1586364061
transform 1 0 12972 0 -1 32096
box -38 -48 1142 592
use scs8hd_decap_3  PHY_109
timestamp 1586364061
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use scs8hd_decap_4  FILLER_54_141
timestamp 1586364061
transform 1 0 14076 0 -1 32096
box -38 -48 406 592
use scs8hd_fill_1  FILLER_54_145
timestamp 1586364061
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use scs8hd_decap_3  PHY_110
timestamp 1586364061
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use scs8hd_decap_12  FILLER_55_3
timestamp 1586364061
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_15
timestamp 1586364061
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_27
timestamp 1586364061
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_39
timestamp 1586364061
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_51
timestamp 1586364061
transform 1 0 5796 0 1 32096
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use scs8hd_fill_2  FILLER_55_59
timestamp 1586364061
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use scs8hd_decap_12  FILLER_55_62
timestamp 1586364061
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_74
timestamp 1586364061
transform 1 0 7912 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_86
timestamp 1586364061
transform 1 0 9016 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_98
timestamp 1586364061
transform 1 0 10120 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_55_110
timestamp 1586364061
transform 1 0 11224 0 1 32096
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use scs8hd_decap_12  FILLER_55_123
timestamp 1586364061
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_55_135
timestamp 1586364061
transform 1 0 13524 0 1 32096
box -38 -48 774 592
use scs8hd_decap_3  PHY_111
timestamp 1586364061
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  FILLER_55_143
timestamp 1586364061
transform 1 0 14260 0 1 32096
box -38 -48 314 592
use scs8hd_decap_3  PHY_112
timestamp 1586364061
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_56_3
timestamp 1586364061
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_15
timestamp 1586364061
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_56_27
timestamp 1586364061
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_32
timestamp 1586364061
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_44
timestamp 1586364061
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_56
timestamp 1586364061
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_68
timestamp 1586364061
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_80
timestamp 1586364061
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_12  FILLER_56_93
timestamp 1586364061
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_105
timestamp 1586364061
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_117
timestamp 1586364061
transform 1 0 11868 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_56_129
timestamp 1586364061
transform 1 0 12972 0 -1 33184
box -38 -48 1142 592
use scs8hd_decap_3  PHY_113
timestamp 1586364061
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use scs8hd_decap_4  FILLER_56_141
timestamp 1586364061
transform 1 0 14076 0 -1 33184
box -38 -48 406 592
use scs8hd_fill_1  FILLER_56_145
timestamp 1586364061
transform 1 0 14444 0 -1 33184
box -38 -48 130 592
use scs8hd_decap_3  PHY_114
timestamp 1586364061
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use scs8hd_decap_12  FILLER_57_3
timestamp 1586364061
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_15
timestamp 1586364061
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_27
timestamp 1586364061
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_39
timestamp 1586364061
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_51
timestamp 1586364061
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use scs8hd_fill_2  FILLER_57_59
timestamp 1586364061
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_62
timestamp 1586364061
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 8096 0 1 33184
box -38 -48 222 592
use scs8hd_fill_2  FILLER_57_74
timestamp 1586364061
transform 1 0 7912 0 1 33184
box -38 -48 222 592
use scs8hd_decap_12  FILLER_57_78
timestamp 1586364061
transform 1 0 8280 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_90
timestamp 1586364061
transform 1 0 9384 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_57_102
timestamp 1586364061
transform 1 0 10488 0 1 33184
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use scs8hd_decap_8  FILLER_57_114
timestamp 1586364061
transform 1 0 11592 0 1 33184
box -38 -48 774 592
use scs8hd_decap_12  FILLER_57_123
timestamp 1586364061
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_57_135
timestamp 1586364061
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use scs8hd_decap_3  PHY_115
timestamp 1586364061
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  FILLER_57_143
timestamp 1586364061
transform 1 0 14260 0 1 33184
box -38 -48 314 592
use scs8hd_decap_3  PHY_116
timestamp 1586364061
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_12  FILLER_58_3
timestamp 1586364061
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_15
timestamp 1586364061
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_58_27
timestamp 1586364061
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_32
timestamp 1586364061
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_44
timestamp 1586364061
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_56
timestamp 1586364061
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_58_68
timestamp 1586364061
transform 1 0 7360 0 -1 34272
box -38 -48 774 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 8096 0 -1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_58_80
timestamp 1586364061
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_12  FILLER_58_93
timestamp 1586364061
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_105
timestamp 1586364061
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_117
timestamp 1586364061
transform 1 0 11868 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_58_129
timestamp 1586364061
transform 1 0 12972 0 -1 34272
box -38 -48 1142 592
use scs8hd_decap_3  PHY_117
timestamp 1586364061
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use scs8hd_decap_4  FILLER_58_141
timestamp 1586364061
transform 1 0 14076 0 -1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_58_145
timestamp 1586364061
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use scs8hd_decap_3  PHY_118
timestamp 1586364061
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_120
timestamp 1586364061
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_59_3
timestamp 1586364061
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_3
timestamp 1586364061
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_59_15
timestamp 1586364061
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_59_27
timestamp 1586364061
transform 1 0 3588 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_15
timestamp 1586364061
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_60_27
timestamp 1586364061
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 4508 0 1 34272
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_35
timestamp 1586364061
transform 1 0 4324 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_41
timestamp 1586364061
transform 1 0 4876 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_60_32
timestamp 1586364061
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 5060 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_45
timestamp 1586364061
transform 1 0 5244 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_44
timestamp 1586364061
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _191_
timestamp 1586364061
transform 1 0 6808 0 1 34272
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_57
timestamp 1586364061
transform 1 0 6348 0 1 34272
box -38 -48 222 592
use scs8hd_decap_4  FILLER_59_66
timestamp 1586364061
transform 1 0 7176 0 1 34272
box -38 -48 406 592
use scs8hd_decap_12  FILLER_60_56
timestamp 1586364061
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_60_68
timestamp 1586364061
transform 1 0 7360 0 -1 35360
box -38 -48 314 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 8280 0 1 34272
box -38 -48 406 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 7636 0 -1 35360
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 7636 0 1 34272
box -38 -48 222 592
use scs8hd_fill_1  FILLER_59_70
timestamp 1586364061
transform 1 0 7544 0 1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_59_73
timestamp 1586364061
transform 1 0 7820 0 1 34272
box -38 -48 406 592
use scs8hd_fill_1  FILLER_59_77
timestamp 1586364061
transform 1 0 8188 0 1 34272
box -38 -48 130 592
use scs8hd_fill_2  FILLER_59_82
timestamp 1586364061
transform 1 0 8648 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_60_75
timestamp 1586364061
transform 1 0 8004 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 9660 0 1 34272
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 8832 0 1 34272
box -38 -48 222 592
use scs8hd_decap_6  FILLER_59_86
timestamp 1586364061
transform 1 0 9016 0 1 34272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_59_92
timestamp 1586364061
transform 1 0 9568 0 1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_60_87
timestamp 1586364061
transform 1 0 9108 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_60_91
timestamp 1586364061
transform 1 0 9476 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_60_93
timestamp 1586364061
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 10212 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_97
timestamp 1586364061
transform 1 0 10028 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_59_101
timestamp 1586364061
transform 1 0 10396 0 1 34272
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_60_105
timestamp 1586364061
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_113
timestamp 1586364061
transform 1 0 11500 0 1 34272
box -38 -48 774 592
use scs8hd_fill_1  FILLER_59_121
timestamp 1586364061
transform 1 0 12236 0 1 34272
box -38 -48 130 592
use scs8hd_decap_8  FILLER_59_123
timestamp 1586364061
transform 1 0 12420 0 1 34272
box -38 -48 774 592
use scs8hd_decap_12  FILLER_60_117
timestamp 1586364061
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use scs8hd_buf_2  _190_
timestamp 1586364061
transform 1 0 13156 0 1 34272
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 13708 0 1 34272
box -38 -48 222 592
use scs8hd_fill_2  FILLER_59_135
timestamp 1586364061
transform 1 0 13524 0 1 34272
box -38 -48 222 592
use scs8hd_decap_12  FILLER_60_129
timestamp 1586364061
transform 1 0 12972 0 -1 35360
box -38 -48 1142 592
use scs8hd_decap_3  PHY_119
timestamp 1586364061
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use scs8hd_decap_3  PHY_121
timestamp 1586364061
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use scs8hd_decap_6  FILLER_59_139
timestamp 1586364061
transform 1 0 13892 0 1 34272
box -38 -48 590 592
use scs8hd_fill_1  FILLER_59_145
timestamp 1586364061
transform 1 0 14444 0 1 34272
box -38 -48 130 592
use scs8hd_decap_4  FILLER_60_141
timestamp 1586364061
transform 1 0 14076 0 -1 35360
box -38 -48 406 592
use scs8hd_fill_1  FILLER_60_145
timestamp 1586364061
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use scs8hd_decap_3  PHY_122
timestamp 1586364061
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use scs8hd_decap_12  FILLER_61_3
timestamp 1586364061
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_15
timestamp 1586364061
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_27
timestamp 1586364061
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_39
timestamp 1586364061
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_51
timestamp 1586364061
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use scs8hd_fill_2  FILLER_61_59
timestamp 1586364061
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use scs8hd_decap_12  FILLER_61_62
timestamp 1586364061
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_74
timestamp 1586364061
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_86
timestamp 1586364061
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_98
timestamp 1586364061
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_61_110
timestamp 1586364061
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use scs8hd_decap_12  FILLER_61_123
timestamp 1586364061
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_61_135
timestamp 1586364061
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use scs8hd_decap_3  PHY_123
timestamp 1586364061
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  FILLER_61_143
timestamp 1586364061
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use scs8hd_decap_3  PHY_124
timestamp 1586364061
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_62_3
timestamp 1586364061
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_15
timestamp 1586364061
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_62_27
timestamp 1586364061
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_32
timestamp 1586364061
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_44
timestamp 1586364061
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_56
timestamp 1586364061
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_68
timestamp 1586364061
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_80
timestamp 1586364061
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_62_93
timestamp 1586364061
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_105
timestamp 1586364061
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_117
timestamp 1586364061
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_62_129
timestamp 1586364061
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use scs8hd_decap_3  PHY_125
timestamp 1586364061
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use scs8hd_decap_4  FILLER_62_141
timestamp 1586364061
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use scs8hd_fill_1  FILLER_62_145
timestamp 1586364061
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use scs8hd_decap_3  PHY_126
timestamp 1586364061
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use scs8hd_decap_12  FILLER_63_3
timestamp 1586364061
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_15
timestamp 1586364061
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_27
timestamp 1586364061
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_39
timestamp 1586364061
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_51
timestamp 1586364061
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use scs8hd_fill_2  FILLER_63_59
timestamp 1586364061
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use scs8hd_decap_12  FILLER_63_62
timestamp 1586364061
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_74
timestamp 1586364061
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_86
timestamp 1586364061
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_98
timestamp 1586364061
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_63_110
timestamp 1586364061
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use scs8hd_decap_12  FILLER_63_123
timestamp 1586364061
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_63_135
timestamp 1586364061
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use scs8hd_decap_3  PHY_127
timestamp 1586364061
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  FILLER_63_143
timestamp 1586364061
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use scs8hd_decap_3  PHY_128
timestamp 1586364061
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use scs8hd_decap_12  FILLER_64_3
timestamp 1586364061
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_15
timestamp 1586364061
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_64_27
timestamp 1586364061
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_12  FILLER_64_32
timestamp 1586364061
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_44
timestamp 1586364061
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_56
timestamp 1586364061
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_63
timestamp 1586364061
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_75
timestamp 1586364061
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_87
timestamp 1586364061
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_94
timestamp 1586364061
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_64_106
timestamp 1586364061
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use scs8hd_decap_6  FILLER_64_118
timestamp 1586364061
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use scs8hd_decap_12  FILLER_64_125
timestamp 1586364061
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_64_137
timestamp 1586364061
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use scs8hd_decap_3  PHY_129
timestamp 1586364061
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use scs8hd_fill_1  FILLER_64_145
timestamp 1586364061
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal2 s 6182 0 6238 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 6734 0 6790 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 7378 0 7434 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 7930 0 7986 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 8574 0 8630 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 9126 0 9182 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 9770 0 9826 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 294 0 350 480 6 chany_bottom_in[0]
port 7 nsew default input
rlabel metal2 s 846 0 902 480 6 chany_bottom_in[1]
port 8 nsew default input
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_in[2]
port 9 nsew default input
rlabel metal2 s 2042 0 2098 480 6 chany_bottom_in[3]
port 10 nsew default input
rlabel metal2 s 2594 0 2650 480 6 chany_bottom_in[4]
port 11 nsew default input
rlabel metal2 s 3238 0 3294 480 6 chany_bottom_in[5]
port 12 nsew default input
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_in[6]
port 13 nsew default input
rlabel metal2 s 4434 0 4490 480 6 chany_bottom_in[7]
port 14 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[8]
port 15 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_out[0]
port 16 nsew default tristate
rlabel metal2 s 11518 0 11574 480 6 chany_bottom_out[1]
port 17 nsew default tristate
rlabel metal2 s 12070 0 12126 480 6 chany_bottom_out[2]
port 18 nsew default tristate
rlabel metal2 s 12714 0 12770 480 6 chany_bottom_out[3]
port 19 nsew default tristate
rlabel metal2 s 13266 0 13322 480 6 chany_bottom_out[4]
port 20 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_out[5]
port 21 nsew default tristate
rlabel metal2 s 14462 0 14518 480 6 chany_bottom_out[6]
port 22 nsew default tristate
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_out[7]
port 23 nsew default tristate
rlabel metal2 s 15658 0 15714 480 6 chany_bottom_out[8]
port 24 nsew default tristate
rlabel metal2 s 386 39520 442 40000 6 chany_top_in[0]
port 25 nsew default input
rlabel metal2 s 1214 39520 1270 40000 6 chany_top_in[1]
port 26 nsew default input
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_in[2]
port 27 nsew default input
rlabel metal2 s 3054 39520 3110 40000 6 chany_top_in[3]
port 28 nsew default input
rlabel metal2 s 3882 39520 3938 40000 6 chany_top_in[4]
port 29 nsew default input
rlabel metal2 s 4802 39520 4858 40000 6 chany_top_in[5]
port 30 nsew default input
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_in[6]
port 31 nsew default input
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_in[7]
port 32 nsew default input
rlabel metal2 s 7470 39520 7526 40000 6 chany_top_in[8]
port 33 nsew default input
rlabel metal2 s 8390 39520 8446 40000 6 chany_top_out[0]
port 34 nsew default tristate
rlabel metal2 s 9218 39520 9274 40000 6 chany_top_out[1]
port 35 nsew default tristate
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_out[2]
port 36 nsew default tristate
rlabel metal2 s 11058 39520 11114 40000 6 chany_top_out[3]
port 37 nsew default tristate
rlabel metal2 s 11886 39520 11942 40000 6 chany_top_out[4]
port 38 nsew default tristate
rlabel metal2 s 12806 39520 12862 40000 6 chany_top_out[5]
port 39 nsew default tristate
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_out[6]
port 40 nsew default tristate
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_out[7]
port 41 nsew default tristate
rlabel metal2 s 15474 39520 15530 40000 6 chany_top_out[8]
port 42 nsew default tristate
rlabel metal2 s 10322 0 10378 480 6 data_in
port 43 nsew default input
rlabel metal2 s 5630 0 5686 480 6 enable
port 44 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_grid_pin_0_
port 45 nsew default tristate
rlabel metal3 s 0 27344 480 27464 6 left_grid_pin_10_
port 46 nsew default tristate
rlabel metal3 s 0 32376 480 32496 6 left_grid_pin_12_
port 47 nsew default tristate
rlabel metal3 s 0 37408 480 37528 6 left_grid_pin_14_
port 48 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 left_grid_pin_2_
port 49 nsew default tristate
rlabel metal3 s 0 12384 480 12504 6 left_grid_pin_4_
port 50 nsew default tristate
rlabel metal3 s 0 17416 480 17536 6 left_grid_pin_6_
port 51 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 left_grid_pin_8_
port 52 nsew default tristate
rlabel metal3 s 15520 9936 16000 10056 6 right_grid_pin_3_
port 53 nsew default tristate
rlabel metal3 s 15520 29928 16000 30048 6 right_grid_pin_7_
port 54 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 vpwr
port 55 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 vgnd
port 56 nsew default input
<< end >>
