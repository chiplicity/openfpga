* NGSPICE file created from cbx_1__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

.subckt cbx_1__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_grid_pin_0_ bottom_grid_pin_4_ bottom_grid_pin_8_ chanx_left_in[0]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1] chanx_right_in[2]
+ chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6] chanx_right_in[7]
+ chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ data_in enable top_grid_pin_0_ top_grid_pin_10_ top_grid_pin_12_ top_grid_pin_14_
+ top_grid_pin_2_ top_grid_pin_4_ top_grid_pin_6_ top_grid_pin_8_ vpwr vgnd
XFILLER_10_328 vgnd vpwr scs8hd_decap_8
XFILLER_7_7 vpwr vgnd scs8hd_fill_2
XFILLER_18_406 vgnd vpwr scs8hd_fill_1
XFILLER_13_199 vgnd vpwr scs8hd_decap_3
XFILLER_13_177 vpwr vgnd scs8hd_fill_2
XANTENNA__113__B _149_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_1_.latch data_in mem_bottom_ipin_2.LATCH_1_.latch/Q _179_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_158 vpwr vgnd scs8hd_fill_2
XFILLER_10_169 vpwr vgnd scs8hd_fill_2
XFILLER_12_10 vpwr vgnd scs8hd_fill_2
XFILLER_2_357 vgnd vpwr scs8hd_decap_12
XFILLER_2_335 vgnd vpwr scs8hd_fill_1
XFILLER_2_313 vgnd vpwr scs8hd_decap_4
XFILLER_12_98 vgnd vpwr scs8hd_decap_3
XFILLER_18_258 vgnd vpwr scs8hd_decap_3
XANTENNA__108__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_162 vpwr vgnd scs8hd_fill_2
XANTENNA__124__A _124_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_4_.latch data_in mem_bottom_ipin_4.LATCH_4_.latch/Q _102_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__209__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
X_200_ chanx_right_in[0] chanx_left_out[0] vgnd vpwr scs8hd_buf_2
X_131_ _077_/A _077_/B _077_/C _113_/A _131_/X vgnd vpwr scs8hd_or4_4
XFILLER_2_154 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _107_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_20 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_114_ _113_/X _115_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_279 vpwr vgnd scs8hd_fill_2
XFILLER_11_297 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_2_.latch/Q mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__121__B _077_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_87 vgnd vpwr scs8hd_decap_6
XANTENNA__116__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__132__A _131_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_172 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _181_/HI mem_bottom_ipin_0.LATCH_5_.latch/Q
+ mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_13_315 vpwr vgnd scs8hd_fill_2
XFILLER_15_87 vpwr vgnd scs8hd_fill_2
XFILLER_13_359 vgnd vpwr scs8hd_fill_1
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_142 vgnd vpwr scs8hd_decap_8
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_10_ vgnd vpwr scs8hd_inv_1
XFILLER_8_396 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_5.LATCH_0_.latch data_in mem_bottom_ipin_5.LATCH_0_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_123 vpwr vgnd scs8hd_fill_2
XFILLER_9_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_369 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_7.LATCH_3_.latch data_in mem_bottom_ipin_7.LATCH_3_.latch/Q _135_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_215 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_391 vgnd vpwr scs8hd_decap_12
XANTENNA__140__A _139_/X vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_0_ vgnd vpwr scs8hd_inv_1
X_130_ _148_/A _125_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__119__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA__135__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_23 vpwr vgnd scs8hd_fill_2
XFILLER_9_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_221 vgnd vpwr scs8hd_decap_12
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
X_113_ _113_/A _149_/A _113_/X vgnd vpwr scs8hd_or2_4
XFILLER_11_254 vpwr vgnd scs8hd_fill_2
XFILLER_19_310 vpwr vgnd scs8hd_fill_2
XFILLER_15_7 vpwr vgnd scs8hd_fill_2
XANTENNA__121__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_6_280 vpwr vgnd scs8hd_fill_2
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_4_206 vgnd vpwr scs8hd_decap_8
XFILLER_16_324 vgnd vpwr scs8hd_decap_12
XFILLER_6_35 vpwr vgnd scs8hd_fill_2
XFILLER_3_272 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_66 vgnd vpwr scs8hd_decap_4
XFILLER_15_11 vpwr vgnd scs8hd_fill_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _125_/B vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_176 vgnd vpwr scs8hd_decap_8
XFILLER_16_154 vpwr vgnd scs8hd_fill_2
XANTENNA__143__A _125_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_4_.latch data_in mem_top_ipin_0.LATCH_4_.latch/Q _144_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_157 vpwr vgnd scs8hd_fill_2
XFILLER_5_301 vpwr vgnd scs8hd_fill_2
XFILLER_5_323 vpwr vgnd scs8hd_fill_2
XFILLER_5_345 vgnd vpwr scs8hd_fill_1
XFILLER_5_389 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A _148_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_105 vpwr vgnd scs8hd_fill_2
XFILLER_10_127 vgnd vpwr scs8hd_fill_1
XFILLER_10_149 vgnd vpwr scs8hd_decap_4
XFILLER_12_23 vgnd vpwr scs8hd_decap_6
XFILLER_12_45 vgnd vpwr scs8hd_decap_4
XFILLER_12_78 vpwr vgnd scs8hd_fill_2
XFILLER_2_337 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _153_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_120 vpwr vgnd scs8hd_fill_2
XFILLER_5_131 vpwr vgnd scs8hd_fill_2
XFILLER_5_175 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_293 vpwr vgnd scs8hd_fill_2
XFILLER_17_282 vpwr vgnd scs8hd_fill_2
XFILLER_15_208 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_252 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_285 vpwr vgnd scs8hd_fill_2
XANTENNA__135__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_46 vpwr vgnd scs8hd_fill_2
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__151__A _173_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_233 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_0.LATCH_4_.latch data_in mem_bottom_ipin_0.LATCH_4_.latch/Q _160_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_112_ _111_/X _149_/A vgnd vpwr scs8hd_buf_1
XFILLER_11_222 vpwr vgnd scs8hd_fill_2
XFILLER_19_377 vpwr vgnd scs8hd_fill_2
XANTENNA__146__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_91 vgnd vpwr scs8hd_fill_1
XFILLER_20_56 vgnd vpwr scs8hd_decap_6
XFILLER_4_229 vpwr vgnd scs8hd_fill_2
XFILLER_16_314 vgnd vpwr scs8hd_fill_1
XFILLER_6_25 vpwr vgnd scs8hd_fill_2
XFILLER_19_196 vgnd vpwr scs8hd_decap_6
Xmem_top_ipin_1.LATCH_0_.latch data_in _154_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_391 vgnd vpwr scs8hd_decap_4
XFILLER_15_380 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_15_56 vpwr vgnd scs8hd_fill_2
XFILLER_15_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_16_111 vgnd vpwr scs8hd_decap_4
XFILLER_0_298 vpwr vgnd scs8hd_fill_2
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_332 vgnd vpwr scs8hd_decap_4
XFILLER_12_383 vpwr vgnd scs8hd_fill_2
XANTENNA__143__B _145_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_365 vpwr vgnd scs8hd_fill_2
XFILLER_8_398 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_136 vpwr vgnd scs8hd_fill_2
XFILLER_5_357 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__154__A _154_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_162 vgnd vpwr scs8hd_fill_1
XFILLER_8_195 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_139 vgnd vpwr scs8hd_decap_8
XFILLER_2_327 vgnd vpwr scs8hd_decap_8
XFILLER_2_305 vgnd vpwr scs8hd_decap_6
XFILLER_5_7 vgnd vpwr scs8hd_fill_1
XFILLER_12_57 vgnd vpwr scs8hd_decap_6
XFILLER_18_206 vgnd vpwr scs8hd_decap_8
XFILLER_1_360 vgnd vpwr scs8hd_decap_6
Xmem_bottom_ipin_1.LATCH_0_.latch data_in mem_bottom_ipin_1.LATCH_0_.latch/Q _172_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A _149_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_404 vgnd vpwr scs8hd_decap_3
XFILLER_4_80 vpwr vgnd scs8hd_fill_2
XFILLER_2_113 vgnd vpwr scs8hd_decap_4
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_3.LATCH_3_.latch data_in mem_bottom_ipin_3.LATCH_3_.latch/Q _086_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__151__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_245 vgnd vpwr scs8hd_decap_3
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _155_/A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_201 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_111_ _077_/A address[4] _077_/C _111_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_227 vgnd vpwr scs8hd_decap_4
XFILLER_11_278 vpwr vgnd scs8hd_fill_2
XFILLER_19_367 vgnd vpwr scs8hd_decap_6
XANTENNA__146__B _145_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_293 vgnd vpwr scs8hd_decap_12
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__072__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_SLEEPB _104_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_252 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_120 vpwr vgnd scs8hd_fill_2
XFILLER_3_296 vpwr vgnd scs8hd_fill_2
XFILLER_3_285 vpwr vgnd scs8hd_fill_2
XFILLER_10_90 vpwr vgnd scs8hd_fill_2
XFILLER_19_153 vpwr vgnd scs8hd_fill_2
XANTENNA__157__A _077_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_2_.latch/Q mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__067__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_211 vgnd vpwr scs8hd_decap_6
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_311 vpwr vgnd scs8hd_fill_2
XFILLER_8_388 vgnd vpwr scs8hd_decap_8
XFILLER_12_351 vpwr vgnd scs8hd_fill_2
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_336 vgnd vpwr scs8hd_decap_3
XFILLER_8_174 vgnd vpwr scs8hd_decap_8
XFILLER_12_192 vgnd vpwr scs8hd_decap_3
XFILLER_4_380 vgnd vpwr scs8hd_decap_12
XANTENNA__170__A _089_/B vgnd vpwr scs8hd_diode_2
XANTENNA__080__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_2_317 vgnd vpwr scs8hd_fill_1
XFILLER_5_144 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB _176_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_199 vpwr vgnd scs8hd_fill_2
XFILLER_17_240 vgnd vpwr scs8hd_decap_4
XANTENNA__149__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__165__A _165_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_6.LATCH_2_.latch data_in mem_bottom_ipin_6.LATCH_2_.latch/Q _128_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_405 vpwr vgnd scs8hd_fill_2
XANTENNA__075__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_2_169 vgnd vpwr scs8hd_fill_1
XFILLER_14_243 vgnd vpwr scs8hd_decap_6
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__151__C _069_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_180 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_18_35 vgnd vpwr scs8hd_decap_12
X_110_ _148_/A _110_/B _110_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_235 vgnd vpwr scs8hd_decap_3
XFILLER_7_206 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _181_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__162__B _158_/X vgnd vpwr scs8hd_diode_2
XFILLER_1_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_404 vgnd vpwr scs8hd_decap_3
XFILLER_16_349 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__157__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_319 vgnd vpwr scs8hd_decap_4
XANTENNA__083__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_16_102 vgnd vpwr scs8hd_decap_3
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_341 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__168__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__078__A _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_39 vgnd vpwr scs8hd_fill_1
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _153_/A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__170__B _171_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_392 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__080__B _067_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_219 vgnd vpwr scs8hd_decap_8
XFILLER_5_101 vpwr vgnd scs8hd_fill_2
XFILLER_5_112 vpwr vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vpwr scs8hd_fill_1
XFILLER_17_252 vpwr vgnd scs8hd_fill_2
XANTENNA__149__C _069_/C vgnd vpwr scs8hd_diode_2
XANTENNA__165__B _149_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_4
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_159 vpwr vgnd scs8hd_fill_2
XFILLER_2_137 vgnd vpwr scs8hd_decap_3
XFILLER_2_126 vpwr vgnd scs8hd_fill_2
XFILLER_9_27 vpwr vgnd scs8hd_fill_2
X_186_ _186_/HI _186_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_91 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__176__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_281 vpwr vgnd scs8hd_fill_2
XFILLER_18_47 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_258 vgnd vpwr scs8hd_decap_3
XFILLER_1_3 vgnd vpwr scs8hd_decap_8
XFILLER_19_314 vgnd vpwr scs8hd_decap_12
XFILLER_19_303 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_251 vpwr vgnd scs8hd_fill_2
XFILLER_6_262 vpwr vgnd scs8hd_fill_2
X_169_ _103_/A _171_/B _169_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_291 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_380 vgnd vpwr scs8hd_decap_12
XFILLER_1_83 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_0_.latch/Q mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_17 vpwr vgnd scs8hd_fill_2
XFILLER_6_39 vpwr vgnd scs8hd_fill_2
XANTENNA__157__C address[3] vgnd vpwr scs8hd_diode_2
XANTENNA__173__B _173_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_48 vgnd vpwr scs8hd_decap_8
XFILLER_15_15 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vgnd vpwr scs8hd_decap_8
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_324 vpwr vgnd scs8hd_fill_2
XFILLER_8_346 vpwr vgnd scs8hd_fill_2
XFILLER_12_364 vgnd vpwr scs8hd_decap_3
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _171_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XANTENNA__094__A _093_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_29 vpwr vgnd scs8hd_fill_2
XFILLER_3_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_154 vgnd vpwr scs8hd_decap_6
XANTENNA__179__A _107_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_109 vpwr vgnd scs8hd_fill_2
XFILLER_12_49 vgnd vpwr scs8hd_fill_1
XANTENNA__080__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__089__A _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_17_297 vgnd vpwr scs8hd_decap_8
XFILLER_17_286 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_7 vpwr vgnd scs8hd_fill_2
XFILLER_14_289 vgnd vpwr scs8hd_decap_4
XFILLER_14_267 vpwr vgnd scs8hd_fill_2
X_185_ _185_/HI _185_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_215 vpwr vgnd scs8hd_fill_2
XANTENNA__176__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA__192__A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__086__B _103_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_2.LATCH_2_.latch data_in mem_bottom_ipin_2.LATCH_2_.latch/Q _178_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_326 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
X_168_ _101_/A _171_/B _168_/Y vgnd vpwr scs8hd_nor2_4
X_099_ _098_/X _110_/B vgnd vpwr scs8hd_buf_1
XFILLER_18_392 vgnd vpwr scs8hd_decap_4
XFILLER_1_62 vgnd vpwr scs8hd_decap_4
XFILLER_1_95 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _182_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_5_.latch data_in mem_bottom_ipin_4.LATCH_5_.latch/Q _100_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__097__A address[5] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_3_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
XFILLER_6_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_3
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XFILLER_19_112 vgnd vpwr scs8hd_decap_8
XFILLER_19_91 vgnd vpwr scs8hd_decap_12
XFILLER_15_351 vpwr vgnd scs8hd_fill_2
XFILLER_15_340 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__157__D _165_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_38 vgnd vpwr scs8hd_fill_1
XFILLER_16_115 vgnd vpwr scs8hd_fill_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_159 vpwr vgnd scs8hd_fill_2
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_332 vgnd vpwr scs8hd_decap_4
XFILLER_12_387 vpwr vgnd scs8hd_fill_2
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_369 vpwr vgnd scs8hd_fill_2
XFILLER_12_398 vgnd vpwr scs8hd_decap_8
XFILLER_15_170 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_7_380 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_118 vpwr vgnd scs8hd_fill_2
XFILLER_5_306 vpwr vgnd scs8hd_fill_2
XFILLER_8_133 vgnd vpwr scs8hd_decap_8
XFILLER_8_144 vgnd vpwr scs8hd_decap_3
XFILLER_12_173 vgnd vpwr scs8hd_fill_1
XFILLER_4_350 vgnd vpwr scs8hd_decap_4
XFILLER_4_361 vgnd vpwr scs8hd_fill_1
XFILLER_8_199 vgnd vpwr scs8hd_decap_4
XANTENNA__179__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA__195__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__089__B _089_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_320 vpwr vgnd scs8hd_fill_2
XFILLER_5_158 vpwr vgnd scs8hd_fill_2
XFILLER_17_265 vpwr vgnd scs8hd_fill_2
XFILLER_17_232 vgnd vpwr scs8hd_decap_6
XFILLER_4_40 vgnd vpwr scs8hd_fill_1
XFILLER_4_84 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_0_.latch/Q mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_257 vgnd vpwr scs8hd_fill_1
X_184_ _184_/HI _184_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_161 vpwr vgnd scs8hd_fill_2
XFILLER_1_172 vgnd vpwr scs8hd_decap_8
Xmem_bottom_ipin_5.LATCH_1_.latch data_in mem_bottom_ipin_5.LATCH_1_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_249 vgnd vpwr scs8hd_decap_12
XFILLER_9_294 vgnd vpwr scs8hd_decap_4
XFILLER_11_205 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_338 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
X_098_ _077_/A address[4] address[3] _113_/A _098_/X vgnd vpwr scs8hd_or4_4
Xmem_bottom_ipin_7.LATCH_4_.latch data_in mem_bottom_ipin_7.LATCH_4_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_167_ _159_/A _171_/B _167_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_2_ vgnd vpwr scs8hd_inv_1
XANTENNA__097__B _097_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_289 vpwr vgnd scs8hd_fill_2
XFILLER_3_256 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_19_157 vgnd vpwr scs8hd_decap_4
XFILLER_19_135 vgnd vpwr scs8hd_decap_12
XFILLER_19_70 vgnd vpwr scs8hd_decap_8
XFILLER_15_363 vgnd vpwr scs8hd_decap_3
XANTENNA__198__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_15_28 vgnd vpwr scs8hd_decap_4
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_7 vpwr vgnd scs8hd_fill_2
XFILLER_15_193 vpwr vgnd scs8hd_fill_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_7_392 vgnd vpwr scs8hd_decap_4
XFILLER_17_403 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_185 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ _156_/A mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB _179_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_406 vgnd vpwr scs8hd_fill_1
XFILLER_17_211 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_183_ _183_/HI _183_/LO vgnd vpwr scs8hd_conb_1
XFILLER_13_83 vpwr vgnd scs8hd_fill_2
Xmem_top_ipin_0.LATCH_5_.latch data_in mem_top_ipin_0.LATCH_5_.latch/Q _143_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_9_240 vpwr vgnd scs8hd_fill_2
XFILLER_9_262 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_166_ _165_/X _171_/B vgnd vpwr scs8hd_buf_1
XFILLER_6_232 vgnd vpwr scs8hd_decap_8
XFILLER_6_276 vpwr vgnd scs8hd_fill_2
X_097_ address[5] _097_/B _113_/A vgnd vpwr scs8hd_nand2_4
XFILLER_1_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _183_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_309 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_268 vpwr vgnd scs8hd_fill_2
XFILLER_3_224 vpwr vgnd scs8hd_fill_2
XFILLER_3_202 vgnd vpwr scs8hd_fill_1
XFILLER_19_147 vgnd vpwr scs8hd_decap_3
XFILLER_19_103 vpwr vgnd scs8hd_fill_2
XFILLER_10_84 vgnd vpwr scs8hd_decap_4
X_149_ _149_/A _149_/B _069_/C _149_/Y vgnd vpwr scs8hd_nor3_4
Xmux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_249 vgnd vpwr scs8hd_decap_12
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_312 vgnd vpwr scs8hd_fill_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_0.LATCH_5_.latch data_in mem_bottom_ipin_0.LATCH_5_.latch/Q _159_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_345 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_0_.latch/Q mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_3 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_319 vpwr vgnd scs8hd_fill_2
XFILLER_16_72 vgnd vpwr scs8hd_decap_3
XFILLER_8_102 vgnd vpwr scs8hd_decap_3
XFILLER_8_113 vpwr vgnd scs8hd_fill_2
XFILLER_4_396 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_1.LATCH_1_.latch data_in _153_/A _149_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_105 vgnd vpwr scs8hd_decap_4
XFILLER_5_116 vpwr vgnd scs8hd_fill_2
XFILLER_5_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_182_ _182_/HI _182_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_226 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_62 vpwr vgnd scs8hd_fill_2
XFILLER_13_95 vgnd vpwr scs8hd_decap_4
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XANTENNA__100__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_207 vgnd vpwr scs8hd_decap_8
XFILLER_13_292 vgnd vpwr scs8hd_fill_1
XFILLER_9_230 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_SLEEPB _137_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_218 vpwr vgnd scs8hd_fill_2
XFILLER_10_262 vgnd vpwr scs8hd_fill_1
XFILLER_10_273 vpwr vgnd scs8hd_fill_2
X_165_ _165_/A _149_/A _165_/X vgnd vpwr scs8hd_or2_4
X_096_ address[6] _097_/B vgnd vpwr scs8hd_inv_8
XFILLER_6_255 vpwr vgnd scs8hd_fill_2
XFILLER_6_266 vgnd vpwr scs8hd_decap_8
Xmem_bottom_ipin_1.LATCH_1_.latch data_in mem_bottom_ipin_1.LATCH_1_.latch/Q _171_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_3_236 vgnd vpwr scs8hd_fill_1
XFILLER_10_41 vpwr vgnd scs8hd_fill_2
XFILLER_10_63 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ _154_/A mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_15_398 vpwr vgnd scs8hd_fill_2
XFILLER_15_387 vpwr vgnd scs8hd_fill_2
XFILLER_15_376 vpwr vgnd scs8hd_fill_2
X_148_ _148_/A _145_/B _148_/Y vgnd vpwr scs8hd_nor2_4
X_079_ _125_/A _079_/B _079_/Y vgnd vpwr scs8hd_nor2_4
Xmem_bottom_ipin_3.LATCH_4_.latch data_in mem_bottom_ipin_3.LATCH_4_.latch/Q _082_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_107 vpwr vgnd scs8hd_fill_2
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_324 vpwr vgnd scs8hd_fill_2
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_328 vpwr vgnd scs8hd_fill_2
XFILLER_15_151 vpwr vgnd scs8hd_fill_2
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_42 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
XFILLER_7_361 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_SLEEPB _118_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_84 vgnd vpwr scs8hd_decap_3
XFILLER_12_165 vpwr vgnd scs8hd_fill_2
XFILLER_4_320 vgnd vpwr scs8hd_decap_6
XFILLER_4_364 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _103_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_367 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_8
XFILLER_4_21 vgnd vpwr scs8hd_decap_8
XFILLER_4_76 vpwr vgnd scs8hd_fill_2
XFILLER_4_183 vpwr vgnd scs8hd_fill_2
XFILLER_4_194 vgnd vpwr scs8hd_decap_8
Xmux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _155_/Y mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_109 vpwr vgnd scs8hd_fill_2
X_181_ _181_/HI _181_/LO vgnd vpwr scs8hd_conb_1
XFILLER_14_249 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__100__B _110_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__201__A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_0_.latch/Q mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_0_.latch data_in mem_bottom_ipin_4.LATCH_0_.latch/Q _110_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_241 vgnd vpwr scs8hd_decap_4
XFILLER_10_285 vgnd vpwr scs8hd_decap_4
X_164_ _148_/A _158_/X _164_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
X_095_ _079_/B _095_/B _095_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__111__A _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_99 vpwr vgnd scs8hd_fill_2
XFILLER_18_396 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _184_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_248 vpwr vgnd scs8hd_fill_2
XFILLER_10_53 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_6.LATCH_3_.latch data_in mem_bottom_ipin_6.LATCH_3_.latch/Q _127_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_19_62 vgnd vpwr scs8hd_fill_1
XFILLER_15_355 vpwr vgnd scs8hd_fill_2
XFILLER_15_344 vpwr vgnd scs8hd_fill_2
X_147_ _107_/X _145_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A _162_/A vgnd vpwr scs8hd_diode_2
X_078_ _078_/A _079_/B vgnd vpwr scs8hd_buf_1
XFILLER_18_3 vgnd vpwr scs8hd_decap_6
XFILLER_18_171 vgnd vpwr scs8hd_decap_12
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_307 vpwr vgnd scs8hd_fill_2
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_369 vgnd vpwr scs8hd_decap_3
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_174 vgnd vpwr scs8hd_decap_3
XFILLER_11_380 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_41 vpwr vgnd scs8hd_fill_2
XFILLER_16_30 vgnd vpwr scs8hd_fill_1
XFILLER_4_310 vgnd vpwr scs8hd_fill_1
XFILLER_4_398 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__204__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_1_324 vgnd vpwr scs8hd_decap_12
XFILLER_1_379 vgnd vpwr scs8hd_decap_12
XFILLER_17_269 vpwr vgnd scs8hd_fill_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_8
XFILLER_4_11 vgnd vpwr scs8hd_fill_1
XANTENNA__114__A _113_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_99 vgnd vpwr scs8hd_decap_4
XFILLER_4_140 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_0_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_206 vgnd vpwr scs8hd_decap_6
X_180_ _095_/B _178_/B _180_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_13_53 vgnd vpwr scs8hd_decap_6
XFILLER_1_132 vgnd vpwr scs8hd_decap_8
XFILLER_1_143 vpwr vgnd scs8hd_fill_2
XFILLER_1_165 vgnd vpwr scs8hd_decap_4
XFILLER_13_250 vpwr vgnd scs8hd_fill_2
XANTENNA__109__A _095_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_210 vgnd vpwr scs8hd_fill_1
XFILLER_9_298 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
X_163_ _107_/X _158_/X _163_/Y vgnd vpwr scs8hd_nor2_4
X_094_ _093_/X _095_/B vgnd vpwr scs8hd_buf_1
XANTENNA__111__B address[4] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_8_ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_353 vgnd vpwr scs8hd_fill_1
XFILLER_18_331 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_205 vgnd vpwr scs8hd_decap_12
XFILLER_10_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_7.LATCH_3_.latch/Q mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_323 vpwr vgnd scs8hd_fill_2
XANTENNA__106__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA__122__A _121_/X vgnd vpwr scs8hd_diode_2
X_077_ _077_/A _077_/B _077_/C _165_/A _078_/A vgnd vpwr scs8hd_or4_4
X_146_ _162_/A _145_/B _146_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_293 vgnd vpwr scs8hd_decap_12
XFILLER_18_183 vgnd vpwr scs8hd_decap_12
XANTENNA__207__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_337 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _153_/Y mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_142 vpwr vgnd scs8hd_fill_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_197 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_11 vgnd vpwr scs8hd_decap_3
XFILLER_7_88 vpwr vgnd scs8hd_fill_2
XANTENNA__117__A _145_/A vgnd vpwr scs8hd_diode_2
X_129_ _107_/X _125_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_4_300 vgnd vpwr scs8hd_decap_8
XFILLER_8_149 vgnd vpwr scs8hd_decap_4
XFILLER_12_134 vgnd vpwr scs8hd_decap_8
XFILLER_12_145 vgnd vpwr scs8hd_decap_6
XFILLER_12_189 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_333 vgnd vpwr scs8hd_fill_1
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_0_.latch/Q mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_336 vgnd vpwr scs8hd_decap_12
XFILLER_17_248 vpwr vgnd scs8hd_fill_2
XFILLER_4_152 vgnd vpwr scs8hd_fill_1
XFILLER_4_163 vgnd vpwr scs8hd_decap_3
XANTENNA__130__A _148_/A vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_0_.latch data_in mem_top_ipin_0.LATCH_0_.latch/Q _148_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_406 vgnd vpwr scs8hd_fill_1
XFILLER_13_21 vgnd vpwr scs8hd_decap_4
XFILLER_13_32 vpwr vgnd scs8hd_fill_2
XFILLER_1_155 vgnd vpwr scs8hd_fill_1
XFILLER_13_295 vpwr vgnd scs8hd_fill_2
XFILLER_13_273 vpwr vgnd scs8hd_fill_2
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
XFILLER_9_277 vpwr vgnd scs8hd_fill_2
XANTENNA__125__A _125_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_SLEEPB _126_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_1_.latch/Q mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
X_162_ _162_/A _158_/X _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_265 vgnd vpwr scs8hd_decap_8
X_093_ address[1] address[2] address[0] _093_/X vgnd vpwr scs8hd_or3_4
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__111__C _077_/C vgnd vpwr scs8hd_diode_2
XFILLER_1_13 vgnd vpwr scs8hd_decap_12
XFILLER_18_398 vgnd vpwr scs8hd_decap_8
XFILLER_1_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_280 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _185_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_239 vgnd vpwr scs8hd_decap_3
XFILLER_3_228 vgnd vpwr scs8hd_decap_8
XFILLER_3_217 vpwr vgnd scs8hd_fill_2
X_145_ _145_/A _145_/B _145_/Y vgnd vpwr scs8hd_nor2_4
X_076_ address[5] address[6] _165_/A vgnd vpwr scs8hd_or2_4
XFILLER_2_261 vgnd vpwr scs8hd_decap_12
XFILLER_2_250 vgnd vpwr scs8hd_decap_8
Xmem_bottom_ipin_0.LATCH_0_.latch data_in mem_bottom_ipin_0.LATCH_0_.latch/Q _164_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_18_195 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vpwr scs8hd_decap_3
X_128_ _162_/A _125_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__133__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_342 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_2.LATCH_3_.latch data_in mem_bottom_ipin_2.LATCH_3_.latch/Q _177_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__117__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_393 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_117 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__128__A _162_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_348 vgnd vpwr scs8hd_decap_12
XANTENNA__130__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_293 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_6.LATCH_3_.latch/Q mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__125__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_234 vgnd vpwr scs8hd_decap_4
XFILLER_9_245 vpwr vgnd scs8hd_fill_2
XANTENNA__141__A _077_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_ipin_0.LATCH_4_.latch/Q mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr
+ scs8hd_ebufn_2
X_161_ _145_/A _158_/X _161_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_215 vpwr vgnd scs8hd_fill_2
XFILLER_10_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_10_299 vgnd vpwr scs8hd_fill_1
X_092_ _079_/B _107_/A _092_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_25 vgnd vpwr scs8hd_decap_12
XANTENNA__136__A _162_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _156_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_10_23 vpwr vgnd scs8hd_fill_2
XFILLER_10_45 vgnd vpwr scs8hd_decap_8
XFILLER_10_67 vpwr vgnd scs8hd_fill_2
XFILLER_19_108 vpwr vgnd scs8hd_fill_2
X_144_ _144_/A _145_/B _144_/Y vgnd vpwr scs8hd_nor2_4
X_075_ address[3] _077_/C vgnd vpwr scs8hd_inv_8
XFILLER_2_273 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_5.LATCH_2_.latch data_in mem_bottom_ipin_5.LATCH_2_.latch/Q _118_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_328 vpwr vgnd scs8hd_fill_2
XFILLER_15_100 vpwr vgnd scs8hd_fill_2
XFILLER_15_166 vpwr vgnd scs8hd_fill_2
XFILLER_15_111 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
X_127_ _145_/A _125_/B _127_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_46 vpwr vgnd scs8hd_fill_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_7_321 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_376 vpwr vgnd scs8hd_fill_2
XFILLER_16_3 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_7.LATCH_5_.latch data_in mem_bottom_ipin_7.LATCH_5_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_22 vgnd vpwr scs8hd_decap_6
XFILLER_8_107 vgnd vpwr scs8hd_decap_3
XFILLER_12_103 vgnd vpwr scs8hd_decap_3
XFILLER_12_169 vgnd vpwr scs8hd_decap_4
XFILLER_4_346 vpwr vgnd scs8hd_fill_2
XFILLER_4_357 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_368 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _125_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_151 vgnd vpwr scs8hd_decap_4
XFILLER_7_173 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_1_.latch/Q mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_291 vgnd vpwr scs8hd_decap_12
XFILLER_17_228 vpwr vgnd scs8hd_fill_2
XFILLER_9_405 vpwr vgnd scs8hd_fill_2
XFILLER_4_187 vgnd vpwr scs8hd_decap_4
XANTENNA__139__A address[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_9_213 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__141__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_091_ _091_/A _107_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_160_ _144_/A _158_/X _160_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_37 vgnd vpwr scs8hd_decap_12
XFILLER_1_59 vpwr vgnd scs8hd_fill_2
XANTENNA__136__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _173_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_271 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _186_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_66 vpwr vgnd scs8hd_fill_2
XFILLER_15_359 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_143_ _125_/A _145_/B _143_/Y vgnd vpwr scs8hd_nor2_4
X_074_ address[4] _077_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__147__A _107_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_373 vgnd vpwr scs8hd_decap_12
XFILLER_15_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_7_25 vpwr vgnd scs8hd_fill_2
XFILLER_7_300 vpwr vgnd scs8hd_fill_2
XFILLER_11_340 vpwr vgnd scs8hd_fill_2
XFILLER_11_362 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_5.LATCH_3_.latch/Q mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
X_126_ _144_/A _125_/B _126_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_388 vpwr vgnd scs8hd_fill_2
XFILLER_7_399 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ _156_/Y mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_89 vgnd vpwr scs8hd_decap_3
XFILLER_16_67 vgnd vpwr scs8hd_decap_3
XFILLER_16_45 vgnd vpwr scs8hd_decap_12
XANTENNA__144__B _145_/B vgnd vpwr scs8hd_diode_2
X_109_ _095_/B _148_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__160__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_1_306 vgnd vpwr scs8hd_decap_12
XFILLER_8_90 vpwr vgnd scs8hd_fill_2
XANTENNA__070__A _069_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_59 vgnd vpwr scs8hd_decap_6
XFILLER_4_144 vgnd vpwr scs8hd_decap_8
XANTENNA__139__B _097_/B vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _155_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_79 vpwr vgnd scs8hd_fill_2
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_1_147 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_6 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_0_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_169 vgnd vpwr scs8hd_fill_1
XFILLER_13_254 vpwr vgnd scs8hd_fill_2
XFILLER_9_258 vpwr vgnd scs8hd_fill_2
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XANTENNA__141__C address[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_14_ vgnd vpwr scs8hd_inv_1
X_090_ address[1] address[2] _069_/C _091_/A vgnd vpwr scs8hd_or3_4
XFILLER_6_206 vgnd vpwr scs8hd_decap_6
XFILLER_10_202 vpwr vgnd scs8hd_fill_2
XFILLER_10_224 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vpwr vgnd scs8hd_fill_2
XFILLER_18_368 vgnd vpwr scs8hd_decap_12
XFILLER_18_357 vgnd vpwr scs8hd_decap_8
XFILLER_18_335 vgnd vpwr scs8hd_fill_1
XFILLER_1_49 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__152__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_261 vgnd vpwr scs8hd_fill_1
XFILLER_19_78 vpwr vgnd scs8hd_fill_2
XFILLER_19_23 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_327 vpwr vgnd scs8hd_fill_2
X_142_ _142_/A _145_/B vgnd vpwr scs8hd_buf_1
X_073_ _121_/A _077_/A vgnd vpwr scs8hd_buf_1
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_1_.latch/Q mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_8
XANTENNA__147__B _145_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_371 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A _107_/X vgnd vpwr scs8hd_diode_2
XFILLER_2_81 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_308 vgnd vpwr scs8hd_decap_4
XFILLER_20_385 vgnd vpwr scs8hd_decap_12
XANTENNA__073__A _121_/A vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_8_ vgnd vpwr scs8hd_inv_1
X_125_ _125_/A _125_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_15_179 vpwr vgnd scs8hd_fill_2
XANTENNA__158__A _157_/X vgnd vpwr scs8hd_diode_2
XFILLER_14_190 vpwr vgnd scs8hd_fill_2
XFILLER_16_57 vgnd vpwr scs8hd_fill_1
XANTENNA__068__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_4_326 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_1.LATCH_2_.latch data_in mem_bottom_ipin_1.LATCH_2_.latch/Q _170_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_108_ _107_/X _110_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_197 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_160 vpwr vgnd scs8hd_fill_2
XANTENNA__160__B _158_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_3.LATCH_5_.latch data_in mem_bottom_ipin_3.LATCH_5_.latch/Q _079_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_112 vpwr vgnd scs8hd_fill_2
XFILLER_4_123 vpwr vgnd scs8hd_fill_2
XFILLER_0_373 vgnd vpwr scs8hd_decap_12
XFILLER_16_241 vgnd vpwr scs8hd_decap_3
XFILLER_16_285 vgnd vpwr scs8hd_decap_8
XFILLER_16_252 vgnd vpwr scs8hd_decap_3
XANTENNA__171__A _107_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_0_.latch/Q mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_406 vgnd vpwr scs8hd_fill_1
XFILLER_13_36 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__081__A _080_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_299 vgnd vpwr scs8hd_decap_4
XFILLER_13_288 vgnd vpwr scs8hd_decap_4
XFILLER_9_226 vpwr vgnd scs8hd_fill_2
XANTENNA__141__D _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__166__A _165_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__076__A address[5] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_4.LATCH_3_.latch/Q mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_247 vpwr vgnd scs8hd_fill_2
XFILLER_10_258 vgnd vpwr scs8hd_decap_4
Xmux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ _154_/Y mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__152__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_284 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_391 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_35 vgnd vpwr scs8hd_decap_12
XFILLER_15_306 vgnd vpwr scs8hd_decap_4
X_141_ _077_/A address[4] address[3] _149_/B _142_/A vgnd vpwr scs8hd_or4_4
X_072_ enable _121_/A vgnd vpwr scs8hd_inv_8
XFILLER_18_133 vgnd vpwr scs8hd_decap_12
XFILLER_18_122 vpwr vgnd scs8hd_fill_2
XFILLER_18_111 vgnd vpwr scs8hd_decap_8
XFILLER_2_276 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__163__B _158_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_6
XFILLER_2_60 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_342 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_397 vgnd vpwr scs8hd_decap_6
XFILLER_15_147 vpwr vgnd scs8hd_fill_2
XFILLER_7_346 vpwr vgnd scs8hd_fill_2
XFILLER_7_357 vpwr vgnd scs8hd_fill_2
X_124_ _124_/A _125_/B vgnd vpwr scs8hd_buf_1
XFILLER_11_397 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_91 vpwr vgnd scs8hd_fill_2
XANTENNA__174__A _173_/X vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_1_.latch data_in mem_bottom_ipin_4.LATCH_1_.latch/Q _108_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_117 vgnd vpwr scs8hd_decap_8
XANTENNA__084__A _084_/A vgnd vpwr scs8hd_diode_2
X_107_ _107_/A _107_/X vgnd vpwr scs8hd_buf_1
XFILLER_3_371 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_6.LATCH_4_.latch data_in mem_bottom_ipin_6.LATCH_4_.latch/Q _126_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
XANTENNA__169__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_81 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_385 vgnd vpwr scs8hd_decap_12
XFILLER_4_168 vgnd vpwr scs8hd_decap_6
XFILLER_16_264 vgnd vpwr scs8hd_decap_3
XFILLER_16_297 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _155_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__171__B _171_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_1_.latch/Q mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_13_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB _177_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_82 vpwr vgnd scs8hd_fill_2
XANTENNA__076__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_6_219 vpwr vgnd scs8hd_fill_2
XANTENNA__092__A _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_337 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _103_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vpwr vgnd scs8hd_fill_2
XFILLER_19_47 vgnd vpwr scs8hd_decap_12
XANTENNA__087__A _084_/A vgnd vpwr scs8hd_diode_2
X_140_ _139_/X _149_/B vgnd vpwr scs8hd_buf_1
X_071_ _159_/A _125_/A vgnd vpwr scs8hd_buf_1
XFILLER_2_288 vgnd vpwr scs8hd_decap_3
XFILLER_18_145 vgnd vpwr scs8hd_decap_8
XFILLER_18_101 vgnd vpwr scs8hd_fill_1
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_354 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_7.LATCH_0_.latch data_in mem_bottom_ipin_7.LATCH_0_.latch/Q _138_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_115 vgnd vpwr scs8hd_decap_4
XFILLER_15_104 vpwr vgnd scs8hd_fill_2
XFILLER_11_321 vpwr vgnd scs8hd_fill_2
X_123_ _113_/A _173_/B _124_/A vgnd vpwr scs8hd_or2_4
XFILLER_7_325 vpwr vgnd scs8hd_fill_2
XFILLER_11_376 vpwr vgnd scs8hd_fill_2
XFILLER_11_70 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_7 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_0_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_162 vgnd vpwr scs8hd_fill_1
XANTENNA__084__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB _160_/Y vgnd vpwr scs8hd_diode_2
X_106_ _162_/A _110_/B _106_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_155 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_184 vgnd vpwr scs8hd_decap_4
XFILLER_3_383 vgnd vpwr scs8hd_decap_12
XANTENNA__169__B _171_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_1_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_3.LATCH_3_.latch/Q mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__079__B _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_405 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__095__A _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_4_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_397 vgnd vpwr scs8hd_decap_6
XFILLER_0_342 vgnd vpwr scs8hd_decap_12
XFILLER_16_221 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_3_191 vpwr vgnd scs8hd_fill_2
XFILLER_3_180 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_0_ vgnd vpwr scs8hd_inv_1
XFILLER_1_106 vgnd vpwr scs8hd_decap_6
XFILLER_13_49 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_224 vpwr vgnd scs8hd_fill_2
XFILLER_5_401 vgnd vpwr scs8hd_decap_6
XFILLER_9_206 vgnd vpwr scs8hd_decap_4
XANTENNA__092__B _107_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_7.LATCH_4_.latch/Q mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_349 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_242 vpwr vgnd scs8hd_fill_2
XFILLER_14_81 vpwr vgnd scs8hd_fill_2
XFILLER_5_297 vpwr vgnd scs8hd_fill_2
XFILLER_17_371 vgnd vpwr scs8hd_fill_1
XANTENNA__177__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA__193__A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _188_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__087__B address[2] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_1_.latch data_in mem_top_ipin_0.LATCH_1_.latch/Q _147_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_070_ _069_/X _159_/A vgnd vpwr scs8hd_buf_1
XFILLER_4_3 vgnd vpwr scs8hd_decap_8
XFILLER_14_396 vgnd vpwr scs8hd_fill_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
X_199_ chanx_right_in[1] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_366 vgnd vpwr scs8hd_decap_6
XFILLER_20_311 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__098__A _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_138 vpwr vgnd scs8hd_fill_2
XFILLER_7_304 vgnd vpwr scs8hd_fill_1
XFILLER_11_344 vgnd vpwr scs8hd_decap_3
X_122_ _121_/X _173_/B vgnd vpwr scs8hd_buf_1
XFILLER_7_29 vpwr vgnd scs8hd_fill_2
XFILLER_14_171 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_1_.latch/Q mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__084__C _069_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_185 vgnd vpwr scs8hd_fill_1
XFILLER_4_329 vgnd vpwr scs8hd_decap_4
X_105_ _089_/B _162_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_112 vgnd vpwr scs8hd_decap_4
XFILLER_7_134 vpwr vgnd scs8hd_fill_2
XFILLER_3_395 vgnd vpwr scs8hd_decap_12
XFILLER_19_230 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_1_.latch data_in mem_bottom_ipin_0.LATCH_1_.latch/Q _163_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__095__B _095_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_354 vgnd vpwr scs8hd_decap_12
XFILLER_16_233 vgnd vpwr scs8hd_decap_8
XFILLER_3_170 vgnd vpwr scs8hd_decap_4
XANTENNA__196__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_4_.latch data_in mem_bottom_ipin_2.LATCH_4_.latch/Q _176_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_17 vpwr vgnd scs8hd_fill_2
XFILLER_13_28 vpwr vgnd scs8hd_fill_2
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_2_.latch/Q mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_236 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_13_269 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_4
XFILLER_8_251 vpwr vgnd scs8hd_fill_2
XFILLER_10_206 vgnd vpwr scs8hd_decap_3
XFILLER_10_228 vpwr vgnd scs8hd_fill_2
XFILLER_6_7 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_0_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_60 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_254 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__087__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_213 vgnd vpwr scs8hd_fill_1
XFILLER_14_375 vpwr vgnd scs8hd_fill_2
XPHY_70 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ chanx_right_in[2] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_2.LATCH_3_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
XFILLER_20_323 vgnd vpwr scs8hd_decap_12
XFILLER_17_180 vgnd vpwr scs8hd_decap_3
XANTENNA__098__B address[4] vgnd vpwr scs8hd_diode_2
X_121_ _121_/A _077_/B address[3] _121_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_338 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_194 vgnd vpwr scs8hd_decap_3
XFILLER_6_360 vpwr vgnd scs8hd_fill_2
XFILLER_6_371 vgnd vpwr scs8hd_decap_8
XANTENNA__199__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_6_382 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _156_/Y vgnd vpwr
+ scs8hd_diode_2
X_104_ _145_/A _110_/B _104_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_175 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_3.LATCH_0_.latch data_in mem_bottom_ipin_3.LATCH_0_.latch/Q _095_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_330 vpwr vgnd scs8hd_fill_2
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XFILLER_19_264 vpwr vgnd scs8hd_fill_2
XFILLER_19_242 vpwr vgnd scs8hd_fill_2
XFILLER_19_220 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_6.LATCH_4_.latch/Q mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_311 vgnd vpwr scs8hd_decap_12
XFILLER_4_116 vpwr vgnd scs8hd_fill_2
XFILLER_4_127 vpwr vgnd scs8hd_fill_2
XFILLER_16_201 vpwr vgnd scs8hd_fill_2
XFILLER_0_366 vgnd vpwr scs8hd_decap_6
Xmem_bottom_ipin_5.LATCH_3_.latch data_in mem_bottom_ipin_5.LATCH_3_.latch/Q _117_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _189_/HI mem_top_ipin_0.LATCH_5_.latch/Q
+ mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_8_230 vgnd vpwr scs8hd_decap_4
XFILLER_8_285 vpwr vgnd scs8hd_fill_2
XFILLER_2_406 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_307 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_211 vpwr vgnd scs8hd_fill_2
XFILLER_5_277 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_362 vgnd vpwr scs8hd_decap_4
XFILLER_2_247 vgnd vpwr scs8hd_fill_1
XFILLER_2_258 vgnd vpwr scs8hd_fill_1
XFILLER_18_126 vgnd vpwr scs8hd_decap_4
XFILLER_14_354 vpwr vgnd scs8hd_fill_2
XPHY_71 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_60 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ chanx_right_in[3] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_14_398 vgnd vpwr scs8hd_decap_8
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_64 vpwr vgnd scs8hd_fill_2
XFILLER_20_335 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_380 vpwr vgnd scs8hd_fill_2
XANTENNA__098__C address[3] vgnd vpwr scs8hd_diode_2
Xmux_top_ipin_2.INVTX1_0_.scs8hd_inv_1 chanx_left_in[1] mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_306 vgnd vpwr scs8hd_decap_4
X_120_ _148_/A _115_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_350 vgnd vpwr scs8hd_decap_4
XFILLER_6_394 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_2_.latch/Q mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_18 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_187 vgnd vpwr scs8hd_decap_12
XFILLER_20_165 vgnd vpwr scs8hd_decap_12
X_103_ _103_/A _145_/A vgnd vpwr scs8hd_buf_1
XFILLER_7_158 vpwr vgnd scs8hd_fill_2
XFILLER_11_143 vpwr vgnd scs8hd_fill_2
XFILLER_8_41 vgnd vpwr scs8hd_decap_8
XFILLER_8_85 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_0_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_323 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_3.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB _180_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_1.LATCH_3_.latch/Q mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_120 vgnd vpwr scs8hd_decap_4
XFILLER_0_153 vpwr vgnd scs8hd_fill_2
XFILLER_8_297 vgnd vpwr scs8hd_fill_1
XFILLER_12_271 vpwr vgnd scs8hd_fill_2
XFILLER_5_20 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vpwr vgnd scs8hd_fill_2
XFILLER_5_86 vpwr vgnd scs8hd_fill_2
XFILLER_18_319 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_223 vpwr vgnd scs8hd_fill_2
XANTENNA__101__A _101_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_352 vgnd vpwr scs8hd_fill_1
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_14_388 vgnd vpwr scs8hd_decap_8
XFILLER_14_333 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_61 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_196_ chanx_right_in[4] chanx_left_out[4] vgnd vpwr scs8hd_buf_2
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_5.LATCH_4_.latch/Q mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_1_281 vgnd vpwr scs8hd_decap_12
XFILLER_2_54 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__D _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_119 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_ipin_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_325 vpwr vgnd scs8hd_fill_2
XFILLER_11_358 vpwr vgnd scs8hd_fill_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_8
XFILLER_11_52 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_152 vgnd vpwr scs8hd_fill_1
X_179_ _107_/A _178_/B _179_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_199 vgnd vpwr scs8hd_decap_6
XFILLER_20_177 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_406 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_102_ _144_/A _110_/B _102_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_ipin_0.INVTX1_0_.scs8hd_inv_1 chanx_left_in[3] mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_365 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_64 vpwr vgnd scs8hd_fill_2
XFILLER_6_192 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_1_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_335 vgnd vpwr scs8hd_decap_6
XFILLER_0_302 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_62 vgnd vpwr scs8hd_decap_6
XFILLER_16_269 vgnd vpwr scs8hd_decap_4
XFILLER_16_247 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_6_ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__104__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_280 vpwr vgnd scs8hd_fill_2
XFILLER_13_228 vgnd vpwr scs8hd_decap_3
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_5_10 vgnd vpwr scs8hd_fill_1
XFILLER_8_210 vpwr vgnd scs8hd_fill_2
XFILLER_8_243 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_1.LATCH_3_.latch data_in mem_bottom_ipin_1.LATCH_3_.latch/Q _169_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_43 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_52 vgnd vpwr scs8hd_decap_8
XFILLER_14_85 vgnd vpwr scs8hd_decap_4
XFILLER_14_96 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_2_.latch/Q mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_375 vpwr vgnd scs8hd_fill_2
XFILLER_19_19 vpwr vgnd scs8hd_fill_2
XFILLER_4_290 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XANTENNA__202__A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_SLEEPB _138_/Y vgnd vpwr scs8hd_diode_2
XPHY_40 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_62 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_51 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_195_ chanx_right_in[5] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_2_44 vgnd vpwr scs8hd_decap_8
XFILLER_1_293 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A _111_/X vgnd vpwr scs8hd_diode_2
XFILLER_17_194 vpwr vgnd scs8hd_fill_2
XFILLER_17_172 vpwr vgnd scs8hd_fill_2
XFILLER_2_99 vgnd vpwr scs8hd_fill_1
XFILLER_20_304 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_0_.latch/Q mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_393 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__107__A _107_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_186 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_178_ _089_/B _178_/B _178_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_20_112 vgnd vpwr scs8hd_fill_1
XFILLER_20_156 vgnd vpwr scs8hd_decap_6
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_0.LATCH_3_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_105 vgnd vpwr scs8hd_decap_4
XFILLER_7_138 vpwr vgnd scs8hd_fill_2
XFILLER_11_112 vgnd vpwr scs8hd_decap_4
XFILLER_11_123 vgnd vpwr scs8hd_decap_4
XFILLER_11_156 vpwr vgnd scs8hd_fill_2
X_101_ _101_/A _144_/A vgnd vpwr scs8hd_buf_1
XFILLER_3_300 vgnd vpwr scs8hd_decap_3
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_19_234 vgnd vpwr scs8hd_decap_8
XFILLER_6_171 vgnd vpwr scs8hd_decap_6
XFILLER_8_10 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_1_.latch/Q mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_96 vpwr vgnd scs8hd_fill_2
XFILLER_17_41 vgnd vpwr scs8hd_decap_4
XFILLER_16_215 vgnd vpwr scs8hd_decap_4
XANTENNA__104__B _110_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _148_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_4.LATCH_2_.latch data_in mem_bottom_ipin_4.LATCH_2_.latch/Q _106_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_4.LATCH_4_.latch/Q mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__205__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_133 vgnd vpwr scs8hd_decap_12
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_255 vgnd vpwr scs8hd_decap_3
XANTENNA__115__A _125_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_284 vpwr vgnd scs8hd_fill_2
XFILLER_5_66 vgnd vpwr scs8hd_fill_1
Xmem_bottom_ipin_6.LATCH_5_.latch data_in mem_bottom_ipin_6.LATCH_5_.latch/Q _125_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_203 vgnd vpwr scs8hd_fill_1
XFILLER_5_236 vgnd vpwr scs8hd_decap_4
XFILLER_5_258 vgnd vpwr scs8hd_fill_1
XFILLER_14_64 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _155_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_239 vgnd vpwr scs8hd_decap_8
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_14_302 vgnd vpwr scs8hd_decap_12
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_63 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_52 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_194_ chanx_right_in[6] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_2_89 vgnd vpwr scs8hd_decap_3
XFILLER_17_184 vgnd vpwr scs8hd_decap_8
XFILLER_17_140 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_32 vpwr vgnd scs8hd_fill_2
XFILLER_11_87 vpwr vgnd scs8hd_fill_2
XFILLER_19_405 vpwr vgnd scs8hd_fill_2
XFILLER_14_143 vgnd vpwr scs8hd_fill_1
XFILLER_14_154 vpwr vgnd scs8hd_fill_2
X_177_ _103_/A _178_/B _177_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_331 vgnd vpwr scs8hd_decap_4
XANTENNA__123__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_191 vpwr vgnd scs8hd_fill_2
X_100_ _125_/A _110_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__208__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_11_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_367 vpwr vgnd scs8hd_fill_2
XFILLER_3_334 vpwr vgnd scs8hd_fill_2
XFILLER_19_279 vgnd vpwr scs8hd_decap_12
XFILLER_19_268 vgnd vpwr scs8hd_decap_4
XFILLER_19_257 vgnd vpwr scs8hd_decap_3
XFILLER_19_202 vgnd vpwr scs8hd_fill_1
XANTENNA__118__A _162_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_2_.latch/Q mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_20 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_3_153 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_7.LATCH_1_.latch data_in mem_bottom_ipin_7.LATCH_1_.latch/Q _137_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_15_293 vpwr vgnd scs8hd_fill_2
XFILLER_0_112 vgnd vpwr scs8hd_fill_1
XFILLER_0_145 vgnd vpwr scs8hd_decap_8
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_0_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_252 vpwr vgnd scs8hd_fill_2
XFILLER_8_267 vgnd vpwr scs8hd_decap_6
XFILLER_8_289 vgnd vpwr scs8hd_decap_8
XANTENNA__115__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _077_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_21 vpwr vgnd scs8hd_fill_2
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__126__A _144_/A vgnd vpwr scs8hd_diode_2
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_14_314 vgnd vpwr scs8hd_fill_1
XPHY_64 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_53 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_42 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_20 vgnd vpwr scs8hd_decap_3
XFILLER_14_358 vpwr vgnd scs8hd_fill_2
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_193_ chanx_right_in[7] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_2_68 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_1_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_362 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_306 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_11 vgnd vpwr scs8hd_decap_4
XFILLER_11_66 vpwr vgnd scs8hd_fill_2
XFILLER_14_100 vgnd vpwr scs8hd_decap_4
XFILLER_14_122 vpwr vgnd scs8hd_fill_2
X_176_ _101_/A _178_/B _176_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__123__B _173_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_398 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_125 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_3.LATCH_4_.latch/Q mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_ipin_0.LATCH_2_.latch/Q mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_3_313 vpwr vgnd scs8hd_fill_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_19_214 vgnd vpwr scs8hd_decap_4
Xmem_top_ipin_0.LATCH_2_.latch data_in mem_top_ipin_0.LATCH_2_.latch/Q _146_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__118__B _115_/B vgnd vpwr scs8hd_diode_2
XFILLER_8_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
X_159_ _159_/A _158_/X _159_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__134__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_180 vgnd vpwr scs8hd_decap_8
XFILLER_18_291 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
XFILLER_3_198 vgnd vpwr scs8hd_decap_4
XFILLER_3_187 vpwr vgnd scs8hd_fill_2
XFILLER_3_176 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _107_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_209 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _188_/HI mem_bottom_ipin_7.LATCH_5_.latch/Q
+ mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_0_102 vpwr vgnd scs8hd_fill_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
XFILLER_5_24 vgnd vpwr scs8hd_decap_4
XFILLER_5_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__131__B _077_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_0.LATCH_2_.latch data_in mem_bottom_ipin_0.LATCH_2_.latch/Q _162_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_367 vpwr vgnd scs8hd_fill_2
XANTENNA__126__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_ipin_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _142_/A vgnd vpwr scs8hd_diode_2
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_14_337 vgnd vpwr scs8hd_decap_6
XPHY_65 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_54 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_43 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_bottom_ipin_2.LATCH_5_.latch data_in mem_bottom_ipin_2.LATCH_5_.latch/Q _175_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_21 vgnd vpwr scs8hd_decap_3
X_192_ chanx_right_in[8] chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_14 vpwr vgnd scs8hd_fill_2
XFILLER_13_381 vgnd vpwr scs8hd_decap_3
XANTENNA__137__A _107_/X vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_2_.latch/Q mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_56 vgnd vpwr scs8hd_decap_3
XFILLER_14_167 vpwr vgnd scs8hd_fill_2
X_175_ _159_/A _178_/B _175_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_20_137 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_0_.latch/Q mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_104 vpwr vgnd scs8hd_fill_2
XFILLER_3_347 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_68 vpwr vgnd scs8hd_fill_2
X_158_ _157_/X _158_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_152 vgnd vpwr scs8hd_fill_1
XFILLER_6_163 vpwr vgnd scs8hd_fill_2
XFILLER_6_196 vgnd vpwr scs8hd_fill_1
XANTENNA__134__B _134_/B vgnd vpwr scs8hd_diode_2
X_089_ _079_/B _089_/B _089_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__150__A _149_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_12_ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_1.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_406 vgnd vpwr scs8hd_fill_1
XFILLER_3_166 vpwr vgnd scs8hd_fill_2
XFILLER_15_240 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__129__B _125_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_1_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_247 vpwr vgnd scs8hd_fill_2
XFILLER_12_298 vgnd vpwr scs8hd_decap_8
XANTENNA__131__C _077_/C vgnd vpwr scs8hd_diode_2
XFILLER_10_6 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_3.LATCH_1_.latch data_in mem_bottom_ipin_3.LATCH_1_.latch/Q _092_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1 mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ bottom_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_14_89 vgnd vpwr scs8hd_fill_1
XFILLER_17_379 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_2.LATCH_4_.latch/Q mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_261 vgnd vpwr scs8hd_fill_1
XFILLER_4_283 vgnd vpwr scs8hd_decap_4
Xmem_bottom_ipin_5.LATCH_4_.latch data_in mem_bottom_ipin_5.LATCH_4_.latch/Q _116_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_209 vgnd vpwr scs8hd_decap_4
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_55 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_44 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_17_176 vpwr vgnd scs8hd_fill_2
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XFILLER_17_198 vpwr vgnd scs8hd_fill_2
XFILLER_13_393 vpwr vgnd scs8hd_fill_2
XANTENNA__137__B _134_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _153_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB _175_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_146 vgnd vpwr scs8hd_decap_6
X_174_ _173_/X _178_/B vgnd vpwr scs8hd_buf_1
XFILLER_6_323 vgnd vpwr scs8hd_decap_6
XFILLER_6_356 vpwr vgnd scs8hd_fill_2
XFILLER_10_363 vpwr vgnd scs8hd_fill_2
XFILLER_10_396 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__148__A _148_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_149 vgnd vpwr scs8hd_decap_6
XFILLER_20_116 vgnd vpwr scs8hd_decap_8
Xmux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _187_/HI mem_bottom_ipin_6.LATCH_5_.latch/Q
+ mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_7_109 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_127 vgnd vpwr scs8hd_fill_1
XFILLER_3_359 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_8_58 vgnd vpwr scs8hd_decap_4
X_157_ _077_/A address[4] address[3] _165_/A _157_/X vgnd vpwr scs8hd_or4_4
XANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_381 vgnd vpwr scs8hd_decap_12
X_088_ _087_/X _089_/B vgnd vpwr scs8hd_buf_1
XANTENNA__150__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_56 vgnd vpwr scs8hd_decap_3
XFILLER_3_101 vpwr vgnd scs8hd_fill_2
XFILLER_15_263 vpwr vgnd scs8hd_fill_2
XANTENNA__145__B _145_/B vgnd vpwr scs8hd_diode_2
X_209_ chanx_left_in[0] chanx_right_out[0] vgnd vpwr scs8hd_buf_2
XANTENNA__161__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_92 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__071__A _159_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_6.LATCH_0_.latch data_in mem_bottom_ipin_6.LATCH_0_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_12_233 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_2_.latch/Q mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_8_226 vpwr vgnd scs8hd_fill_2
XFILLER_12_288 vgnd vpwr scs8hd_fill_1
XFILLER_5_48 vpwr vgnd scs8hd_fill_2
XANTENNA__131__D _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA__156__A _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_292 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_207 vpwr vgnd scs8hd_fill_2
XFILLER_14_68 vpwr vgnd scs8hd_fill_2
Xmux_top_ipin_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_17_358 vpwr vgnd scs8hd_fill_2
XFILLER_17_336 vgnd vpwr scs8hd_decap_12
XFILLER_17_325 vpwr vgnd scs8hd_fill_2
XFILLER_4_240 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_0_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_12 vgnd vpwr scs8hd_decap_3
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_14_328 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_45 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_56 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
Xmux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_17_155 vpwr vgnd scs8hd_fill_2
XFILLER_17_144 vpwr vgnd scs8hd_fill_2
XFILLER_17_100 vpwr vgnd scs8hd_fill_2
XFILLER_9_321 vgnd vpwr scs8hd_decap_3
XFILLER_9_343 vpwr vgnd scs8hd_fill_2
XFILLER_9_376 vpwr vgnd scs8hd_fill_2
XFILLER_11_47 vgnd vpwr scs8hd_decap_3
X_173_ _165_/A _173_/B _173_/X vgnd vpwr scs8hd_or2_4
XFILLER_6_335 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_6
XANTENNA__148__B _145_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_162 vpwr vgnd scs8hd_fill_2
XANTENNA__164__A _148_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_92 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_1_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _154_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__074__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_11_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
X_087_ _084_/A address[2] address[0] _087_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_110 vgnd vpwr scs8hd_decap_4
XFILLER_6_121 vpwr vgnd scs8hd_fill_2
X_156_ _156_/A _156_/Y vgnd vpwr scs8hd_inv_8
XFILLER_12_90 vpwr vgnd scs8hd_fill_2
XFILLER_2_393 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__150__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__159__A _159_/A vgnd vpwr scs8hd_diode_2
XANTENNA__069__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_79 vgnd vpwr scs8hd_decap_6
XFILLER_17_24 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_ipin_1.LATCH_4_.latch/Q mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_297 vgnd vpwr scs8hd_decap_8
XFILLER_15_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__161__B _158_/X vgnd vpwr scs8hd_diode_2
X_139_ address[5] _097_/B _139_/X vgnd vpwr scs8hd_or2_4
X_208_ chanx_left_in[1] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_0_71 vgnd vpwr scs8hd_fill_1
XFILLER_9_80 vpwr vgnd scs8hd_fill_2
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_12_223 vgnd vpwr scs8hd_fill_1
XFILLER_12_267 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_5.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _095_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_260 vpwr vgnd scs8hd_fill_2
XFILLER_14_14 vgnd vpwr scs8hd_decap_4
XFILLER_14_25 vgnd vpwr scs8hd_decap_6
XFILLER_14_36 vgnd vpwr scs8hd_decap_3
XFILLER_5_219 vpwr vgnd scs8hd_fill_2
XANTENNA__082__A _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_403 vgnd vpwr scs8hd_decap_4
XFILLER_17_348 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _186_/HI mem_bottom_ipin_5.LATCH_5_.latch/Q
+ mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_381 vgnd vpwr scs8hd_decap_12
XFILLER_16_370 vpwr vgnd scs8hd_fill_2
XANTENNA__167__A _159_/A vgnd vpwr scs8hd_diode_2
XPHY_35 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_46 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_13 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _077_/A vgnd vpwr scs8hd_diode_2
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_57 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_3 vgnd vpwr scs8hd_decap_3
XFILLER_13_362 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_1.LATCH_4_.latch data_in mem_bottom_ipin_1.LATCH_4_.latch/Q _168_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_104 vgnd vpwr scs8hd_fill_1
XFILLER_14_137 vgnd vpwr scs8hd_decap_6
X_172_ _095_/B _171_/B _172_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_376 vgnd vpwr scs8hd_decap_8
XFILLER_10_398 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_181 vpwr vgnd scs8hd_fill_2
XANTENNA__164__B _158_/X vgnd vpwr scs8hd_diode_2
XANTENNA__180__A _095_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_2_.latch/Q mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_3_317 vpwr vgnd scs8hd_fill_2
XFILLER_15_402 vgnd vpwr scs8hd_decap_4
XFILLER_8_27 vpwr vgnd scs8hd_fill_2
X_086_ _079_/B _103_/A _086_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_155_ _155_/A _155_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_144 vgnd vpwr scs8hd_decap_8
XFILLER_6_188 vpwr vgnd scs8hd_fill_2
XFILLER_10_173 vgnd vpwr scs8hd_decap_4
XFILLER_18_295 vgnd vpwr scs8hd_decap_12
XFILLER_18_273 vpwr vgnd scs8hd_fill_2
XANTENNA__159__B _158_/X vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_2.LATCH_0_.latch data_in _156_/A _152_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__175__A _159_/A vgnd vpwr scs8hd_diode_2
XANTENNA__069__B _067_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__085__A _084_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_136 vpwr vgnd scs8hd_fill_2
X_207_ chanx_left_in[2] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_15_276 vpwr vgnd scs8hd_fill_2
X_069_ address[1] _067_/Y _069_/C _069_/X vgnd vpwr scs8hd_or3_4
X_138_ _148_/A _134_/B _138_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_94 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_106 vgnd vpwr scs8hd_decap_6
XFILLER_8_206 vpwr vgnd scs8hd_fill_2
XFILLER_12_279 vgnd vpwr scs8hd_decap_3
XFILLER_5_39 vpwr vgnd scs8hd_fill_2
XANTENNA__172__B _171_/B vgnd vpwr scs8hd_diode_2
XANTENNA__082__B _101_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_ipin_2.LATCH_0_.latch data_in mem_bottom_ipin_2.LATCH_0_.latch/Q _180_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_264 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_3.LATCH_1_.latch/Q mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_393 vgnd vpwr scs8hd_decap_4
XANTENNA__167__B _171_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_60 vpwr vgnd scs8hd_fill_2
XFILLER_6_93 vpwr vgnd scs8hd_fill_2
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_69 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_58 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_47 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _077_/B vgnd vpwr scs8hd_diode_2
XPHY_25 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__093__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
XFILLER_2_18 vgnd vpwr scs8hd_decap_12
Xmem_bottom_ipin_4.LATCH_3_.latch data_in mem_bottom_ipin_4.LATCH_3_.latch/Q _104_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_301 vpwr vgnd scs8hd_fill_2
XANTENNA__178__A _089_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_ipin_0.LATCH_4_.latch/Q mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__088__A _087_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_171_ _107_/A _171_/B _171_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_337 vpwr vgnd scs8hd_fill_2
XFILLER_10_311 vpwr vgnd scs8hd_fill_2
XFILLER_10_388 vgnd vpwr scs8hd_decap_8
XFILLER_13_193 vgnd vpwr scs8hd_decap_4
XFILLER_9_142 vgnd vpwr scs8hd_decap_3
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XANTENNA__180__B _178_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_370 vgnd vpwr scs8hd_decap_8
XFILLER_5_381 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_7.LATCH_2_.latch/Q mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_108 vpwr vgnd scs8hd_fill_2
XANTENNA__090__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_085_ _084_/X _103_/A vgnd vpwr scs8hd_buf_1
X_154_ _154_/A _154_/Y vgnd vpwr scs8hd_inv_8
XFILLER_6_167 vpwr vgnd scs8hd_fill_2
XFILLER_18_241 vgnd vpwr scs8hd_decap_12
XFILLER_18_230 vgnd vpwr scs8hd_decap_8
XANTENNA__175__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA__069__C _069_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_17_48 vgnd vpwr scs8hd_decap_8
XFILLER_17_37 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _185_/HI mem_bottom_ipin_4.LATCH_5_.latch/Q
+ mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_406 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_137_ _107_/X _134_/B _137_/Y vgnd vpwr scs8hd_nor2_4
X_206_ chanx_left_in[3] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_192 vgnd vpwr scs8hd_decap_3
X_068_ address[0] _069_/C vgnd vpwr scs8hd_inv_8
XFILLER_17_3 vpwr vgnd scs8hd_fill_2
XFILLER_0_129 vpwr vgnd scs8hd_fill_2
XANTENNA__096__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_20_280 vgnd vpwr scs8hd_decap_12
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
XFILLER_17_306 vgnd vpwr scs8hd_decap_12
XFILLER_4_276 vgnd vpwr scs8hd_decap_4
XFILLER_4_287 vgnd vpwr scs8hd_fill_1
Xmux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_2_.latch/Q mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_6_83 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_7.LATCH_2_.latch data_in mem_bottom_ipin_7.LATCH_2_.latch/Q _136_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_59 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_48 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_15 vgnd vpwr scs8hd_decap_3
XANTENNA__077__C _077_/C vgnd vpwr scs8hd_diode_2
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB _178_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_136 vgnd vpwr scs8hd_decap_4
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_397 vgnd vpwr scs8hd_decap_8
XFILLER_13_342 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__178__B _178_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__194__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_11_28 vpwr vgnd scs8hd_fill_2
X_170_ _089_/B _171_/B _170_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_305 vgnd vpwr scs8hd_decap_3
XFILLER_13_172 vgnd vpwr scs8hd_decap_3
XFILLER_9_187 vpwr vgnd scs8hd_fill_2
XFILLER_3_73 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vpwr vgnd scs8hd_fill_2
XANTENNA__090__C _069_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__099__A _098_/X vgnd vpwr scs8hd_diode_2
X_153_ _153_/A _153_/Y vgnd vpwr scs8hd_inv_8
XFILLER_10_120 vgnd vpwr scs8hd_decap_4
X_084_ _084_/A address[2] _069_/C _084_/X vgnd vpwr scs8hd_or3_4
XFILLER_2_341 vpwr vgnd scs8hd_fill_2
XFILLER_12_82 vgnd vpwr scs8hd_decap_8
XFILLER_12_93 vpwr vgnd scs8hd_fill_2
XFILLER_18_253 vgnd vpwr scs8hd_decap_3
XFILLER_3_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_2.LATCH_1_.latch/Q mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_245 vpwr vgnd scs8hd_fill_2
XFILLER_15_223 vpwr vgnd scs8hd_fill_2
X_205_ chanx_left_in[4] chanx_right_out[4] vgnd vpwr scs8hd_buf_2
X_136_ _162_/A _134_/B _136_/Y vgnd vpwr scs8hd_nor2_4
X_067_ address[2] _067_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_63 vgnd vpwr scs8hd_decap_8
XFILLER_0_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_215 vpwr vgnd scs8hd_fill_2
XFILLER_20_292 vgnd vpwr scs8hd_decap_12
XFILLER_12_248 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_ipin_0.INVTX1_2_.scs8hd_inv_1 chanx_left_in[7] mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_7_296 vpwr vgnd scs8hd_fill_2
X_119_ _107_/X _115_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_381 vgnd vpwr scs8hd_decap_12
XANTENNA__197__A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmem_top_ipin_0.LATCH_3_.latch data_in mem_top_ipin_0.LATCH_3_.latch/Q _145_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_329 vgnd vpwr scs8hd_decap_4
XFILLER_17_318 vgnd vpwr scs8hd_decap_4
XFILLER_4_222 vgnd vpwr scs8hd_decap_4
XFILLER_4_233 vgnd vpwr scs8hd_decap_4
XFILLER_4_244 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_6.LATCH_2_.latch/Q mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _153_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_16 vgnd vpwr scs8hd_decap_3
XANTENNA__077__D _165_/A vgnd vpwr scs8hd_diode_2
XANTENNA__093__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_1_269 vgnd vpwr scs8hd_decap_12
XFILLER_17_159 vpwr vgnd scs8hd_fill_2
XFILLER_17_148 vgnd vpwr scs8hd_decap_4
XFILLER_17_104 vgnd vpwr scs8hd_fill_1
XFILLER_15_60 vgnd vpwr scs8hd_fill_1
XFILLER_13_376 vgnd vpwr scs8hd_decap_3
XFILLER_9_358 vpwr vgnd scs8hd_fill_2
XFILLER_0_280 vgnd vpwr scs8hd_decap_12
Xmux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _184_/HI mem_bottom_ipin_3.LATCH_5_.latch/Q
+ mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_14_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_13_140 vpwr vgnd scs8hd_fill_2
Xmem_bottom_ipin_0.LATCH_3_.latch data_in mem_bottom_ipin_0.LATCH_3_.latch/Q _161_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_361 vgnd vpwr scs8hd_fill_1
XFILLER_3_309 vpwr vgnd scs8hd_fill_2
X_152_ _173_/B _149_/B address[0] _152_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_125 vpwr vgnd scs8hd_fill_2
XFILLER_10_154 vpwr vgnd scs8hd_fill_2
X_083_ address[1] _084_/A vgnd vpwr scs8hd_inv_8
XFILLER_18_265 vgnd vpwr scs8hd_decap_8
X_204_ chanx_left_in[5] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_135_ _145_/A _134_/B _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_150 vgnd vpwr scs8hd_decap_3
XFILLER_0_86 vgnd vpwr scs8hd_decap_6
XFILLER_9_62 vgnd vpwr scs8hd_decap_3
XFILLER_9_84 vpwr vgnd scs8hd_fill_2
XFILLER_18_93 vgnd vpwr scs8hd_decap_8
XFILLER_11_293 vpwr vgnd scs8hd_fill_2
XFILLER_7_275 vpwr vgnd scs8hd_fill_2
X_118_ _162_/A _115_/B _118_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_393 vgnd vpwr scs8hd_decap_12
XFILLER_14_18 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_94 vgnd vpwr scs8hd_decap_12
XFILLER_16_374 vpwr vgnd scs8hd_fill_2
XFILLER_16_341 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_15_83 vpwr vgnd scs8hd_fill_2
XFILLER_13_355 vgnd vpwr scs8hd_decap_4
XFILLER_9_315 vgnd vpwr scs8hd_decap_4
XFILLER_9_337 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_0_292 vpwr vgnd scs8hd_fill_2
XFILLER_16_193 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_1.LATCH_1_.latch/Q mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_358 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_3.LATCH_2_.latch data_in mem_bottom_ipin_3.LATCH_2_.latch/Q _089_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1 mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A
+ top_grid_pin_4_ vgnd vpwr scs8hd_inv_1
XFILLER_9_101 vpwr vgnd scs8hd_fill_2
XFILLER_9_134 vpwr vgnd scs8hd_fill_2
XFILLER_9_156 vgnd vpwr scs8hd_decap_4
XFILLER_3_97 vpwr vgnd scs8hd_fill_2
XFILLER_3_53 vpwr vgnd scs8hd_fill_2
XFILLER_3_42 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_ipin_5.LATCH_5_.latch data_in mem_bottom_ipin_5.LATCH_5_.latch/Q _115_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_406 vgnd vpwr scs8hd_fill_1
X_151_ _173_/B _149_/B _069_/C _151_/Y vgnd vpwr scs8hd_nor3_4
X_082_ _079_/B _101_/A _082_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_188 vgnd vpwr scs8hd_decap_3
XFILLER_2_398 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_6.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_SLEEPB _082_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_5.LATCH_2_.latch/Q mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_236 vpwr vgnd scs8hd_fill_2
X_203_ chanx_left_in[6] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
X_134_ _144_/A _134_/B _134_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_184 vgnd vpwr scs8hd_decap_8
XFILLER_2_173 vgnd vpwr scs8hd_decap_8
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_98 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_206 vgnd vpwr scs8hd_decap_8
XFILLER_20_261 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_ipin_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _183_/HI mem_bottom_ipin_2.LATCH_5_.latch/Q
+ mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_7_210 vpwr vgnd scs8hd_fill_2
XFILLER_7_254 vgnd vpwr scs8hd_decap_4
X_117_ _145_/A _115_/B _117_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_350 vgnd vpwr scs8hd_decap_12
XFILLER_4_202 vgnd vpwr scs8hd_fill_1
XFILLER_4_257 vgnd vpwr scs8hd_decap_4
XFILLER_4_268 vgnd vpwr scs8hd_decap_6
XFILLER_16_353 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_64 vgnd vpwr scs8hd_decap_4
XFILLER_19_180 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_9_8 vpwr vgnd scs8hd_fill_2
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_150 vgnd vpwr scs8hd_decap_3
Xmem_bottom_ipin_6.LATCH_1_.latch data_in mem_bottom_ipin_6.LATCH_1_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_6_319 vpwr vgnd scs8hd_fill_2
XFILLER_10_315 vpwr vgnd scs8hd_fill_2
XFILLER_10_337 vgnd vpwr scs8hd_decap_8
XFILLER_13_153 vpwr vgnd scs8hd_fill_2
XFILLER_5_341 vgnd vpwr scs8hd_decap_4
XFILLER_5_385 vpwr vgnd scs8hd_fill_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_150_ _149_/A _149_/B address[0] _150_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_138 vgnd vpwr scs8hd_decap_4
X_081_ _080_/X _101_/A vgnd vpwr scs8hd_buf_1
XFILLER_12_41 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_193 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB _146_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_259 vpwr vgnd scs8hd_fill_2
XFILLER_15_204 vpwr vgnd scs8hd_fill_2
XANTENNA__200__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_202_ chanx_left_in[7] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
X_133_ _125_/A _134_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_403 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_163 vgnd vpwr scs8hd_decap_6
XFILLER_2_130 vpwr vgnd scs8hd_fill_2
XFILLER_17_7 vpwr vgnd scs8hd_fill_2
XFILLER_0_44 vgnd vpwr scs8hd_decap_12
XANTENNA__110__A _148_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_42 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_9_97 vpwr vgnd scs8hd_fill_2
XFILLER_20_273 vgnd vpwr scs8hd_decap_6
XFILLER_4_406 vgnd vpwr scs8hd_fill_1
XFILLER_18_62 vgnd vpwr scs8hd_decap_8
XFILLER_18_84 vgnd vpwr scs8hd_decap_8
XFILLER_18_73 vgnd vpwr scs8hd_decap_8
XANTENNA__105__A _089_/B vgnd vpwr scs8hd_diode_2
X_116_ _144_/A _115_/B _116_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _154_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_362 vgnd vpwr scs8hd_decap_4
Xmux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_ipin_0.LATCH_1_.latch/Q mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_63 vgnd vpwr scs8hd_decap_12
XFILLER_16_398 vgnd vpwr scs8hd_decap_8
XFILLER_6_21 vpwr vgnd scs8hd_fill_2
XFILLER_6_43 vgnd vpwr scs8hd_decap_3
XFILLER_6_87 vgnd vpwr scs8hd_decap_3
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XANTENNA__102__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_261 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_350 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_ipin_4.LATCH_2_.latch/Q mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__203__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_110 vpwr vgnd scs8hd_fill_2
XFILLER_3_22 vgnd vpwr scs8hd_decap_4
XFILLER_3_11 vpwr vgnd scs8hd_fill_2
XFILLER_5_364 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_77 vpwr vgnd scs8hd_fill_2
XFILLER_3_33 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_191 vpwr vgnd scs8hd_fill_2
Xmux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _182_/HI mem_bottom_ipin_1.LATCH_5_.latch/Q
+ mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_080_ address[1] _067_/Y address[0] _080_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_106 vpwr vgnd scs8hd_fill_2
XFILLER_10_124 vgnd vpwr scs8hd_fill_1
XFILLER_2_345 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_18_279 vgnd vpwr scs8hd_decap_12
XANTENNA__108__A _107_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_150 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_249 vgnd vpwr scs8hd_fill_1
XFILLER_15_227 vpwr vgnd scs8hd_fill_2
X_201_ chanx_left_in[8] chanx_right_out[8] vgnd vpwr scs8hd_buf_2
X_132_ _131_/X _134_/B vgnd vpwr scs8hd_buf_1
Xmem_bottom_ipin_1.LATCH_5_.latch data_in mem_bottom_ipin_1.LATCH_5_.latch/Q _167_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_197 vgnd vpwr scs8hd_decap_12
XFILLER_2_142 vgnd vpwr scs8hd_decap_8
XFILLER_0_56 vgnd vpwr scs8hd_decap_6
XANTENNA__110__B _110_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_271 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_4.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_219 vpwr vgnd scs8hd_fill_2
XFILLER_18_30 vgnd vpwr scs8hd_fill_1
XFILLER_7_223 vpwr vgnd scs8hd_fill_2
XFILLER_11_274 vpwr vgnd scs8hd_fill_2
X_115_ _125_/A _115_/B _115_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__121__A _121_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_top_ipin_2.LATCH_1_.latch data_in _155_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_7.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vgnd vpwr scs8hd_decap_4
XFILLER_4_226 vgnd vpwr scs8hd_fill_1
XANTENNA__206__A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_20_75 vgnd vpwr scs8hd_decap_12
XANTENNA__116__A _144_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_6_55 vgnd vpwr scs8hd_decap_3
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_13_336 vgnd vpwr scs8hd_decap_4
XFILLER_0_273 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_ipin_2.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_16_163 vpwr vgnd scs8hd_fill_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_384 vpwr vgnd scs8hd_fill_2
XFILLER_12_391 vgnd vpwr scs8hd_decap_6
.ends

