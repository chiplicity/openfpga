magic
tech sky130A
magscale 1 2
timestamp 1604667884
<< viali >>
rect 23949 19087 23983 19121
rect 24501 19087 24535 19121
rect 24133 18951 24167 18985
rect 16681 18747 16715 18781
rect 20637 18747 20671 18781
rect 8852 18679 8886 18713
rect 8585 18611 8619 18645
rect 15557 18611 15591 18645
rect 20453 18611 20487 18645
rect 23949 18611 23983 18645
rect 25053 18611 25087 18645
rect 15301 18543 15335 18577
rect 9965 18407 9999 18441
rect 24133 18407 24167 18441
rect 25237 18407 25271 18441
rect 8677 18203 8711 18237
rect 15485 18203 15519 18237
rect 25053 18203 25087 18237
rect 8953 18135 8987 18169
rect 23765 18135 23799 18169
rect 23949 17999 23983 18033
rect 24501 17999 24535 18033
rect 15853 17931 15887 17965
rect 20453 17863 20487 17897
rect 24133 17863 24167 17897
rect 23949 17523 23983 17557
rect 24133 17319 24167 17353
rect 18061 17115 18095 17149
rect 24041 17115 24075 17149
rect 17969 16979 18003 17013
rect 18705 16979 18739 17013
rect 18521 16843 18555 16877
rect 17509 16775 17543 16809
rect 18429 16775 18463 16809
rect 14381 16571 14415 16605
rect 18337 16571 18371 16605
rect 13001 16435 13035 16469
rect 13268 16435 13302 16469
rect 7021 16027 7055 16061
rect 13001 16027 13035 16061
rect 24501 16027 24535 16061
rect 7113 15891 7147 15925
rect 23949 15823 23983 15857
rect 7358 15755 7392 15789
rect 8493 15687 8527 15721
rect 13461 15687 13495 15721
rect 24133 15687 24167 15721
rect 7205 15483 7239 15517
rect 23949 15347 23983 15381
rect 18613 15143 18647 15177
rect 24133 15143 24167 15177
rect 18521 14939 18555 14973
rect 24041 14939 24075 14973
rect 18337 14803 18371 14837
rect 19073 14803 19107 14837
rect 18889 14667 18923 14701
rect 18981 14599 19015 14633
rect 18613 14395 18647 14429
rect 19441 14395 19475 14429
rect 19809 14259 19843 14293
rect 19901 14191 19935 14225
rect 20085 14191 20119 14225
rect 19625 13647 19659 13681
rect 19901 13647 19935 13681
rect 19073 13511 19107 13545
rect 20361 13511 20395 13545
rect 13553 13307 13587 13341
rect 20085 13307 20119 13341
rect 1409 13171 1443 13205
rect 13921 13171 13955 13205
rect 20177 13171 20211 13205
rect 14013 13103 14047 13137
rect 14197 13103 14231 13137
rect 20361 13103 20395 13137
rect 19717 13035 19751 13069
rect 1593 12967 1627 13001
rect 13093 12967 13127 13001
rect 14197 12763 14231 12797
rect 20085 12763 20119 12797
rect 13093 12695 13127 12729
rect 13737 12627 13771 12661
rect 1409 12559 1443 12593
rect 1961 12559 1995 12593
rect 12909 12559 12943 12593
rect 13461 12559 13495 12593
rect 13553 12491 13587 12525
rect 1593 12423 1627 12457
rect 19717 12423 19751 12457
rect 20453 12423 20487 12457
rect 1593 12219 1627 12253
rect 13921 12219 13955 12253
rect 13185 12151 13219 12185
rect 8309 12083 8343 12117
rect 8401 12015 8435 12049
rect 8585 12015 8619 12049
rect 7941 11947 7975 11981
rect 13645 11947 13679 11981
rect 12081 11879 12115 11913
rect 8033 11675 8067 11709
rect 11897 11675 11931 11709
rect 12081 11675 12115 11709
rect 24133 11607 24167 11641
rect 12633 11539 12667 11573
rect 1409 11471 1443 11505
rect 1961 11471 1995 11505
rect 23949 11471 23983 11505
rect 24501 11471 24535 11505
rect 12449 11403 12483 11437
rect 1593 11335 1627 11369
rect 8309 11335 8343 11369
rect 8677 11335 8711 11369
rect 12541 11335 12575 11369
rect 7757 11131 7791 11165
rect 12081 11131 12115 11165
rect 1409 10995 1443 11029
rect 8125 10995 8159 11029
rect 23949 10995 23983 11029
rect 8217 10927 8251 10961
rect 8401 10927 8435 10961
rect 1593 10859 1627 10893
rect 24133 10859 24167 10893
rect 2053 10587 2087 10621
rect 2421 10587 2455 10621
rect 7941 10587 7975 10621
rect 8953 10587 8987 10621
rect 24041 10587 24075 10621
rect 7113 10519 7147 10553
rect 8585 10451 8619 10485
rect 1409 10383 1443 10417
rect 8309 10315 8343 10349
rect 1593 10247 1627 10281
rect 7389 10247 7423 10281
rect 7849 10247 7883 10281
rect 8401 10247 8435 10281
rect 8033 10043 8067 10077
rect 8401 10043 8435 10077
rect 1409 9907 1443 9941
rect 1593 9703 1627 9737
rect 2053 9499 2087 9533
rect 2421 9431 2455 9465
rect 1409 9295 1443 9329
rect 23949 9295 23983 9329
rect 24501 9295 24535 9329
rect 1593 9159 1627 9193
rect 24133 9159 24167 9193
rect 1409 8819 1443 8853
rect 23949 8819 23983 8853
rect 1593 8615 1627 8649
rect 24133 8615 24167 8649
rect 1593 8411 1627 8445
rect 23857 8411 23891 8445
rect 24133 8343 24167 8377
rect 23949 8207 23983 8241
rect 24501 8207 24535 8241
rect 24133 7867 24167 7901
rect 23949 7731 23983 7765
rect 22661 7323 22695 7357
rect 23121 7323 23155 7357
rect 18889 7255 18923 7289
rect 18705 7119 18739 7153
rect 19257 7119 19291 7153
rect 22477 7119 22511 7153
rect 23949 7119 23983 7153
rect 10885 6643 10919 6677
rect 14657 6643 14691 6677
rect 23949 6643 23983 6677
rect 24133 6507 24167 6541
rect 11069 6439 11103 6473
rect 14841 6439 14875 6473
rect 10885 6235 10919 6269
rect 14657 6235 14691 6269
rect 23949 6235 23983 6269
rect 12817 5691 12851 5725
rect 4813 5555 4847 5589
rect 12633 5555 12667 5589
rect 4997 5419 5031 5453
rect 4813 5147 4847 5181
rect 12633 5147 12667 5181
rect 13921 5147 13955 5181
rect 13737 4943 13771 4977
rect 14289 4943 14323 4977
rect 23949 4943 23983 4977
rect 24501 4943 24535 4977
rect 24133 4807 24167 4841
rect 16313 4467 16347 4501
rect 20729 4467 20763 4501
rect 16497 4331 16531 4365
rect 20913 4331 20947 4365
rect 21097 4059 21131 4093
rect 16405 3991 16439 4025
rect 21465 3855 21499 3889
rect 23949 3855 23983 3889
rect 24501 3855 24535 3889
rect 21649 3719 21683 3753
rect 22109 3719 22143 3753
rect 24133 3719 24167 3753
rect 23949 3379 23983 3413
rect 24133 3243 24167 3277
rect 23857 2971 23891 3005
rect 1409 2767 1443 2801
rect 1961 2767 1995 2801
rect 23949 2767 23983 2801
rect 24501 2767 24535 2801
rect 1593 2631 1627 2665
rect 24133 2631 24167 2665
rect 24225 2427 24259 2461
rect 1409 2291 1443 2325
rect 2053 2291 2087 2325
rect 24041 2291 24075 2325
rect 24593 2291 24627 2325
rect 25145 2291 25179 2325
rect 25697 2291 25731 2325
rect 1593 2087 1627 2121
rect 25329 2087 25363 2121
<< metal1 >>
rect 1104 21612 28888 21634
rect 1104 21560 5982 21612
rect 6034 21560 6046 21612
rect 6098 21560 6110 21612
rect 6162 21560 6174 21612
rect 6226 21560 15982 21612
rect 16034 21560 16046 21612
rect 16098 21560 16110 21612
rect 16162 21560 16174 21612
rect 16226 21560 25982 21612
rect 26034 21560 26046 21612
rect 26098 21560 26110 21612
rect 26162 21560 26174 21612
rect 26226 21560 28888 21612
rect 1104 21538 28888 21560
rect 1104 21068 28888 21090
rect 1104 21016 10982 21068
rect 11034 21016 11046 21068
rect 11098 21016 11110 21068
rect 11162 21016 11174 21068
rect 11226 21016 20982 21068
rect 21034 21016 21046 21068
rect 21098 21016 21110 21068
rect 21162 21016 21174 21068
rect 21226 21016 28888 21068
rect 1104 20994 28888 21016
rect 3418 20574 3424 20626
rect 3476 20614 3482 20626
rect 19794 20614 19800 20626
rect 3476 20586 19800 20614
rect 3476 20574 3482 20586
rect 19794 20574 19800 20586
rect 19852 20574 19858 20626
rect 20162 20574 20168 20626
rect 20220 20614 20226 20626
rect 24854 20614 24860 20626
rect 20220 20586 24860 20614
rect 20220 20574 20226 20586
rect 24854 20574 24860 20586
rect 24912 20574 24918 20626
rect 1104 20524 28888 20546
rect 1104 20472 5982 20524
rect 6034 20472 6046 20524
rect 6098 20472 6110 20524
rect 6162 20472 6174 20524
rect 6226 20472 15982 20524
rect 16034 20472 16046 20524
rect 16098 20472 16110 20524
rect 16162 20472 16174 20524
rect 16226 20472 25982 20524
rect 26034 20472 26046 20524
rect 26098 20472 26110 20524
rect 26162 20472 26174 20524
rect 26226 20472 28888 20524
rect 1104 20450 28888 20472
rect 1104 19980 28888 20002
rect 1104 19928 10982 19980
rect 11034 19928 11046 19980
rect 11098 19928 11110 19980
rect 11162 19928 11174 19980
rect 11226 19928 20982 19980
rect 21034 19928 21046 19980
rect 21098 19928 21110 19980
rect 21162 19928 21174 19980
rect 21226 19928 28888 19980
rect 1104 19906 28888 19928
rect 1104 19436 28888 19458
rect 1104 19384 5982 19436
rect 6034 19384 6046 19436
rect 6098 19384 6110 19436
rect 6162 19384 6174 19436
rect 6226 19384 15982 19436
rect 16034 19384 16046 19436
rect 16098 19384 16110 19436
rect 16162 19384 16174 19436
rect 16226 19384 25982 19436
rect 26034 19384 26046 19436
rect 26098 19384 26110 19436
rect 26162 19384 26174 19436
rect 26226 19384 28888 19436
rect 1104 19362 28888 19384
rect 23934 19118 23940 19130
rect 23895 19090 23940 19118
rect 23934 19078 23940 19090
rect 23992 19118 23998 19130
rect 24489 19121 24547 19127
rect 24489 19118 24501 19121
rect 23992 19090 24501 19118
rect 23992 19078 23998 19090
rect 24489 19087 24501 19090
rect 24535 19087 24547 19121
rect 24489 19081 24547 19087
rect 24121 18985 24179 18991
rect 24121 18951 24133 18985
rect 24167 18982 24179 18985
rect 24670 18982 24676 18994
rect 24167 18954 24676 18982
rect 24167 18951 24179 18954
rect 24121 18945 24179 18951
rect 24670 18942 24676 18954
rect 24728 18942 24734 18994
rect 1104 18892 28888 18914
rect 1104 18840 10982 18892
rect 11034 18840 11046 18892
rect 11098 18840 11110 18892
rect 11162 18840 11174 18892
rect 11226 18840 20982 18892
rect 21034 18840 21046 18892
rect 21098 18840 21110 18892
rect 21162 18840 21174 18892
rect 21226 18840 28888 18892
rect 1104 18818 28888 18840
rect 16666 18778 16672 18790
rect 16627 18750 16672 18778
rect 16666 18738 16672 18750
rect 16724 18738 16730 18790
rect 20622 18778 20628 18790
rect 20583 18750 20628 18778
rect 20622 18738 20628 18750
rect 20680 18738 20686 18790
rect 8846 18719 8852 18722
rect 8840 18710 8852 18719
rect 8807 18682 8852 18710
rect 8840 18673 8852 18682
rect 8846 18670 8852 18673
rect 8904 18670 8910 18722
rect 8570 18642 8576 18654
rect 8531 18614 8576 18642
rect 8570 18602 8576 18614
rect 8628 18602 8634 18654
rect 15194 18602 15200 18654
rect 15252 18642 15258 18654
rect 15545 18645 15603 18651
rect 15545 18642 15557 18645
rect 15252 18614 15557 18642
rect 15252 18602 15258 18614
rect 15545 18611 15557 18614
rect 15591 18611 15603 18645
rect 20438 18642 20444 18654
rect 20399 18614 20444 18642
rect 15545 18605 15603 18611
rect 20438 18602 20444 18614
rect 20496 18602 20502 18654
rect 23750 18602 23756 18654
rect 23808 18642 23814 18654
rect 23937 18645 23995 18651
rect 23937 18642 23949 18645
rect 23808 18614 23949 18642
rect 23808 18602 23814 18614
rect 23937 18611 23949 18614
rect 23983 18611 23995 18645
rect 25038 18642 25044 18654
rect 24999 18614 25044 18642
rect 23937 18605 23995 18611
rect 25038 18602 25044 18614
rect 25096 18602 25102 18654
rect 15286 18574 15292 18586
rect 15247 18546 15292 18574
rect 15286 18534 15292 18546
rect 15344 18534 15350 18586
rect 9950 18438 9956 18450
rect 9911 18410 9956 18438
rect 9950 18398 9956 18410
rect 10008 18398 10014 18450
rect 24118 18438 24124 18450
rect 24079 18410 24124 18438
rect 24118 18398 24124 18410
rect 24176 18398 24182 18450
rect 25225 18441 25283 18447
rect 25225 18407 25237 18441
rect 25271 18438 25283 18441
rect 25314 18438 25320 18450
rect 25271 18410 25320 18438
rect 25271 18407 25283 18410
rect 25225 18401 25283 18407
rect 25314 18398 25320 18410
rect 25372 18398 25378 18450
rect 1104 18348 28888 18370
rect 1104 18296 5982 18348
rect 6034 18296 6046 18348
rect 6098 18296 6110 18348
rect 6162 18296 6174 18348
rect 6226 18296 15982 18348
rect 16034 18296 16046 18348
rect 16098 18296 16110 18348
rect 16162 18296 16174 18348
rect 16226 18296 25982 18348
rect 26034 18296 26046 18348
rect 26098 18296 26110 18348
rect 26162 18296 26174 18348
rect 26226 18296 28888 18348
rect 1104 18274 28888 18296
rect 8665 18237 8723 18243
rect 8665 18203 8677 18237
rect 8711 18234 8723 18237
rect 8846 18234 8852 18246
rect 8711 18206 8852 18234
rect 8711 18203 8723 18206
rect 8665 18197 8723 18203
rect 8846 18194 8852 18206
rect 8904 18194 8910 18246
rect 15286 18194 15292 18246
rect 15344 18234 15350 18246
rect 15473 18237 15531 18243
rect 15473 18234 15485 18237
rect 15344 18206 15485 18234
rect 15344 18194 15350 18206
rect 15473 18203 15485 18206
rect 15519 18203 15531 18237
rect 25038 18234 25044 18246
rect 24999 18206 25044 18234
rect 15473 18197 15531 18203
rect 25038 18194 25044 18206
rect 25096 18194 25102 18246
rect 8570 18126 8576 18178
rect 8628 18166 8634 18178
rect 8941 18169 8999 18175
rect 8941 18166 8953 18169
rect 8628 18138 8953 18166
rect 8628 18126 8634 18138
rect 8941 18135 8953 18138
rect 8987 18135 8999 18169
rect 23750 18166 23756 18178
rect 23711 18138 23756 18166
rect 8941 18129 8999 18135
rect 23750 18126 23756 18138
rect 23808 18126 23814 18178
rect 23934 18030 23940 18042
rect 23895 18002 23940 18030
rect 23934 17990 23940 18002
rect 23992 18030 23998 18042
rect 24489 18033 24547 18039
rect 24489 18030 24501 18033
rect 23992 18002 24501 18030
rect 23992 17990 23998 18002
rect 24489 17999 24501 18002
rect 24535 17999 24547 18033
rect 24489 17993 24547 17999
rect 15194 17922 15200 17974
rect 15252 17962 15258 17974
rect 15841 17965 15899 17971
rect 15841 17962 15853 17965
rect 15252 17934 15853 17962
rect 15252 17922 15258 17934
rect 15841 17931 15853 17934
rect 15887 17931 15899 17965
rect 15841 17925 15899 17931
rect 19334 17854 19340 17906
rect 19392 17894 19398 17906
rect 20438 17894 20444 17906
rect 19392 17866 20444 17894
rect 19392 17854 19398 17866
rect 20438 17854 20444 17866
rect 20496 17854 20502 17906
rect 24121 17897 24179 17903
rect 24121 17863 24133 17897
rect 24167 17894 24179 17897
rect 24210 17894 24216 17906
rect 24167 17866 24216 17894
rect 24167 17863 24179 17866
rect 24121 17857 24179 17863
rect 24210 17854 24216 17866
rect 24268 17854 24274 17906
rect 1104 17804 28888 17826
rect 1104 17752 10982 17804
rect 11034 17752 11046 17804
rect 11098 17752 11110 17804
rect 11162 17752 11174 17804
rect 11226 17752 20982 17804
rect 21034 17752 21046 17804
rect 21098 17752 21110 17804
rect 21162 17752 21174 17804
rect 21226 17752 28888 17804
rect 1104 17730 28888 17752
rect 23937 17557 23995 17563
rect 23937 17523 23949 17557
rect 23983 17554 23995 17557
rect 24302 17554 24308 17566
rect 23983 17526 24308 17554
rect 23983 17523 23995 17526
rect 23937 17517 23995 17523
rect 24302 17514 24308 17526
rect 24360 17514 24366 17566
rect 23474 17310 23480 17362
rect 23532 17350 23538 17362
rect 24121 17353 24179 17359
rect 24121 17350 24133 17353
rect 23532 17322 24133 17350
rect 23532 17310 23538 17322
rect 24121 17319 24133 17322
rect 24167 17319 24179 17353
rect 24121 17313 24179 17319
rect 1104 17260 28888 17282
rect 1104 17208 5982 17260
rect 6034 17208 6046 17260
rect 6098 17208 6110 17260
rect 6162 17208 6174 17260
rect 6226 17208 15982 17260
rect 16034 17208 16046 17260
rect 16098 17208 16110 17260
rect 16162 17208 16174 17260
rect 16226 17208 25982 17260
rect 26034 17208 26046 17260
rect 26098 17208 26110 17260
rect 26162 17208 26174 17260
rect 26226 17208 28888 17260
rect 1104 17186 28888 17208
rect 18049 17149 18107 17155
rect 18049 17115 18061 17149
rect 18095 17146 18107 17149
rect 19242 17146 19248 17158
rect 18095 17118 19248 17146
rect 18095 17115 18107 17118
rect 18049 17109 18107 17115
rect 19242 17106 19248 17118
rect 19300 17106 19306 17158
rect 24029 17149 24087 17155
rect 24029 17115 24041 17149
rect 24075 17146 24087 17149
rect 24302 17146 24308 17158
rect 24075 17118 24308 17146
rect 24075 17115 24087 17118
rect 24029 17109 24087 17115
rect 24302 17106 24308 17118
rect 24360 17106 24366 17158
rect 17957 17013 18015 17019
rect 17957 16979 17969 17013
rect 18003 17010 18015 17013
rect 18690 17010 18696 17022
rect 18003 16982 18696 17010
rect 18003 16979 18015 16982
rect 17957 16973 18015 16979
rect 18690 16970 18696 16982
rect 18748 16970 18754 17022
rect 18509 16877 18567 16883
rect 18509 16874 18521 16877
rect 17512 16846 18521 16874
rect 17512 16818 17540 16846
rect 18509 16843 18521 16846
rect 18555 16843 18567 16877
rect 18509 16837 18567 16843
rect 17494 16806 17500 16818
rect 17455 16778 17500 16806
rect 17494 16766 17500 16778
rect 17552 16766 17558 16818
rect 18322 16766 18328 16818
rect 18380 16806 18386 16818
rect 18417 16809 18475 16815
rect 18417 16806 18429 16809
rect 18380 16778 18429 16806
rect 18380 16766 18386 16778
rect 18417 16775 18429 16778
rect 18463 16775 18475 16809
rect 18417 16769 18475 16775
rect 1104 16716 28888 16738
rect 1104 16664 10982 16716
rect 11034 16664 11046 16716
rect 11098 16664 11110 16716
rect 11162 16664 11174 16716
rect 11226 16664 20982 16716
rect 21034 16664 21046 16716
rect 21098 16664 21110 16716
rect 21162 16664 21174 16716
rect 21226 16664 28888 16716
rect 1104 16642 28888 16664
rect 14182 16562 14188 16614
rect 14240 16602 14246 16614
rect 14369 16605 14427 16611
rect 14369 16602 14381 16605
rect 14240 16574 14381 16602
rect 14240 16562 14246 16574
rect 14369 16571 14381 16574
rect 14415 16602 14427 16605
rect 15194 16602 15200 16614
rect 14415 16574 15200 16602
rect 14415 16571 14427 16574
rect 14369 16565 14427 16571
rect 15194 16562 15200 16574
rect 15252 16562 15258 16614
rect 18322 16602 18328 16614
rect 18283 16574 18328 16602
rect 18322 16562 18328 16574
rect 18380 16562 18386 16614
rect 12986 16466 12992 16478
rect 12947 16438 12992 16466
rect 12986 16426 12992 16438
rect 13044 16426 13050 16478
rect 13256 16469 13314 16475
rect 13256 16435 13268 16469
rect 13302 16466 13314 16469
rect 13722 16466 13728 16478
rect 13302 16438 13728 16466
rect 13302 16435 13314 16438
rect 13256 16429 13314 16435
rect 13722 16426 13728 16438
rect 13780 16426 13786 16478
rect 1104 16172 28888 16194
rect 1104 16120 5982 16172
rect 6034 16120 6046 16172
rect 6098 16120 6110 16172
rect 6162 16120 6174 16172
rect 6226 16120 15982 16172
rect 16034 16120 16046 16172
rect 16098 16120 16110 16172
rect 16162 16120 16174 16172
rect 16226 16120 25982 16172
rect 26034 16120 26046 16172
rect 26098 16120 26110 16172
rect 26162 16120 26174 16172
rect 26226 16120 28888 16172
rect 1104 16098 28888 16120
rect 7006 16058 7012 16070
rect 6967 16030 7012 16058
rect 7006 16018 7012 16030
rect 7064 16018 7070 16070
rect 12986 16058 12992 16070
rect 12947 16030 12992 16058
rect 12986 16018 12992 16030
rect 13044 16018 13050 16070
rect 24486 16058 24492 16070
rect 24447 16030 24492 16058
rect 24486 16018 24492 16030
rect 24544 16018 24550 16070
rect 7024 15922 7052 16018
rect 7101 15925 7159 15931
rect 7101 15922 7113 15925
rect 7024 15894 7113 15922
rect 7101 15891 7113 15894
rect 7147 15891 7159 15925
rect 7101 15885 7159 15891
rect 23937 15857 23995 15863
rect 23937 15823 23949 15857
rect 23983 15854 23995 15857
rect 24486 15854 24492 15866
rect 23983 15826 24492 15854
rect 23983 15823 23995 15826
rect 23937 15817 23995 15823
rect 24486 15814 24492 15826
rect 24544 15814 24550 15866
rect 7190 15746 7196 15798
rect 7248 15786 7254 15798
rect 7346 15789 7404 15795
rect 7346 15786 7358 15789
rect 7248 15758 7358 15786
rect 7248 15746 7254 15758
rect 7346 15755 7358 15758
rect 7392 15755 7404 15789
rect 7346 15749 7404 15755
rect 8481 15721 8539 15727
rect 8481 15687 8493 15721
rect 8527 15718 8539 15721
rect 8570 15718 8576 15730
rect 8527 15690 8576 15718
rect 8527 15687 8539 15690
rect 8481 15681 8539 15687
rect 8570 15678 8576 15690
rect 8628 15718 8634 15730
rect 13449 15721 13507 15727
rect 13449 15718 13461 15721
rect 8628 15690 13461 15718
rect 8628 15678 8634 15690
rect 13449 15687 13461 15690
rect 13495 15718 13507 15721
rect 13722 15718 13728 15730
rect 13495 15690 13728 15718
rect 13495 15687 13507 15690
rect 13449 15681 13507 15687
rect 13722 15678 13728 15690
rect 13780 15678 13786 15730
rect 23658 15678 23664 15730
rect 23716 15718 23722 15730
rect 24121 15721 24179 15727
rect 24121 15718 24133 15721
rect 23716 15690 24133 15718
rect 23716 15678 23722 15690
rect 24121 15687 24133 15690
rect 24167 15687 24179 15721
rect 24121 15681 24179 15687
rect 1104 15628 28888 15650
rect 1104 15576 10982 15628
rect 11034 15576 11046 15628
rect 11098 15576 11110 15628
rect 11162 15576 11174 15628
rect 11226 15576 20982 15628
rect 21034 15576 21046 15628
rect 21098 15576 21110 15628
rect 21162 15576 21174 15628
rect 21226 15576 28888 15628
rect 1104 15554 28888 15576
rect 7190 15514 7196 15526
rect 7151 15486 7196 15514
rect 7190 15474 7196 15486
rect 7248 15474 7254 15526
rect 23937 15381 23995 15387
rect 23937 15347 23949 15381
rect 23983 15378 23995 15381
rect 24026 15378 24032 15390
rect 23983 15350 24032 15378
rect 23983 15347 23995 15350
rect 23937 15341 23995 15347
rect 24026 15338 24032 15350
rect 24084 15378 24090 15390
rect 24762 15378 24768 15390
rect 24084 15350 24768 15378
rect 24084 15338 24090 15350
rect 24762 15338 24768 15350
rect 24820 15338 24826 15390
rect 18598 15174 18604 15186
rect 18559 15146 18604 15174
rect 18598 15134 18604 15146
rect 18656 15134 18662 15186
rect 23750 15134 23756 15186
rect 23808 15174 23814 15186
rect 24121 15177 24179 15183
rect 24121 15174 24133 15177
rect 23808 15146 24133 15174
rect 23808 15134 23814 15146
rect 24121 15143 24133 15146
rect 24167 15143 24179 15177
rect 24121 15137 24179 15143
rect 1104 15084 28888 15106
rect 1104 15032 5982 15084
rect 6034 15032 6046 15084
rect 6098 15032 6110 15084
rect 6162 15032 6174 15084
rect 6226 15032 15982 15084
rect 16034 15032 16046 15084
rect 16098 15032 16110 15084
rect 16162 15032 16174 15084
rect 16226 15032 25982 15084
rect 26034 15032 26046 15084
rect 26098 15032 26110 15084
rect 26162 15032 26174 15084
rect 26226 15032 28888 15084
rect 1104 15010 28888 15032
rect 18322 14930 18328 14982
rect 18380 14970 18386 14982
rect 18509 14973 18567 14979
rect 18509 14970 18521 14973
rect 18380 14942 18521 14970
rect 18380 14930 18386 14942
rect 18509 14939 18521 14942
rect 18555 14939 18567 14973
rect 24026 14970 24032 14982
rect 23987 14942 24032 14970
rect 18509 14933 18567 14939
rect 24026 14930 24032 14942
rect 24084 14930 24090 14982
rect 18322 14834 18328 14846
rect 18283 14806 18328 14834
rect 18322 14794 18328 14806
rect 18380 14834 18386 14846
rect 19061 14837 19119 14843
rect 19061 14834 19073 14837
rect 18380 14806 19073 14834
rect 18380 14794 18386 14806
rect 19061 14803 19073 14806
rect 19107 14803 19119 14837
rect 19061 14797 19119 14803
rect 18598 14658 18604 14710
rect 18656 14698 18662 14710
rect 18877 14701 18935 14707
rect 18877 14698 18889 14701
rect 18656 14670 18889 14698
rect 18656 14658 18662 14670
rect 18877 14667 18889 14670
rect 18923 14698 18935 14701
rect 19242 14698 19248 14710
rect 18923 14670 19248 14698
rect 18923 14667 18935 14670
rect 18877 14661 18935 14667
rect 19242 14658 19248 14670
rect 19300 14658 19306 14710
rect 18966 14630 18972 14642
rect 18927 14602 18972 14630
rect 18966 14590 18972 14602
rect 19024 14590 19030 14642
rect 1104 14540 28888 14562
rect 1104 14488 10982 14540
rect 11034 14488 11046 14540
rect 11098 14488 11110 14540
rect 11162 14488 11174 14540
rect 11226 14488 20982 14540
rect 21034 14488 21046 14540
rect 21098 14488 21110 14540
rect 21162 14488 21174 14540
rect 21226 14488 28888 14540
rect 1104 14466 28888 14488
rect 18601 14429 18659 14435
rect 18601 14395 18613 14429
rect 18647 14426 18659 14429
rect 18966 14426 18972 14438
rect 18647 14398 18972 14426
rect 18647 14395 18659 14398
rect 18601 14389 18659 14395
rect 18966 14386 18972 14398
rect 19024 14426 19030 14438
rect 19429 14429 19487 14435
rect 19429 14426 19441 14429
rect 19024 14398 19441 14426
rect 19024 14386 19030 14398
rect 19429 14395 19441 14398
rect 19475 14395 19487 14429
rect 19429 14389 19487 14395
rect 19610 14250 19616 14302
rect 19668 14290 19674 14302
rect 19794 14290 19800 14302
rect 19668 14262 19800 14290
rect 19668 14250 19674 14262
rect 19794 14250 19800 14262
rect 19852 14250 19858 14302
rect 19886 14222 19892 14234
rect 19847 14194 19892 14222
rect 19886 14182 19892 14194
rect 19944 14182 19950 14234
rect 20073 14225 20131 14231
rect 20073 14191 20085 14225
rect 20119 14222 20131 14225
rect 20438 14222 20444 14234
rect 20119 14194 20444 14222
rect 20119 14191 20131 14194
rect 20073 14185 20131 14191
rect 20438 14182 20444 14194
rect 20496 14182 20502 14234
rect 1104 13996 28888 14018
rect 1104 13944 5982 13996
rect 6034 13944 6046 13996
rect 6098 13944 6110 13996
rect 6162 13944 6174 13996
rect 6226 13944 15982 13996
rect 16034 13944 16046 13996
rect 16098 13944 16110 13996
rect 16162 13944 16174 13996
rect 16226 13944 25982 13996
rect 26034 13944 26046 13996
rect 26098 13944 26110 13996
rect 26162 13944 26174 13996
rect 26226 13944 28888 13996
rect 1104 13922 28888 13944
rect 24854 13842 24860 13894
rect 24912 13882 24918 13894
rect 25314 13882 25320 13894
rect 24912 13854 25320 13882
rect 24912 13842 24918 13854
rect 25314 13842 25320 13854
rect 25372 13842 25378 13894
rect 19610 13678 19616 13690
rect 19571 13650 19616 13678
rect 19610 13638 19616 13650
rect 19668 13638 19674 13690
rect 19886 13678 19892 13690
rect 19847 13650 19892 13678
rect 19886 13638 19892 13650
rect 19944 13638 19950 13690
rect 24210 13638 24216 13690
rect 24268 13678 24274 13690
rect 24762 13678 24768 13690
rect 24268 13650 24768 13678
rect 24268 13638 24274 13650
rect 24762 13638 24768 13650
rect 24820 13638 24826 13690
rect 19058 13542 19064 13554
rect 19019 13514 19064 13542
rect 19058 13502 19064 13514
rect 19116 13502 19122 13554
rect 20349 13545 20407 13551
rect 20349 13511 20361 13545
rect 20395 13542 20407 13545
rect 20438 13542 20444 13554
rect 20395 13514 20444 13542
rect 20395 13511 20407 13514
rect 20349 13505 20407 13511
rect 20438 13502 20444 13514
rect 20496 13502 20502 13554
rect 1104 13452 28888 13474
rect 1104 13400 10982 13452
rect 11034 13400 11046 13452
rect 11098 13400 11110 13452
rect 11162 13400 11174 13452
rect 11226 13400 20982 13452
rect 21034 13400 21046 13452
rect 21098 13400 21110 13452
rect 21162 13400 21174 13452
rect 21226 13400 28888 13452
rect 1104 13378 28888 13400
rect 13538 13338 13544 13350
rect 13499 13310 13544 13338
rect 13538 13298 13544 13310
rect 13596 13298 13602 13350
rect 19058 13298 19064 13350
rect 19116 13338 19122 13350
rect 20070 13338 20076 13350
rect 19116 13310 20076 13338
rect 19116 13298 19122 13310
rect 20070 13298 20076 13310
rect 20128 13298 20134 13350
rect 1397 13205 1455 13211
rect 1397 13171 1409 13205
rect 1443 13202 1455 13205
rect 1486 13202 1492 13214
rect 1443 13174 1492 13202
rect 1443 13171 1455 13174
rect 1397 13165 1455 13171
rect 1486 13162 1492 13174
rect 1544 13162 1550 13214
rect 13906 13202 13912 13214
rect 13867 13174 13912 13202
rect 13906 13162 13912 13174
rect 13964 13162 13970 13214
rect 19702 13162 19708 13214
rect 19760 13202 19766 13214
rect 20162 13202 20168 13214
rect 19760 13174 20168 13202
rect 19760 13162 19766 13174
rect 20162 13162 20168 13174
rect 20220 13162 20226 13214
rect 13814 13094 13820 13146
rect 13872 13134 13878 13146
rect 14001 13137 14059 13143
rect 14001 13134 14013 13137
rect 13872 13106 14013 13134
rect 13872 13094 13878 13106
rect 14001 13103 14013 13106
rect 14047 13103 14059 13137
rect 14182 13134 14188 13146
rect 14143 13106 14188 13134
rect 14001 13097 14059 13103
rect 14182 13094 14188 13106
rect 14240 13094 14246 13146
rect 20349 13137 20407 13143
rect 20349 13103 20361 13137
rect 20395 13134 20407 13137
rect 20438 13134 20444 13146
rect 20395 13106 20444 13134
rect 20395 13103 20407 13106
rect 20349 13097 20407 13103
rect 20438 13094 20444 13106
rect 20496 13094 20502 13146
rect 19334 13026 19340 13078
rect 19392 13066 19398 13078
rect 19705 13069 19763 13075
rect 19705 13066 19717 13069
rect 19392 13038 19717 13066
rect 19392 13026 19398 13038
rect 19705 13035 19717 13038
rect 19751 13035 19763 13069
rect 19705 13029 19763 13035
rect 1581 13001 1639 13007
rect 1581 12967 1593 13001
rect 1627 12998 1639 13001
rect 2130 12998 2136 13010
rect 1627 12970 2136 12998
rect 1627 12967 1639 12970
rect 1581 12961 1639 12967
rect 2130 12958 2136 12970
rect 2188 12958 2194 13010
rect 13078 12998 13084 13010
rect 13039 12970 13084 12998
rect 13078 12958 13084 12970
rect 13136 12958 13142 13010
rect 1104 12908 28888 12930
rect 1104 12856 5982 12908
rect 6034 12856 6046 12908
rect 6098 12856 6110 12908
rect 6162 12856 6174 12908
rect 6226 12856 15982 12908
rect 16034 12856 16046 12908
rect 16098 12856 16110 12908
rect 16162 12856 16174 12908
rect 16226 12856 25982 12908
rect 26034 12856 26046 12908
rect 26098 12856 26110 12908
rect 26162 12856 26174 12908
rect 26226 12856 28888 12908
rect 1104 12834 28888 12856
rect 14182 12794 14188 12806
rect 14143 12766 14188 12794
rect 14182 12754 14188 12766
rect 14240 12754 14246 12806
rect 20070 12794 20076 12806
rect 20031 12766 20076 12794
rect 20070 12754 20076 12766
rect 20128 12754 20134 12806
rect 13081 12729 13139 12735
rect 13081 12695 13093 12729
rect 13127 12726 13139 12729
rect 13906 12726 13912 12738
rect 13127 12698 13912 12726
rect 13127 12695 13139 12698
rect 13081 12689 13139 12695
rect 13906 12686 13912 12698
rect 13964 12686 13970 12738
rect 13722 12658 13728 12670
rect 13683 12630 13728 12658
rect 13722 12618 13728 12630
rect 13780 12618 13786 12670
rect 1394 12590 1400 12602
rect 1355 12562 1400 12590
rect 1394 12550 1400 12562
rect 1452 12590 1458 12602
rect 1949 12593 2007 12599
rect 1949 12590 1961 12593
rect 1452 12562 1961 12590
rect 1452 12550 1458 12562
rect 1949 12559 1961 12562
rect 1995 12559 2007 12593
rect 12894 12590 12900 12602
rect 12855 12562 12900 12590
rect 1949 12553 2007 12559
rect 12894 12550 12900 12562
rect 12952 12590 12958 12602
rect 13449 12593 13507 12599
rect 13449 12590 13461 12593
rect 12952 12562 13461 12590
rect 12952 12550 12958 12562
rect 13449 12559 13461 12562
rect 13495 12559 13507 12593
rect 13449 12553 13507 12559
rect 12434 12482 12440 12534
rect 12492 12522 12498 12534
rect 13078 12522 13084 12534
rect 12492 12494 13084 12522
rect 12492 12482 12498 12494
rect 13078 12482 13084 12494
rect 13136 12522 13142 12534
rect 13541 12525 13599 12531
rect 13541 12522 13553 12525
rect 13136 12494 13553 12522
rect 13136 12482 13142 12494
rect 13541 12491 13553 12494
rect 13587 12491 13599 12525
rect 13541 12485 13599 12491
rect 1486 12414 1492 12466
rect 1544 12454 1550 12466
rect 1581 12457 1639 12463
rect 1581 12454 1593 12457
rect 1544 12426 1593 12454
rect 1544 12414 1550 12426
rect 1581 12423 1593 12426
rect 1627 12423 1639 12457
rect 19702 12454 19708 12466
rect 19663 12426 19708 12454
rect 1581 12417 1639 12423
rect 19702 12414 19708 12426
rect 19760 12414 19766 12466
rect 20438 12454 20444 12466
rect 20399 12426 20444 12454
rect 20438 12414 20444 12426
rect 20496 12414 20502 12466
rect 1104 12364 28888 12386
rect 1104 12312 10982 12364
rect 11034 12312 11046 12364
rect 11098 12312 11110 12364
rect 11162 12312 11174 12364
rect 11226 12312 20982 12364
rect 21034 12312 21046 12364
rect 21098 12312 21110 12364
rect 21162 12312 21174 12364
rect 21226 12312 28888 12364
rect 1104 12290 28888 12312
rect 1578 12250 1584 12262
rect 1539 12222 1584 12250
rect 1578 12210 1584 12222
rect 1636 12210 1642 12262
rect 3602 12210 3608 12262
rect 3660 12250 3666 12262
rect 3878 12250 3884 12262
rect 3660 12222 3884 12250
rect 3660 12210 3666 12222
rect 3878 12210 3884 12222
rect 3936 12210 3942 12262
rect 13906 12250 13912 12262
rect 13867 12222 13912 12250
rect 13906 12210 13912 12222
rect 13964 12210 13970 12262
rect 13173 12185 13231 12191
rect 13173 12151 13185 12185
rect 13219 12182 13231 12185
rect 13722 12182 13728 12194
rect 13219 12154 13728 12182
rect 13219 12151 13231 12154
rect 13173 12145 13231 12151
rect 13722 12142 13728 12154
rect 13780 12142 13786 12194
rect 8297 12117 8355 12123
rect 8297 12083 8309 12117
rect 8343 12114 8355 12117
rect 8662 12114 8668 12126
rect 8343 12086 8668 12114
rect 8343 12083 8355 12086
rect 8297 12077 8355 12083
rect 8662 12074 8668 12086
rect 8720 12074 8726 12126
rect 8389 12049 8447 12055
rect 8389 12015 8401 12049
rect 8435 12015 8447 12049
rect 8570 12046 8576 12058
rect 8531 12018 8576 12046
rect 8389 12009 8447 12015
rect 7926 11978 7932 11990
rect 7887 11950 7932 11978
rect 7926 11938 7932 11950
rect 7984 11938 7990 11990
rect 8294 11938 8300 11990
rect 8352 11978 8358 11990
rect 8404 11978 8432 12009
rect 8570 12006 8576 12018
rect 8628 12006 8634 12058
rect 8352 11950 8432 11978
rect 13633 11981 13691 11987
rect 8352 11938 8358 11950
rect 13633 11947 13645 11981
rect 13679 11978 13691 11981
rect 13722 11978 13728 11990
rect 13679 11950 13728 11978
rect 13679 11947 13691 11950
rect 13633 11941 13691 11947
rect 13722 11938 13728 11950
rect 13780 11938 13786 11990
rect 12066 11910 12072 11922
rect 12027 11882 12072 11910
rect 12066 11870 12072 11882
rect 12124 11870 12130 11922
rect 1104 11820 28888 11842
rect 1104 11768 5982 11820
rect 6034 11768 6046 11820
rect 6098 11768 6110 11820
rect 6162 11768 6174 11820
rect 6226 11768 15982 11820
rect 16034 11768 16046 11820
rect 16098 11768 16110 11820
rect 16162 11768 16174 11820
rect 16226 11768 25982 11820
rect 26034 11768 26046 11820
rect 26098 11768 26110 11820
rect 26162 11768 26174 11820
rect 26226 11768 28888 11820
rect 1104 11746 28888 11768
rect 8021 11709 8079 11715
rect 8021 11675 8033 11709
rect 8067 11706 8079 11709
rect 8570 11706 8576 11718
rect 8067 11678 8576 11706
rect 8067 11675 8079 11678
rect 8021 11669 8079 11675
rect 8570 11666 8576 11678
rect 8628 11666 8634 11718
rect 11882 11706 11888 11718
rect 11843 11678 11888 11706
rect 11882 11666 11888 11678
rect 11940 11666 11946 11718
rect 12069 11709 12127 11715
rect 12069 11675 12081 11709
rect 12115 11706 12127 11709
rect 12342 11706 12348 11718
rect 12115 11678 12348 11706
rect 12115 11675 12127 11678
rect 12069 11669 12127 11675
rect 12342 11666 12348 11678
rect 12400 11666 12406 11718
rect 24121 11641 24179 11647
rect 24121 11607 24133 11641
rect 24167 11638 24179 11641
rect 24854 11638 24860 11650
rect 24167 11610 24860 11638
rect 24167 11607 24179 11610
rect 24121 11601 24179 11607
rect 24854 11598 24860 11610
rect 24912 11598 24918 11650
rect 12066 11530 12072 11582
rect 12124 11570 12130 11582
rect 12621 11573 12679 11579
rect 12621 11570 12633 11573
rect 12124 11542 12633 11570
rect 12124 11530 12130 11542
rect 12621 11539 12633 11542
rect 12667 11539 12679 11573
rect 12621 11533 12679 11539
rect 1397 11505 1455 11511
rect 1397 11471 1409 11505
rect 1443 11502 1455 11505
rect 1670 11502 1676 11514
rect 1443 11474 1676 11502
rect 1443 11471 1455 11474
rect 1397 11465 1455 11471
rect 1670 11462 1676 11474
rect 1728 11502 1734 11514
rect 1949 11505 2007 11511
rect 1949 11502 1961 11505
rect 1728 11474 1961 11502
rect 1728 11462 1734 11474
rect 1949 11471 1961 11474
rect 1995 11471 2007 11505
rect 1949 11465 2007 11471
rect 11882 11462 11888 11514
rect 11940 11502 11946 11514
rect 12526 11502 12532 11514
rect 11940 11474 12532 11502
rect 11940 11462 11946 11474
rect 12526 11462 12532 11474
rect 12584 11462 12590 11514
rect 23474 11462 23480 11514
rect 23532 11502 23538 11514
rect 23937 11505 23995 11511
rect 23937 11502 23949 11505
rect 23532 11474 23949 11502
rect 23532 11462 23538 11474
rect 23937 11471 23949 11474
rect 23983 11502 23995 11505
rect 24489 11505 24547 11511
rect 24489 11502 24501 11505
rect 23983 11474 24501 11502
rect 23983 11471 23995 11474
rect 23937 11465 23995 11471
rect 24489 11471 24501 11474
rect 24535 11471 24547 11505
rect 24489 11465 24547 11471
rect 11514 11394 11520 11446
rect 11572 11434 11578 11446
rect 12437 11437 12495 11443
rect 12437 11434 12449 11437
rect 11572 11406 12449 11434
rect 11572 11394 11578 11406
rect 12437 11403 12449 11406
rect 12483 11434 12495 11437
rect 13722 11434 13728 11446
rect 12483 11406 13728 11434
rect 12483 11403 12495 11406
rect 12437 11397 12495 11403
rect 13722 11394 13728 11406
rect 13780 11394 13786 11446
rect 1581 11369 1639 11375
rect 1581 11335 1593 11369
rect 1627 11366 1639 11369
rect 2222 11366 2228 11378
rect 1627 11338 2228 11366
rect 1627 11335 1639 11338
rect 1581 11329 1639 11335
rect 2222 11326 2228 11338
rect 2280 11326 2286 11378
rect 8294 11366 8300 11378
rect 8255 11338 8300 11366
rect 8294 11326 8300 11338
rect 8352 11326 8358 11378
rect 8662 11366 8668 11378
rect 8623 11338 8668 11366
rect 8662 11326 8668 11338
rect 8720 11326 8726 11378
rect 12526 11366 12532 11378
rect 12487 11338 12532 11366
rect 12526 11326 12532 11338
rect 12584 11326 12590 11378
rect 1104 11276 28888 11298
rect 1104 11224 10982 11276
rect 11034 11224 11046 11276
rect 11098 11224 11110 11276
rect 11162 11224 11174 11276
rect 11226 11224 20982 11276
rect 21034 11224 21046 11276
rect 21098 11224 21110 11276
rect 21162 11224 21174 11276
rect 21226 11224 28888 11276
rect 1104 11202 28888 11224
rect 7745 11165 7803 11171
rect 7745 11131 7757 11165
rect 7791 11162 7803 11165
rect 8662 11162 8668 11174
rect 7791 11134 8668 11162
rect 7791 11131 7803 11134
rect 7745 11125 7803 11131
rect 8662 11122 8668 11134
rect 8720 11122 8726 11174
rect 11514 11122 11520 11174
rect 11572 11162 11578 11174
rect 12069 11165 12127 11171
rect 12069 11162 12081 11165
rect 11572 11134 12081 11162
rect 11572 11122 11578 11134
rect 12069 11131 12081 11134
rect 12115 11131 12127 11165
rect 12069 11125 12127 11131
rect 7190 11054 7196 11106
rect 7248 11094 7254 11106
rect 7248 11066 8248 11094
rect 7248 11054 7254 11066
rect 1397 11029 1455 11035
rect 1397 10995 1409 11029
rect 1443 11026 1455 11029
rect 2038 11026 2044 11038
rect 1443 10998 2044 11026
rect 1443 10995 1455 10998
rect 1397 10989 1455 10995
rect 2038 10986 2044 10998
rect 2096 10986 2102 11038
rect 8110 11026 8116 11038
rect 8071 10998 8116 11026
rect 8110 10986 8116 10998
rect 8168 10986 8174 11038
rect 8220 11026 8248 11066
rect 23937 11029 23995 11035
rect 8220 10998 8432 11026
rect 8404 10970 8432 10998
rect 23937 10995 23949 11029
rect 23983 11026 23995 11029
rect 24026 11026 24032 11038
rect 23983 10998 24032 11026
rect 23983 10995 23995 10998
rect 23937 10989 23995 10995
rect 24026 10986 24032 10998
rect 24084 11026 24090 11038
rect 24394 11026 24400 11038
rect 24084 10998 24400 11026
rect 24084 10986 24090 10998
rect 24394 10986 24400 10998
rect 24452 10986 24458 11038
rect 7374 10918 7380 10970
rect 7432 10958 7438 10970
rect 8205 10961 8263 10967
rect 8205 10958 8217 10961
rect 7432 10930 8217 10958
rect 7432 10918 7438 10930
rect 8205 10927 8217 10930
rect 8251 10927 8263 10961
rect 8205 10921 8263 10927
rect 8386 10918 8392 10970
rect 8444 10958 8450 10970
rect 8444 10930 8537 10958
rect 8444 10918 8450 10930
rect 1581 10893 1639 10899
rect 1581 10859 1593 10893
rect 1627 10890 1639 10893
rect 1946 10890 1952 10902
rect 1627 10862 1952 10890
rect 1627 10859 1639 10862
rect 1581 10853 1639 10859
rect 1946 10850 1952 10862
rect 2004 10850 2010 10902
rect 24118 10890 24124 10902
rect 24079 10862 24124 10890
rect 24118 10850 24124 10862
rect 24176 10850 24182 10902
rect 1104 10732 28888 10754
rect 1104 10680 5982 10732
rect 6034 10680 6046 10732
rect 6098 10680 6110 10732
rect 6162 10680 6174 10732
rect 6226 10680 15982 10732
rect 16034 10680 16046 10732
rect 16098 10680 16110 10732
rect 16162 10680 16174 10732
rect 16226 10680 25982 10732
rect 26034 10680 26046 10732
rect 26098 10680 26110 10732
rect 26162 10680 26174 10732
rect 26226 10680 28888 10732
rect 1104 10658 28888 10680
rect 2038 10618 2044 10630
rect 1999 10590 2044 10618
rect 2038 10578 2044 10590
rect 2096 10578 2102 10630
rect 2406 10618 2412 10630
rect 2367 10590 2412 10618
rect 2406 10578 2412 10590
rect 2464 10578 2470 10630
rect 7929 10621 7987 10627
rect 7929 10587 7941 10621
rect 7975 10618 7987 10621
rect 8202 10618 8208 10630
rect 7975 10590 8208 10618
rect 7975 10587 7987 10590
rect 7929 10581 7987 10587
rect 8202 10578 8208 10590
rect 8260 10578 8266 10630
rect 8386 10578 8392 10630
rect 8444 10618 8450 10630
rect 8941 10621 8999 10627
rect 8941 10618 8953 10621
rect 8444 10590 8953 10618
rect 8444 10578 8450 10590
rect 7098 10550 7104 10562
rect 7011 10522 7104 10550
rect 7098 10510 7104 10522
rect 7156 10550 7162 10562
rect 8110 10550 8116 10562
rect 7156 10522 8116 10550
rect 7156 10510 7162 10522
rect 8110 10510 8116 10522
rect 8168 10510 8174 10562
rect 8588 10491 8616 10590
rect 8941 10587 8953 10590
rect 8987 10587 8999 10621
rect 24026 10618 24032 10630
rect 23987 10590 24032 10618
rect 8941 10581 8999 10587
rect 24026 10578 24032 10590
rect 24084 10578 24090 10630
rect 8573 10485 8631 10491
rect 8573 10451 8585 10485
rect 8619 10451 8631 10485
rect 8573 10445 8631 10451
rect 1397 10417 1455 10423
rect 1397 10383 1409 10417
rect 1443 10414 1455 10417
rect 2406 10414 2412 10426
rect 1443 10386 2412 10414
rect 1443 10383 1455 10386
rect 1397 10377 1455 10383
rect 2406 10374 2412 10386
rect 2464 10374 2470 10426
rect 8294 10346 8300 10358
rect 8255 10318 8300 10346
rect 8294 10306 8300 10318
rect 8352 10306 8358 10358
rect 1581 10281 1639 10287
rect 1581 10247 1593 10281
rect 1627 10278 1639 10281
rect 1762 10278 1768 10290
rect 1627 10250 1768 10278
rect 1627 10247 1639 10250
rect 1581 10241 1639 10247
rect 1762 10238 1768 10250
rect 1820 10238 1826 10290
rect 7374 10278 7380 10290
rect 7335 10250 7380 10278
rect 7374 10238 7380 10250
rect 7432 10238 7438 10290
rect 7834 10278 7840 10290
rect 7747 10250 7840 10278
rect 7834 10238 7840 10250
rect 7892 10278 7898 10290
rect 8386 10278 8392 10290
rect 7892 10250 8392 10278
rect 7892 10238 7898 10250
rect 8386 10238 8392 10250
rect 8444 10238 8450 10290
rect 1104 10188 28888 10210
rect 1104 10136 10982 10188
rect 11034 10136 11046 10188
rect 11098 10136 11110 10188
rect 11162 10136 11174 10188
rect 11226 10136 20982 10188
rect 21034 10136 21046 10188
rect 21098 10136 21110 10188
rect 21162 10136 21174 10188
rect 21226 10136 28888 10188
rect 1104 10114 28888 10136
rect 8021 10077 8079 10083
rect 8021 10043 8033 10077
rect 8067 10074 8079 10077
rect 8294 10074 8300 10086
rect 8067 10046 8300 10074
rect 8067 10043 8079 10046
rect 8021 10037 8079 10043
rect 8294 10034 8300 10046
rect 8352 10034 8358 10086
rect 8389 10077 8447 10083
rect 8389 10043 8401 10077
rect 8435 10074 8447 10077
rect 8478 10074 8484 10086
rect 8435 10046 8484 10074
rect 8435 10043 8447 10046
rect 8389 10037 8447 10043
rect 8478 10034 8484 10046
rect 8536 10034 8542 10086
rect 1397 9941 1455 9947
rect 1397 9907 1409 9941
rect 1443 9938 1455 9941
rect 2038 9938 2044 9950
rect 1443 9910 2044 9938
rect 1443 9907 1455 9910
rect 1397 9901 1455 9907
rect 2038 9898 2044 9910
rect 2096 9898 2102 9950
rect 1578 9734 1584 9746
rect 1539 9706 1584 9734
rect 1578 9694 1584 9706
rect 1636 9694 1642 9746
rect 1104 9644 28888 9666
rect 1104 9592 5982 9644
rect 6034 9592 6046 9644
rect 6098 9592 6110 9644
rect 6162 9592 6174 9644
rect 6226 9592 15982 9644
rect 16034 9592 16046 9644
rect 16098 9592 16110 9644
rect 16162 9592 16174 9644
rect 16226 9592 25982 9644
rect 26034 9592 26046 9644
rect 26098 9592 26110 9644
rect 26162 9592 26174 9644
rect 26226 9592 28888 9644
rect 1104 9570 28888 9592
rect 2038 9530 2044 9542
rect 1999 9502 2044 9530
rect 2038 9490 2044 9502
rect 2096 9490 2102 9542
rect 2409 9465 2467 9471
rect 2409 9431 2421 9465
rect 2455 9462 2467 9465
rect 2498 9462 2504 9474
rect 2455 9434 2504 9462
rect 2455 9431 2467 9434
rect 2409 9425 2467 9431
rect 1397 9329 1455 9335
rect 1397 9295 1409 9329
rect 1443 9326 1455 9329
rect 2424 9326 2452 9425
rect 2498 9422 2504 9434
rect 2556 9422 2562 9474
rect 23934 9326 23940 9338
rect 1443 9298 2452 9326
rect 23895 9298 23940 9326
rect 1443 9295 1455 9298
rect 1397 9289 1455 9295
rect 23934 9286 23940 9298
rect 23992 9326 23998 9338
rect 24489 9329 24547 9335
rect 24489 9326 24501 9329
rect 23992 9298 24501 9326
rect 23992 9286 23998 9298
rect 24489 9295 24501 9298
rect 24535 9295 24547 9329
rect 24489 9289 24547 9295
rect 1581 9193 1639 9199
rect 1581 9159 1593 9193
rect 1627 9190 1639 9193
rect 1670 9190 1676 9202
rect 1627 9162 1676 9190
rect 1627 9159 1639 9162
rect 1581 9153 1639 9159
rect 1670 9150 1676 9162
rect 1728 9150 1734 9202
rect 24118 9190 24124 9202
rect 24079 9162 24124 9190
rect 24118 9150 24124 9162
rect 24176 9150 24182 9202
rect 1104 9100 28888 9122
rect 1104 9048 10982 9100
rect 11034 9048 11046 9100
rect 11098 9048 11110 9100
rect 11162 9048 11174 9100
rect 11226 9048 20982 9100
rect 21034 9048 21046 9100
rect 21098 9048 21110 9100
rect 21162 9048 21174 9100
rect 21226 9048 28888 9100
rect 1104 9026 28888 9048
rect 1394 8850 1400 8862
rect 1355 8822 1400 8850
rect 1394 8810 1400 8822
rect 1452 8810 1458 8862
rect 23937 8853 23995 8859
rect 23937 8819 23949 8853
rect 23983 8850 23995 8853
rect 24486 8850 24492 8862
rect 23983 8822 24492 8850
rect 23983 8819 23995 8822
rect 23937 8813 23995 8819
rect 24486 8810 24492 8822
rect 24544 8810 24550 8862
rect 1486 8606 1492 8658
rect 1544 8646 1550 8658
rect 1581 8649 1639 8655
rect 1581 8646 1593 8649
rect 1544 8618 1593 8646
rect 1544 8606 1550 8618
rect 1581 8615 1593 8618
rect 1627 8615 1639 8649
rect 24118 8646 24124 8658
rect 24079 8618 24124 8646
rect 1581 8609 1639 8615
rect 24118 8606 24124 8618
rect 24176 8606 24182 8658
rect 1104 8556 28888 8578
rect 1104 8504 5982 8556
rect 6034 8504 6046 8556
rect 6098 8504 6110 8556
rect 6162 8504 6174 8556
rect 6226 8504 15982 8556
rect 16034 8504 16046 8556
rect 16098 8504 16110 8556
rect 16162 8504 16174 8556
rect 16226 8504 25982 8556
rect 26034 8504 26046 8556
rect 26098 8504 26110 8556
rect 26162 8504 26174 8556
rect 26226 8504 28888 8556
rect 1104 8482 28888 8504
rect 1394 8402 1400 8454
rect 1452 8442 1458 8454
rect 1581 8445 1639 8451
rect 1581 8442 1593 8445
rect 1452 8414 1593 8442
rect 1452 8402 1458 8414
rect 1581 8411 1593 8414
rect 1627 8411 1639 8445
rect 1581 8405 1639 8411
rect 23845 8445 23903 8451
rect 23845 8411 23857 8445
rect 23891 8442 23903 8445
rect 24578 8442 24584 8454
rect 23891 8414 24584 8442
rect 23891 8411 23903 8414
rect 23845 8405 23903 8411
rect 23474 8334 23480 8386
rect 23532 8374 23538 8386
rect 24121 8377 24179 8383
rect 24121 8374 24133 8377
rect 23532 8346 24133 8374
rect 23532 8334 23538 8346
rect 24121 8343 24133 8346
rect 24167 8343 24179 8377
rect 24121 8337 24179 8343
rect 1394 8266 1400 8318
rect 1452 8306 1458 8318
rect 1854 8306 1860 8318
rect 1452 8278 1860 8306
rect 1452 8266 1458 8278
rect 1854 8266 1860 8278
rect 1912 8266 1918 8318
rect 23937 8241 23995 8247
rect 23937 8207 23949 8241
rect 23983 8238 23995 8241
rect 24228 8238 24256 8414
rect 24578 8402 24584 8414
rect 24636 8402 24642 8454
rect 24486 8238 24492 8250
rect 23983 8210 24256 8238
rect 24447 8210 24492 8238
rect 23983 8207 23995 8210
rect 23937 8201 23995 8207
rect 24486 8198 24492 8210
rect 24544 8198 24550 8250
rect 10778 8062 10784 8114
rect 10836 8102 10842 8114
rect 11330 8102 11336 8114
rect 10836 8074 11336 8102
rect 10836 8062 10842 8074
rect 11330 8062 11336 8074
rect 11388 8062 11394 8114
rect 1104 8012 28888 8034
rect 1104 7960 10982 8012
rect 11034 7960 11046 8012
rect 11098 7960 11110 8012
rect 11162 7960 11174 8012
rect 11226 7960 20982 8012
rect 21034 7960 21046 8012
rect 21098 7960 21110 8012
rect 21162 7960 21174 8012
rect 21226 7960 28888 8012
rect 1104 7938 28888 7960
rect 24118 7898 24124 7910
rect 24079 7870 24124 7898
rect 24118 7858 24124 7870
rect 24176 7858 24182 7910
rect 23934 7762 23940 7774
rect 23895 7734 23940 7762
rect 23934 7722 23940 7734
rect 23992 7722 23998 7774
rect 1104 7468 28888 7490
rect 1104 7416 5982 7468
rect 6034 7416 6046 7468
rect 6098 7416 6110 7468
rect 6162 7416 6174 7468
rect 6226 7416 15982 7468
rect 16034 7416 16046 7468
rect 16098 7416 16110 7468
rect 16162 7416 16174 7468
rect 16226 7416 25982 7468
rect 26034 7416 26046 7468
rect 26098 7416 26110 7468
rect 26162 7416 26174 7468
rect 26226 7416 28888 7468
rect 1104 7394 28888 7416
rect 22646 7354 22652 7366
rect 22607 7326 22652 7354
rect 22646 7314 22652 7326
rect 22704 7314 22710 7366
rect 23106 7354 23112 7366
rect 23067 7326 23112 7354
rect 23106 7314 23112 7326
rect 23164 7314 23170 7366
rect 18874 7286 18880 7298
rect 18835 7258 18880 7286
rect 18874 7246 18880 7258
rect 18932 7246 18938 7298
rect 18690 7150 18696 7162
rect 18651 7122 18696 7150
rect 18690 7110 18696 7122
rect 18748 7150 18754 7162
rect 19245 7153 19303 7159
rect 19245 7150 19257 7153
rect 18748 7122 19257 7150
rect 18748 7110 18754 7122
rect 19245 7119 19257 7122
rect 19291 7119 19303 7153
rect 19245 7113 19303 7119
rect 22465 7153 22523 7159
rect 22465 7119 22477 7153
rect 22511 7150 22523 7153
rect 23106 7150 23112 7162
rect 22511 7122 23112 7150
rect 22511 7119 22523 7122
rect 22465 7113 22523 7119
rect 23106 7110 23112 7122
rect 23164 7110 23170 7162
rect 23934 7150 23940 7162
rect 23895 7122 23940 7150
rect 23934 7110 23940 7122
rect 23992 7110 23998 7162
rect 1104 6924 28888 6946
rect 1104 6872 10982 6924
rect 11034 6872 11046 6924
rect 11098 6872 11110 6924
rect 11162 6872 11174 6924
rect 11226 6872 20982 6924
rect 21034 6872 21046 6924
rect 21098 6872 21110 6924
rect 21162 6872 21174 6924
rect 21226 6872 28888 6924
rect 1104 6850 28888 6872
rect 1578 6634 1584 6686
rect 1636 6674 1642 6686
rect 1854 6674 1860 6686
rect 1636 6646 1860 6674
rect 1636 6634 1642 6646
rect 1854 6634 1860 6646
rect 1912 6634 1918 6686
rect 10870 6674 10876 6686
rect 10831 6646 10876 6674
rect 10870 6634 10876 6646
rect 10928 6634 10934 6686
rect 14642 6674 14648 6686
rect 14603 6646 14648 6674
rect 14642 6634 14648 6646
rect 14700 6634 14706 6686
rect 23934 6674 23940 6686
rect 23847 6646 23940 6674
rect 23934 6634 23940 6646
rect 23992 6674 23998 6686
rect 24118 6674 24124 6686
rect 23992 6646 24124 6674
rect 23992 6634 23998 6646
rect 24118 6634 24124 6646
rect 24176 6634 24182 6686
rect 24118 6538 24124 6550
rect 24079 6510 24124 6538
rect 24118 6498 24124 6510
rect 24176 6498 24182 6550
rect 11054 6470 11060 6482
rect 11015 6442 11060 6470
rect 11054 6430 11060 6442
rect 11112 6430 11118 6482
rect 14826 6470 14832 6482
rect 14787 6442 14832 6470
rect 14826 6430 14832 6442
rect 14884 6430 14890 6482
rect 1104 6380 28888 6402
rect 1104 6328 5982 6380
rect 6034 6328 6046 6380
rect 6098 6328 6110 6380
rect 6162 6328 6174 6380
rect 6226 6328 15982 6380
rect 16034 6328 16046 6380
rect 16098 6328 16110 6380
rect 16162 6328 16174 6380
rect 16226 6328 25982 6380
rect 26034 6328 26046 6380
rect 26098 6328 26110 6380
rect 26162 6328 26174 6380
rect 26226 6328 28888 6380
rect 1104 6306 28888 6328
rect 10870 6266 10876 6278
rect 10831 6238 10876 6266
rect 10870 6226 10876 6238
rect 10928 6226 10934 6278
rect 14642 6266 14648 6278
rect 14603 6238 14648 6266
rect 14642 6226 14648 6238
rect 14700 6226 14706 6278
rect 23934 6266 23940 6278
rect 23895 6238 23940 6266
rect 23934 6226 23940 6238
rect 23992 6226 23998 6278
rect 1104 5836 28888 5858
rect 1104 5784 10982 5836
rect 11034 5784 11046 5836
rect 11098 5784 11110 5836
rect 11162 5784 11174 5836
rect 11226 5784 20982 5836
rect 21034 5784 21046 5836
rect 21098 5784 21110 5836
rect 21162 5784 21174 5836
rect 21226 5784 28888 5836
rect 1104 5762 28888 5784
rect 12802 5722 12808 5734
rect 12763 5694 12808 5722
rect 12802 5682 12808 5694
rect 12860 5682 12866 5734
rect 4798 5586 4804 5598
rect 4759 5558 4804 5586
rect 4798 5546 4804 5558
rect 4856 5546 4862 5598
rect 12618 5586 12624 5598
rect 12579 5558 12624 5586
rect 12618 5546 12624 5558
rect 12676 5546 12682 5598
rect 4982 5450 4988 5462
rect 4943 5422 4988 5450
rect 4982 5410 4988 5422
rect 5040 5410 5046 5462
rect 1104 5292 28888 5314
rect 1104 5240 5982 5292
rect 6034 5240 6046 5292
rect 6098 5240 6110 5292
rect 6162 5240 6174 5292
rect 6226 5240 15982 5292
rect 16034 5240 16046 5292
rect 16098 5240 16110 5292
rect 16162 5240 16174 5292
rect 16226 5240 25982 5292
rect 26034 5240 26046 5292
rect 26098 5240 26110 5292
rect 26162 5240 26174 5292
rect 26226 5240 28888 5292
rect 1104 5218 28888 5240
rect 4798 5178 4804 5190
rect 4759 5150 4804 5178
rect 4798 5138 4804 5150
rect 4856 5138 4862 5190
rect 12618 5178 12624 5190
rect 12579 5150 12624 5178
rect 12618 5138 12624 5150
rect 12676 5138 12682 5190
rect 13909 5181 13967 5187
rect 13909 5147 13921 5181
rect 13955 5178 13967 5181
rect 16390 5178 16396 5190
rect 13955 5150 16396 5178
rect 13955 5147 13967 5150
rect 13909 5141 13967 5147
rect 16390 5138 16396 5150
rect 16448 5138 16454 5190
rect 13722 4974 13728 4986
rect 13683 4946 13728 4974
rect 13722 4934 13728 4946
rect 13780 4974 13786 4986
rect 14277 4977 14335 4983
rect 14277 4974 14289 4977
rect 13780 4946 14289 4974
rect 13780 4934 13786 4946
rect 14277 4943 14289 4946
rect 14323 4943 14335 4977
rect 14277 4937 14335 4943
rect 23566 4934 23572 4986
rect 23624 4974 23630 4986
rect 23937 4977 23995 4983
rect 23937 4974 23949 4977
rect 23624 4946 23949 4974
rect 23624 4934 23630 4946
rect 23937 4943 23949 4946
rect 23983 4974 23995 4977
rect 24489 4977 24547 4983
rect 24489 4974 24501 4977
rect 23983 4946 24501 4974
rect 23983 4943 23995 4946
rect 23937 4937 23995 4943
rect 24489 4943 24501 4946
rect 24535 4943 24547 4977
rect 24489 4937 24547 4943
rect 24118 4838 24124 4850
rect 24079 4810 24124 4838
rect 24118 4798 24124 4810
rect 24176 4798 24182 4850
rect 1104 4748 28888 4770
rect 1104 4696 10982 4748
rect 11034 4696 11046 4748
rect 11098 4696 11110 4748
rect 11162 4696 11174 4748
rect 11226 4696 20982 4748
rect 21034 4696 21046 4748
rect 21098 4696 21110 4748
rect 21162 4696 21174 4748
rect 21226 4696 28888 4748
rect 1104 4674 28888 4696
rect 16301 4501 16359 4507
rect 16301 4467 16313 4501
rect 16347 4498 16359 4501
rect 16390 4498 16396 4510
rect 16347 4470 16396 4498
rect 16347 4467 16359 4470
rect 16301 4461 16359 4467
rect 16390 4458 16396 4470
rect 16448 4458 16454 4510
rect 20714 4498 20720 4510
rect 20675 4470 20720 4498
rect 20714 4458 20720 4470
rect 20772 4458 20778 4510
rect 16482 4362 16488 4374
rect 16443 4334 16488 4362
rect 16482 4322 16488 4334
rect 16540 4322 16546 4374
rect 20898 4362 20904 4374
rect 20859 4334 20904 4362
rect 20898 4322 20904 4334
rect 20956 4322 20962 4374
rect 1104 4204 28888 4226
rect 1104 4152 5982 4204
rect 6034 4152 6046 4204
rect 6098 4152 6110 4204
rect 6162 4152 6174 4204
rect 6226 4152 15982 4204
rect 16034 4152 16046 4204
rect 16098 4152 16110 4204
rect 16162 4152 16174 4204
rect 16226 4152 25982 4204
rect 26034 4152 26046 4204
rect 26098 4152 26110 4204
rect 26162 4152 26174 4204
rect 26226 4152 28888 4204
rect 1104 4130 28888 4152
rect 20714 4050 20720 4102
rect 20772 4090 20778 4102
rect 21085 4093 21143 4099
rect 21085 4090 21097 4093
rect 20772 4062 21097 4090
rect 20772 4050 20778 4062
rect 21085 4059 21097 4062
rect 21131 4059 21143 4093
rect 21085 4053 21143 4059
rect 16390 4022 16396 4034
rect 16351 3994 16396 4022
rect 16390 3982 16396 3994
rect 16448 3982 16454 4034
rect 21453 3889 21511 3895
rect 21453 3855 21465 3889
rect 21499 3886 21511 3889
rect 23934 3886 23940 3898
rect 21499 3858 22140 3886
rect 23895 3858 23940 3886
rect 21499 3855 21511 3858
rect 21453 3849 21511 3855
rect 22112 3762 22140 3858
rect 23934 3846 23940 3858
rect 23992 3886 23998 3898
rect 24489 3889 24547 3895
rect 24489 3886 24501 3889
rect 23992 3858 24501 3886
rect 23992 3846 23998 3858
rect 24489 3855 24501 3858
rect 24535 3855 24547 3889
rect 24489 3849 24547 3855
rect 21634 3750 21640 3762
rect 21595 3722 21640 3750
rect 21634 3710 21640 3722
rect 21692 3710 21698 3762
rect 22094 3750 22100 3762
rect 22055 3722 22100 3750
rect 22094 3710 22100 3722
rect 22152 3710 22158 3762
rect 24118 3750 24124 3762
rect 24079 3722 24124 3750
rect 24118 3710 24124 3722
rect 24176 3710 24182 3762
rect 1104 3660 28888 3682
rect 1104 3608 10982 3660
rect 11034 3608 11046 3660
rect 11098 3608 11110 3660
rect 11162 3608 11174 3660
rect 11226 3608 20982 3660
rect 21034 3608 21046 3660
rect 21098 3608 21110 3660
rect 21162 3608 21174 3660
rect 21226 3608 28888 3660
rect 1104 3586 28888 3608
rect 23937 3413 23995 3419
rect 23937 3379 23949 3413
rect 23983 3410 23995 3413
rect 24026 3410 24032 3422
rect 23983 3382 24032 3410
rect 23983 3379 23995 3382
rect 23937 3373 23995 3379
rect 24026 3370 24032 3382
rect 24084 3370 24090 3422
rect 24118 3274 24124 3286
rect 24079 3246 24124 3274
rect 24118 3234 24124 3246
rect 24176 3234 24182 3286
rect 1104 3116 28888 3138
rect 1104 3064 5982 3116
rect 6034 3064 6046 3116
rect 6098 3064 6110 3116
rect 6162 3064 6174 3116
rect 6226 3064 15982 3116
rect 16034 3064 16046 3116
rect 16098 3064 16110 3116
rect 16162 3064 16174 3116
rect 16226 3064 25982 3116
rect 26034 3064 26046 3116
rect 26098 3064 26110 3116
rect 26162 3064 26174 3116
rect 26226 3064 28888 3116
rect 1104 3042 28888 3064
rect 23845 3005 23903 3011
rect 23845 2971 23857 3005
rect 23891 3002 23903 3005
rect 24026 3002 24032 3014
rect 23891 2974 24032 3002
rect 23891 2971 23903 2974
rect 23845 2965 23903 2971
rect 24026 2962 24032 2974
rect 24084 2962 24090 3014
rect 1394 2798 1400 2810
rect 1355 2770 1400 2798
rect 1394 2758 1400 2770
rect 1452 2798 1458 2810
rect 1949 2801 2007 2807
rect 1949 2798 1961 2801
rect 1452 2770 1961 2798
rect 1452 2758 1458 2770
rect 1949 2767 1961 2770
rect 1995 2767 2007 2801
rect 23934 2798 23940 2810
rect 23895 2770 23940 2798
rect 1949 2761 2007 2767
rect 23934 2758 23940 2770
rect 23992 2798 23998 2810
rect 24489 2801 24547 2807
rect 24489 2798 24501 2801
rect 23992 2770 24501 2798
rect 23992 2758 23998 2770
rect 24489 2767 24501 2770
rect 24535 2767 24547 2801
rect 24489 2761 24547 2767
rect 1581 2665 1639 2671
rect 1581 2631 1593 2665
rect 1627 2662 1639 2665
rect 2682 2662 2688 2674
rect 1627 2634 2688 2662
rect 1627 2631 1639 2634
rect 1581 2625 1639 2631
rect 2682 2622 2688 2634
rect 2740 2622 2746 2674
rect 24121 2665 24179 2671
rect 24121 2631 24133 2665
rect 24167 2662 24179 2665
rect 24854 2662 24860 2674
rect 24167 2634 24860 2662
rect 24167 2631 24179 2634
rect 24121 2625 24179 2631
rect 24854 2622 24860 2634
rect 24912 2622 24918 2674
rect 1104 2572 28888 2594
rect 1104 2520 10982 2572
rect 11034 2520 11046 2572
rect 11098 2520 11110 2572
rect 11162 2520 11174 2572
rect 11226 2520 20982 2572
rect 21034 2520 21046 2572
rect 21098 2520 21110 2572
rect 21162 2520 21174 2572
rect 21226 2520 28888 2572
rect 1104 2498 28888 2520
rect 24210 2458 24216 2470
rect 24171 2430 24216 2458
rect 24210 2418 24216 2430
rect 24268 2418 24274 2470
rect 1397 2325 1455 2331
rect 1397 2291 1409 2325
rect 1443 2322 1455 2325
rect 2038 2322 2044 2334
rect 1443 2294 2044 2322
rect 1443 2291 1455 2294
rect 1397 2285 1455 2291
rect 2038 2282 2044 2294
rect 2096 2282 2102 2334
rect 24026 2322 24032 2334
rect 23987 2294 24032 2322
rect 24026 2282 24032 2294
rect 24084 2322 24090 2334
rect 24581 2325 24639 2331
rect 24581 2322 24593 2325
rect 24084 2294 24593 2322
rect 24084 2282 24090 2294
rect 24581 2291 24593 2294
rect 24627 2291 24639 2325
rect 25130 2322 25136 2334
rect 25091 2294 25136 2322
rect 24581 2285 24639 2291
rect 25130 2282 25136 2294
rect 25188 2322 25194 2334
rect 25685 2325 25743 2331
rect 25685 2322 25697 2325
rect 25188 2294 25697 2322
rect 25188 2282 25194 2294
rect 25685 2291 25697 2294
rect 25731 2291 25743 2325
rect 25685 2285 25743 2291
rect 1578 2118 1584 2130
rect 1539 2090 1584 2118
rect 1578 2078 1584 2090
rect 1636 2078 1642 2130
rect 25314 2118 25320 2130
rect 25275 2090 25320 2118
rect 25314 2078 25320 2090
rect 25372 2078 25378 2130
rect 1104 2028 28888 2050
rect 1104 1976 5982 2028
rect 6034 1976 6046 2028
rect 6098 1976 6110 2028
rect 6162 1976 6174 2028
rect 6226 1976 15982 2028
rect 16034 1976 16046 2028
rect 16098 1976 16110 2028
rect 16162 1976 16174 2028
rect 16226 1976 25982 2028
rect 26034 1976 26046 2028
rect 26098 1976 26110 2028
rect 26162 1976 26174 2028
rect 26226 1976 28888 2028
rect 1104 1954 28888 1976
<< via1 >>
rect 5982 21560 6034 21612
rect 6046 21560 6098 21612
rect 6110 21560 6162 21612
rect 6174 21560 6226 21612
rect 15982 21560 16034 21612
rect 16046 21560 16098 21612
rect 16110 21560 16162 21612
rect 16174 21560 16226 21612
rect 25982 21560 26034 21612
rect 26046 21560 26098 21612
rect 26110 21560 26162 21612
rect 26174 21560 26226 21612
rect 10982 21016 11034 21068
rect 11046 21016 11098 21068
rect 11110 21016 11162 21068
rect 11174 21016 11226 21068
rect 20982 21016 21034 21068
rect 21046 21016 21098 21068
rect 21110 21016 21162 21068
rect 21174 21016 21226 21068
rect 3424 20574 3476 20626
rect 19800 20574 19852 20626
rect 20168 20574 20220 20626
rect 24860 20574 24912 20626
rect 5982 20472 6034 20524
rect 6046 20472 6098 20524
rect 6110 20472 6162 20524
rect 6174 20472 6226 20524
rect 15982 20472 16034 20524
rect 16046 20472 16098 20524
rect 16110 20472 16162 20524
rect 16174 20472 16226 20524
rect 25982 20472 26034 20524
rect 26046 20472 26098 20524
rect 26110 20472 26162 20524
rect 26174 20472 26226 20524
rect 10982 19928 11034 19980
rect 11046 19928 11098 19980
rect 11110 19928 11162 19980
rect 11174 19928 11226 19980
rect 20982 19928 21034 19980
rect 21046 19928 21098 19980
rect 21110 19928 21162 19980
rect 21174 19928 21226 19980
rect 5982 19384 6034 19436
rect 6046 19384 6098 19436
rect 6110 19384 6162 19436
rect 6174 19384 6226 19436
rect 15982 19384 16034 19436
rect 16046 19384 16098 19436
rect 16110 19384 16162 19436
rect 16174 19384 16226 19436
rect 25982 19384 26034 19436
rect 26046 19384 26098 19436
rect 26110 19384 26162 19436
rect 26174 19384 26226 19436
rect 23940 19121 23992 19130
rect 23940 19087 23949 19121
rect 23949 19087 23983 19121
rect 23983 19087 23992 19121
rect 23940 19078 23992 19087
rect 24676 18942 24728 18994
rect 10982 18840 11034 18892
rect 11046 18840 11098 18892
rect 11110 18840 11162 18892
rect 11174 18840 11226 18892
rect 20982 18840 21034 18892
rect 21046 18840 21098 18892
rect 21110 18840 21162 18892
rect 21174 18840 21226 18892
rect 16672 18781 16724 18790
rect 16672 18747 16681 18781
rect 16681 18747 16715 18781
rect 16715 18747 16724 18781
rect 16672 18738 16724 18747
rect 20628 18781 20680 18790
rect 20628 18747 20637 18781
rect 20637 18747 20671 18781
rect 20671 18747 20680 18781
rect 20628 18738 20680 18747
rect 8852 18713 8904 18722
rect 8852 18679 8886 18713
rect 8886 18679 8904 18713
rect 8852 18670 8904 18679
rect 8576 18645 8628 18654
rect 8576 18611 8585 18645
rect 8585 18611 8619 18645
rect 8619 18611 8628 18645
rect 8576 18602 8628 18611
rect 15200 18602 15252 18654
rect 20444 18645 20496 18654
rect 20444 18611 20453 18645
rect 20453 18611 20487 18645
rect 20487 18611 20496 18645
rect 20444 18602 20496 18611
rect 23756 18602 23808 18654
rect 25044 18645 25096 18654
rect 25044 18611 25053 18645
rect 25053 18611 25087 18645
rect 25087 18611 25096 18645
rect 25044 18602 25096 18611
rect 15292 18577 15344 18586
rect 15292 18543 15301 18577
rect 15301 18543 15335 18577
rect 15335 18543 15344 18577
rect 15292 18534 15344 18543
rect 9956 18441 10008 18450
rect 9956 18407 9965 18441
rect 9965 18407 9999 18441
rect 9999 18407 10008 18441
rect 9956 18398 10008 18407
rect 24124 18441 24176 18450
rect 24124 18407 24133 18441
rect 24133 18407 24167 18441
rect 24167 18407 24176 18441
rect 24124 18398 24176 18407
rect 25320 18398 25372 18450
rect 5982 18296 6034 18348
rect 6046 18296 6098 18348
rect 6110 18296 6162 18348
rect 6174 18296 6226 18348
rect 15982 18296 16034 18348
rect 16046 18296 16098 18348
rect 16110 18296 16162 18348
rect 16174 18296 16226 18348
rect 25982 18296 26034 18348
rect 26046 18296 26098 18348
rect 26110 18296 26162 18348
rect 26174 18296 26226 18348
rect 8852 18194 8904 18246
rect 15292 18194 15344 18246
rect 25044 18237 25096 18246
rect 25044 18203 25053 18237
rect 25053 18203 25087 18237
rect 25087 18203 25096 18237
rect 25044 18194 25096 18203
rect 8576 18126 8628 18178
rect 23756 18169 23808 18178
rect 23756 18135 23765 18169
rect 23765 18135 23799 18169
rect 23799 18135 23808 18169
rect 23756 18126 23808 18135
rect 23940 18033 23992 18042
rect 23940 17999 23949 18033
rect 23949 17999 23983 18033
rect 23983 17999 23992 18033
rect 23940 17990 23992 17999
rect 15200 17922 15252 17974
rect 19340 17854 19392 17906
rect 20444 17897 20496 17906
rect 20444 17863 20453 17897
rect 20453 17863 20487 17897
rect 20487 17863 20496 17897
rect 20444 17854 20496 17863
rect 24216 17854 24268 17906
rect 10982 17752 11034 17804
rect 11046 17752 11098 17804
rect 11110 17752 11162 17804
rect 11174 17752 11226 17804
rect 20982 17752 21034 17804
rect 21046 17752 21098 17804
rect 21110 17752 21162 17804
rect 21174 17752 21226 17804
rect 24308 17514 24360 17566
rect 23480 17310 23532 17362
rect 5982 17208 6034 17260
rect 6046 17208 6098 17260
rect 6110 17208 6162 17260
rect 6174 17208 6226 17260
rect 15982 17208 16034 17260
rect 16046 17208 16098 17260
rect 16110 17208 16162 17260
rect 16174 17208 16226 17260
rect 25982 17208 26034 17260
rect 26046 17208 26098 17260
rect 26110 17208 26162 17260
rect 26174 17208 26226 17260
rect 19248 17106 19300 17158
rect 24308 17106 24360 17158
rect 18696 17013 18748 17022
rect 18696 16979 18705 17013
rect 18705 16979 18739 17013
rect 18739 16979 18748 17013
rect 18696 16970 18748 16979
rect 17500 16809 17552 16818
rect 17500 16775 17509 16809
rect 17509 16775 17543 16809
rect 17543 16775 17552 16809
rect 17500 16766 17552 16775
rect 18328 16766 18380 16818
rect 10982 16664 11034 16716
rect 11046 16664 11098 16716
rect 11110 16664 11162 16716
rect 11174 16664 11226 16716
rect 20982 16664 21034 16716
rect 21046 16664 21098 16716
rect 21110 16664 21162 16716
rect 21174 16664 21226 16716
rect 14188 16562 14240 16614
rect 15200 16562 15252 16614
rect 18328 16605 18380 16614
rect 18328 16571 18337 16605
rect 18337 16571 18371 16605
rect 18371 16571 18380 16605
rect 18328 16562 18380 16571
rect 12992 16469 13044 16478
rect 12992 16435 13001 16469
rect 13001 16435 13035 16469
rect 13035 16435 13044 16469
rect 12992 16426 13044 16435
rect 13728 16426 13780 16478
rect 5982 16120 6034 16172
rect 6046 16120 6098 16172
rect 6110 16120 6162 16172
rect 6174 16120 6226 16172
rect 15982 16120 16034 16172
rect 16046 16120 16098 16172
rect 16110 16120 16162 16172
rect 16174 16120 16226 16172
rect 25982 16120 26034 16172
rect 26046 16120 26098 16172
rect 26110 16120 26162 16172
rect 26174 16120 26226 16172
rect 7012 16061 7064 16070
rect 7012 16027 7021 16061
rect 7021 16027 7055 16061
rect 7055 16027 7064 16061
rect 7012 16018 7064 16027
rect 12992 16061 13044 16070
rect 12992 16027 13001 16061
rect 13001 16027 13035 16061
rect 13035 16027 13044 16061
rect 12992 16018 13044 16027
rect 24492 16061 24544 16070
rect 24492 16027 24501 16061
rect 24501 16027 24535 16061
rect 24535 16027 24544 16061
rect 24492 16018 24544 16027
rect 24492 15814 24544 15866
rect 7196 15746 7248 15798
rect 8576 15678 8628 15730
rect 13728 15678 13780 15730
rect 23664 15678 23716 15730
rect 10982 15576 11034 15628
rect 11046 15576 11098 15628
rect 11110 15576 11162 15628
rect 11174 15576 11226 15628
rect 20982 15576 21034 15628
rect 21046 15576 21098 15628
rect 21110 15576 21162 15628
rect 21174 15576 21226 15628
rect 7196 15517 7248 15526
rect 7196 15483 7205 15517
rect 7205 15483 7239 15517
rect 7239 15483 7248 15517
rect 7196 15474 7248 15483
rect 24032 15338 24084 15390
rect 24768 15338 24820 15390
rect 18604 15177 18656 15186
rect 18604 15143 18613 15177
rect 18613 15143 18647 15177
rect 18647 15143 18656 15177
rect 18604 15134 18656 15143
rect 23756 15134 23808 15186
rect 5982 15032 6034 15084
rect 6046 15032 6098 15084
rect 6110 15032 6162 15084
rect 6174 15032 6226 15084
rect 15982 15032 16034 15084
rect 16046 15032 16098 15084
rect 16110 15032 16162 15084
rect 16174 15032 16226 15084
rect 25982 15032 26034 15084
rect 26046 15032 26098 15084
rect 26110 15032 26162 15084
rect 26174 15032 26226 15084
rect 18328 14930 18380 14982
rect 24032 14973 24084 14982
rect 24032 14939 24041 14973
rect 24041 14939 24075 14973
rect 24075 14939 24084 14973
rect 24032 14930 24084 14939
rect 18328 14837 18380 14846
rect 18328 14803 18337 14837
rect 18337 14803 18371 14837
rect 18371 14803 18380 14837
rect 18328 14794 18380 14803
rect 18604 14658 18656 14710
rect 19248 14658 19300 14710
rect 18972 14633 19024 14642
rect 18972 14599 18981 14633
rect 18981 14599 19015 14633
rect 19015 14599 19024 14633
rect 18972 14590 19024 14599
rect 10982 14488 11034 14540
rect 11046 14488 11098 14540
rect 11110 14488 11162 14540
rect 11174 14488 11226 14540
rect 20982 14488 21034 14540
rect 21046 14488 21098 14540
rect 21110 14488 21162 14540
rect 21174 14488 21226 14540
rect 18972 14386 19024 14438
rect 19616 14250 19668 14302
rect 19800 14293 19852 14302
rect 19800 14259 19809 14293
rect 19809 14259 19843 14293
rect 19843 14259 19852 14293
rect 19800 14250 19852 14259
rect 19892 14225 19944 14234
rect 19892 14191 19901 14225
rect 19901 14191 19935 14225
rect 19935 14191 19944 14225
rect 19892 14182 19944 14191
rect 20444 14182 20496 14234
rect 5982 13944 6034 13996
rect 6046 13944 6098 13996
rect 6110 13944 6162 13996
rect 6174 13944 6226 13996
rect 15982 13944 16034 13996
rect 16046 13944 16098 13996
rect 16110 13944 16162 13996
rect 16174 13944 16226 13996
rect 25982 13944 26034 13996
rect 26046 13944 26098 13996
rect 26110 13944 26162 13996
rect 26174 13944 26226 13996
rect 24860 13842 24912 13894
rect 25320 13842 25372 13894
rect 19616 13681 19668 13690
rect 19616 13647 19625 13681
rect 19625 13647 19659 13681
rect 19659 13647 19668 13681
rect 19616 13638 19668 13647
rect 19892 13681 19944 13690
rect 19892 13647 19901 13681
rect 19901 13647 19935 13681
rect 19935 13647 19944 13681
rect 19892 13638 19944 13647
rect 24216 13638 24268 13690
rect 24768 13638 24820 13690
rect 19064 13545 19116 13554
rect 19064 13511 19073 13545
rect 19073 13511 19107 13545
rect 19107 13511 19116 13545
rect 19064 13502 19116 13511
rect 20444 13502 20496 13554
rect 10982 13400 11034 13452
rect 11046 13400 11098 13452
rect 11110 13400 11162 13452
rect 11174 13400 11226 13452
rect 20982 13400 21034 13452
rect 21046 13400 21098 13452
rect 21110 13400 21162 13452
rect 21174 13400 21226 13452
rect 13544 13341 13596 13350
rect 13544 13307 13553 13341
rect 13553 13307 13587 13341
rect 13587 13307 13596 13341
rect 13544 13298 13596 13307
rect 19064 13298 19116 13350
rect 20076 13341 20128 13350
rect 20076 13307 20085 13341
rect 20085 13307 20119 13341
rect 20119 13307 20128 13341
rect 20076 13298 20128 13307
rect 1492 13162 1544 13214
rect 13912 13205 13964 13214
rect 13912 13171 13921 13205
rect 13921 13171 13955 13205
rect 13955 13171 13964 13205
rect 13912 13162 13964 13171
rect 19708 13162 19760 13214
rect 20168 13205 20220 13214
rect 20168 13171 20177 13205
rect 20177 13171 20211 13205
rect 20211 13171 20220 13205
rect 20168 13162 20220 13171
rect 13820 13094 13872 13146
rect 14188 13137 14240 13146
rect 14188 13103 14197 13137
rect 14197 13103 14231 13137
rect 14231 13103 14240 13137
rect 14188 13094 14240 13103
rect 20444 13094 20496 13146
rect 19340 13026 19392 13078
rect 2136 12958 2188 13010
rect 13084 13001 13136 13010
rect 13084 12967 13093 13001
rect 13093 12967 13127 13001
rect 13127 12967 13136 13001
rect 13084 12958 13136 12967
rect 5982 12856 6034 12908
rect 6046 12856 6098 12908
rect 6110 12856 6162 12908
rect 6174 12856 6226 12908
rect 15982 12856 16034 12908
rect 16046 12856 16098 12908
rect 16110 12856 16162 12908
rect 16174 12856 16226 12908
rect 25982 12856 26034 12908
rect 26046 12856 26098 12908
rect 26110 12856 26162 12908
rect 26174 12856 26226 12908
rect 14188 12797 14240 12806
rect 14188 12763 14197 12797
rect 14197 12763 14231 12797
rect 14231 12763 14240 12797
rect 14188 12754 14240 12763
rect 20076 12797 20128 12806
rect 20076 12763 20085 12797
rect 20085 12763 20119 12797
rect 20119 12763 20128 12797
rect 20076 12754 20128 12763
rect 13912 12686 13964 12738
rect 13728 12661 13780 12670
rect 13728 12627 13737 12661
rect 13737 12627 13771 12661
rect 13771 12627 13780 12661
rect 13728 12618 13780 12627
rect 1400 12593 1452 12602
rect 1400 12559 1409 12593
rect 1409 12559 1443 12593
rect 1443 12559 1452 12593
rect 1400 12550 1452 12559
rect 12900 12593 12952 12602
rect 12900 12559 12909 12593
rect 12909 12559 12943 12593
rect 12943 12559 12952 12593
rect 12900 12550 12952 12559
rect 12440 12482 12492 12534
rect 13084 12482 13136 12534
rect 1492 12414 1544 12466
rect 19708 12457 19760 12466
rect 19708 12423 19717 12457
rect 19717 12423 19751 12457
rect 19751 12423 19760 12457
rect 19708 12414 19760 12423
rect 20444 12457 20496 12466
rect 20444 12423 20453 12457
rect 20453 12423 20487 12457
rect 20487 12423 20496 12457
rect 20444 12414 20496 12423
rect 10982 12312 11034 12364
rect 11046 12312 11098 12364
rect 11110 12312 11162 12364
rect 11174 12312 11226 12364
rect 20982 12312 21034 12364
rect 21046 12312 21098 12364
rect 21110 12312 21162 12364
rect 21174 12312 21226 12364
rect 1584 12253 1636 12262
rect 1584 12219 1593 12253
rect 1593 12219 1627 12253
rect 1627 12219 1636 12253
rect 1584 12210 1636 12219
rect 3608 12210 3660 12262
rect 3884 12210 3936 12262
rect 13912 12253 13964 12262
rect 13912 12219 13921 12253
rect 13921 12219 13955 12253
rect 13955 12219 13964 12253
rect 13912 12210 13964 12219
rect 13728 12142 13780 12194
rect 8668 12074 8720 12126
rect 8576 12049 8628 12058
rect 7932 11981 7984 11990
rect 7932 11947 7941 11981
rect 7941 11947 7975 11981
rect 7975 11947 7984 11981
rect 7932 11938 7984 11947
rect 8300 11938 8352 11990
rect 8576 12015 8585 12049
rect 8585 12015 8619 12049
rect 8619 12015 8628 12049
rect 8576 12006 8628 12015
rect 13728 11938 13780 11990
rect 12072 11913 12124 11922
rect 12072 11879 12081 11913
rect 12081 11879 12115 11913
rect 12115 11879 12124 11913
rect 12072 11870 12124 11879
rect 5982 11768 6034 11820
rect 6046 11768 6098 11820
rect 6110 11768 6162 11820
rect 6174 11768 6226 11820
rect 15982 11768 16034 11820
rect 16046 11768 16098 11820
rect 16110 11768 16162 11820
rect 16174 11768 16226 11820
rect 25982 11768 26034 11820
rect 26046 11768 26098 11820
rect 26110 11768 26162 11820
rect 26174 11768 26226 11820
rect 8576 11666 8628 11718
rect 11888 11709 11940 11718
rect 11888 11675 11897 11709
rect 11897 11675 11931 11709
rect 11931 11675 11940 11709
rect 11888 11666 11940 11675
rect 12348 11666 12400 11718
rect 24860 11598 24912 11650
rect 12072 11530 12124 11582
rect 1676 11462 1728 11514
rect 11888 11462 11940 11514
rect 12532 11462 12584 11514
rect 23480 11462 23532 11514
rect 11520 11394 11572 11446
rect 13728 11394 13780 11446
rect 2228 11326 2280 11378
rect 8300 11369 8352 11378
rect 8300 11335 8309 11369
rect 8309 11335 8343 11369
rect 8343 11335 8352 11369
rect 8300 11326 8352 11335
rect 8668 11369 8720 11378
rect 8668 11335 8677 11369
rect 8677 11335 8711 11369
rect 8711 11335 8720 11369
rect 8668 11326 8720 11335
rect 12532 11369 12584 11378
rect 12532 11335 12541 11369
rect 12541 11335 12575 11369
rect 12575 11335 12584 11369
rect 12532 11326 12584 11335
rect 10982 11224 11034 11276
rect 11046 11224 11098 11276
rect 11110 11224 11162 11276
rect 11174 11224 11226 11276
rect 20982 11224 21034 11276
rect 21046 11224 21098 11276
rect 21110 11224 21162 11276
rect 21174 11224 21226 11276
rect 8668 11122 8720 11174
rect 11520 11122 11572 11174
rect 7196 11054 7248 11106
rect 2044 10986 2096 11038
rect 8116 11029 8168 11038
rect 8116 10995 8125 11029
rect 8125 10995 8159 11029
rect 8159 10995 8168 11029
rect 8116 10986 8168 10995
rect 24032 10986 24084 11038
rect 24400 10986 24452 11038
rect 7380 10918 7432 10970
rect 8392 10961 8444 10970
rect 8392 10927 8401 10961
rect 8401 10927 8435 10961
rect 8435 10927 8444 10961
rect 8392 10918 8444 10927
rect 1952 10850 2004 10902
rect 24124 10893 24176 10902
rect 24124 10859 24133 10893
rect 24133 10859 24167 10893
rect 24167 10859 24176 10893
rect 24124 10850 24176 10859
rect 5982 10680 6034 10732
rect 6046 10680 6098 10732
rect 6110 10680 6162 10732
rect 6174 10680 6226 10732
rect 15982 10680 16034 10732
rect 16046 10680 16098 10732
rect 16110 10680 16162 10732
rect 16174 10680 16226 10732
rect 25982 10680 26034 10732
rect 26046 10680 26098 10732
rect 26110 10680 26162 10732
rect 26174 10680 26226 10732
rect 2044 10621 2096 10630
rect 2044 10587 2053 10621
rect 2053 10587 2087 10621
rect 2087 10587 2096 10621
rect 2044 10578 2096 10587
rect 2412 10621 2464 10630
rect 2412 10587 2421 10621
rect 2421 10587 2455 10621
rect 2455 10587 2464 10621
rect 2412 10578 2464 10587
rect 8208 10578 8260 10630
rect 8392 10578 8444 10630
rect 7104 10553 7156 10562
rect 7104 10519 7113 10553
rect 7113 10519 7147 10553
rect 7147 10519 7156 10553
rect 7104 10510 7156 10519
rect 8116 10510 8168 10562
rect 24032 10621 24084 10630
rect 24032 10587 24041 10621
rect 24041 10587 24075 10621
rect 24075 10587 24084 10621
rect 24032 10578 24084 10587
rect 2412 10374 2464 10426
rect 8300 10349 8352 10358
rect 8300 10315 8309 10349
rect 8309 10315 8343 10349
rect 8343 10315 8352 10349
rect 8300 10306 8352 10315
rect 1768 10238 1820 10290
rect 7380 10281 7432 10290
rect 7380 10247 7389 10281
rect 7389 10247 7423 10281
rect 7423 10247 7432 10281
rect 7380 10238 7432 10247
rect 7840 10281 7892 10290
rect 7840 10247 7849 10281
rect 7849 10247 7883 10281
rect 7883 10247 7892 10281
rect 8392 10281 8444 10290
rect 7840 10238 7892 10247
rect 8392 10247 8401 10281
rect 8401 10247 8435 10281
rect 8435 10247 8444 10281
rect 8392 10238 8444 10247
rect 10982 10136 11034 10188
rect 11046 10136 11098 10188
rect 11110 10136 11162 10188
rect 11174 10136 11226 10188
rect 20982 10136 21034 10188
rect 21046 10136 21098 10188
rect 21110 10136 21162 10188
rect 21174 10136 21226 10188
rect 8300 10034 8352 10086
rect 8484 10034 8536 10086
rect 2044 9898 2096 9950
rect 1584 9737 1636 9746
rect 1584 9703 1593 9737
rect 1593 9703 1627 9737
rect 1627 9703 1636 9737
rect 1584 9694 1636 9703
rect 5982 9592 6034 9644
rect 6046 9592 6098 9644
rect 6110 9592 6162 9644
rect 6174 9592 6226 9644
rect 15982 9592 16034 9644
rect 16046 9592 16098 9644
rect 16110 9592 16162 9644
rect 16174 9592 16226 9644
rect 25982 9592 26034 9644
rect 26046 9592 26098 9644
rect 26110 9592 26162 9644
rect 26174 9592 26226 9644
rect 2044 9533 2096 9542
rect 2044 9499 2053 9533
rect 2053 9499 2087 9533
rect 2087 9499 2096 9533
rect 2044 9490 2096 9499
rect 2504 9422 2556 9474
rect 23940 9329 23992 9338
rect 23940 9295 23949 9329
rect 23949 9295 23983 9329
rect 23983 9295 23992 9329
rect 23940 9286 23992 9295
rect 1676 9150 1728 9202
rect 24124 9193 24176 9202
rect 24124 9159 24133 9193
rect 24133 9159 24167 9193
rect 24167 9159 24176 9193
rect 24124 9150 24176 9159
rect 10982 9048 11034 9100
rect 11046 9048 11098 9100
rect 11110 9048 11162 9100
rect 11174 9048 11226 9100
rect 20982 9048 21034 9100
rect 21046 9048 21098 9100
rect 21110 9048 21162 9100
rect 21174 9048 21226 9100
rect 1400 8853 1452 8862
rect 1400 8819 1409 8853
rect 1409 8819 1443 8853
rect 1443 8819 1452 8853
rect 1400 8810 1452 8819
rect 24492 8810 24544 8862
rect 1492 8606 1544 8658
rect 24124 8649 24176 8658
rect 24124 8615 24133 8649
rect 24133 8615 24167 8649
rect 24167 8615 24176 8649
rect 24124 8606 24176 8615
rect 5982 8504 6034 8556
rect 6046 8504 6098 8556
rect 6110 8504 6162 8556
rect 6174 8504 6226 8556
rect 15982 8504 16034 8556
rect 16046 8504 16098 8556
rect 16110 8504 16162 8556
rect 16174 8504 16226 8556
rect 25982 8504 26034 8556
rect 26046 8504 26098 8556
rect 26110 8504 26162 8556
rect 26174 8504 26226 8556
rect 1400 8402 1452 8454
rect 23480 8334 23532 8386
rect 1400 8266 1452 8318
rect 1860 8266 1912 8318
rect 24584 8402 24636 8454
rect 24492 8241 24544 8250
rect 24492 8207 24501 8241
rect 24501 8207 24535 8241
rect 24535 8207 24544 8241
rect 24492 8198 24544 8207
rect 10784 8062 10836 8114
rect 11336 8062 11388 8114
rect 10982 7960 11034 8012
rect 11046 7960 11098 8012
rect 11110 7960 11162 8012
rect 11174 7960 11226 8012
rect 20982 7960 21034 8012
rect 21046 7960 21098 8012
rect 21110 7960 21162 8012
rect 21174 7960 21226 8012
rect 24124 7901 24176 7910
rect 24124 7867 24133 7901
rect 24133 7867 24167 7901
rect 24167 7867 24176 7901
rect 24124 7858 24176 7867
rect 23940 7765 23992 7774
rect 23940 7731 23949 7765
rect 23949 7731 23983 7765
rect 23983 7731 23992 7765
rect 23940 7722 23992 7731
rect 5982 7416 6034 7468
rect 6046 7416 6098 7468
rect 6110 7416 6162 7468
rect 6174 7416 6226 7468
rect 15982 7416 16034 7468
rect 16046 7416 16098 7468
rect 16110 7416 16162 7468
rect 16174 7416 16226 7468
rect 25982 7416 26034 7468
rect 26046 7416 26098 7468
rect 26110 7416 26162 7468
rect 26174 7416 26226 7468
rect 22652 7357 22704 7366
rect 22652 7323 22661 7357
rect 22661 7323 22695 7357
rect 22695 7323 22704 7357
rect 22652 7314 22704 7323
rect 23112 7357 23164 7366
rect 23112 7323 23121 7357
rect 23121 7323 23155 7357
rect 23155 7323 23164 7357
rect 23112 7314 23164 7323
rect 18880 7289 18932 7298
rect 18880 7255 18889 7289
rect 18889 7255 18923 7289
rect 18923 7255 18932 7289
rect 18880 7246 18932 7255
rect 18696 7153 18748 7162
rect 18696 7119 18705 7153
rect 18705 7119 18739 7153
rect 18739 7119 18748 7153
rect 18696 7110 18748 7119
rect 23112 7110 23164 7162
rect 23940 7153 23992 7162
rect 23940 7119 23949 7153
rect 23949 7119 23983 7153
rect 23983 7119 23992 7153
rect 23940 7110 23992 7119
rect 10982 6872 11034 6924
rect 11046 6872 11098 6924
rect 11110 6872 11162 6924
rect 11174 6872 11226 6924
rect 20982 6872 21034 6924
rect 21046 6872 21098 6924
rect 21110 6872 21162 6924
rect 21174 6872 21226 6924
rect 1584 6634 1636 6686
rect 1860 6634 1912 6686
rect 10876 6677 10928 6686
rect 10876 6643 10885 6677
rect 10885 6643 10919 6677
rect 10919 6643 10928 6677
rect 10876 6634 10928 6643
rect 14648 6677 14700 6686
rect 14648 6643 14657 6677
rect 14657 6643 14691 6677
rect 14691 6643 14700 6677
rect 14648 6634 14700 6643
rect 23940 6677 23992 6686
rect 23940 6643 23949 6677
rect 23949 6643 23983 6677
rect 23983 6643 23992 6677
rect 23940 6634 23992 6643
rect 24124 6634 24176 6686
rect 24124 6541 24176 6550
rect 24124 6507 24133 6541
rect 24133 6507 24167 6541
rect 24167 6507 24176 6541
rect 24124 6498 24176 6507
rect 11060 6473 11112 6482
rect 11060 6439 11069 6473
rect 11069 6439 11103 6473
rect 11103 6439 11112 6473
rect 11060 6430 11112 6439
rect 14832 6473 14884 6482
rect 14832 6439 14841 6473
rect 14841 6439 14875 6473
rect 14875 6439 14884 6473
rect 14832 6430 14884 6439
rect 5982 6328 6034 6380
rect 6046 6328 6098 6380
rect 6110 6328 6162 6380
rect 6174 6328 6226 6380
rect 15982 6328 16034 6380
rect 16046 6328 16098 6380
rect 16110 6328 16162 6380
rect 16174 6328 16226 6380
rect 25982 6328 26034 6380
rect 26046 6328 26098 6380
rect 26110 6328 26162 6380
rect 26174 6328 26226 6380
rect 10876 6269 10928 6278
rect 10876 6235 10885 6269
rect 10885 6235 10919 6269
rect 10919 6235 10928 6269
rect 10876 6226 10928 6235
rect 14648 6269 14700 6278
rect 14648 6235 14657 6269
rect 14657 6235 14691 6269
rect 14691 6235 14700 6269
rect 14648 6226 14700 6235
rect 23940 6269 23992 6278
rect 23940 6235 23949 6269
rect 23949 6235 23983 6269
rect 23983 6235 23992 6269
rect 23940 6226 23992 6235
rect 10982 5784 11034 5836
rect 11046 5784 11098 5836
rect 11110 5784 11162 5836
rect 11174 5784 11226 5836
rect 20982 5784 21034 5836
rect 21046 5784 21098 5836
rect 21110 5784 21162 5836
rect 21174 5784 21226 5836
rect 12808 5725 12860 5734
rect 12808 5691 12817 5725
rect 12817 5691 12851 5725
rect 12851 5691 12860 5725
rect 12808 5682 12860 5691
rect 4804 5589 4856 5598
rect 4804 5555 4813 5589
rect 4813 5555 4847 5589
rect 4847 5555 4856 5589
rect 4804 5546 4856 5555
rect 12624 5589 12676 5598
rect 12624 5555 12633 5589
rect 12633 5555 12667 5589
rect 12667 5555 12676 5589
rect 12624 5546 12676 5555
rect 4988 5453 5040 5462
rect 4988 5419 4997 5453
rect 4997 5419 5031 5453
rect 5031 5419 5040 5453
rect 4988 5410 5040 5419
rect 5982 5240 6034 5292
rect 6046 5240 6098 5292
rect 6110 5240 6162 5292
rect 6174 5240 6226 5292
rect 15982 5240 16034 5292
rect 16046 5240 16098 5292
rect 16110 5240 16162 5292
rect 16174 5240 16226 5292
rect 25982 5240 26034 5292
rect 26046 5240 26098 5292
rect 26110 5240 26162 5292
rect 26174 5240 26226 5292
rect 4804 5181 4856 5190
rect 4804 5147 4813 5181
rect 4813 5147 4847 5181
rect 4847 5147 4856 5181
rect 4804 5138 4856 5147
rect 12624 5181 12676 5190
rect 12624 5147 12633 5181
rect 12633 5147 12667 5181
rect 12667 5147 12676 5181
rect 12624 5138 12676 5147
rect 16396 5138 16448 5190
rect 13728 4977 13780 4986
rect 13728 4943 13737 4977
rect 13737 4943 13771 4977
rect 13771 4943 13780 4977
rect 13728 4934 13780 4943
rect 23572 4934 23624 4986
rect 24124 4841 24176 4850
rect 24124 4807 24133 4841
rect 24133 4807 24167 4841
rect 24167 4807 24176 4841
rect 24124 4798 24176 4807
rect 10982 4696 11034 4748
rect 11046 4696 11098 4748
rect 11110 4696 11162 4748
rect 11174 4696 11226 4748
rect 20982 4696 21034 4748
rect 21046 4696 21098 4748
rect 21110 4696 21162 4748
rect 21174 4696 21226 4748
rect 16396 4458 16448 4510
rect 20720 4501 20772 4510
rect 20720 4467 20729 4501
rect 20729 4467 20763 4501
rect 20763 4467 20772 4501
rect 20720 4458 20772 4467
rect 16488 4365 16540 4374
rect 16488 4331 16497 4365
rect 16497 4331 16531 4365
rect 16531 4331 16540 4365
rect 16488 4322 16540 4331
rect 20904 4365 20956 4374
rect 20904 4331 20913 4365
rect 20913 4331 20947 4365
rect 20947 4331 20956 4365
rect 20904 4322 20956 4331
rect 5982 4152 6034 4204
rect 6046 4152 6098 4204
rect 6110 4152 6162 4204
rect 6174 4152 6226 4204
rect 15982 4152 16034 4204
rect 16046 4152 16098 4204
rect 16110 4152 16162 4204
rect 16174 4152 16226 4204
rect 25982 4152 26034 4204
rect 26046 4152 26098 4204
rect 26110 4152 26162 4204
rect 26174 4152 26226 4204
rect 20720 4050 20772 4102
rect 16396 4025 16448 4034
rect 16396 3991 16405 4025
rect 16405 3991 16439 4025
rect 16439 3991 16448 4025
rect 16396 3982 16448 3991
rect 23940 3889 23992 3898
rect 23940 3855 23949 3889
rect 23949 3855 23983 3889
rect 23983 3855 23992 3889
rect 23940 3846 23992 3855
rect 21640 3753 21692 3762
rect 21640 3719 21649 3753
rect 21649 3719 21683 3753
rect 21683 3719 21692 3753
rect 21640 3710 21692 3719
rect 22100 3753 22152 3762
rect 22100 3719 22109 3753
rect 22109 3719 22143 3753
rect 22143 3719 22152 3753
rect 22100 3710 22152 3719
rect 24124 3753 24176 3762
rect 24124 3719 24133 3753
rect 24133 3719 24167 3753
rect 24167 3719 24176 3753
rect 24124 3710 24176 3719
rect 10982 3608 11034 3660
rect 11046 3608 11098 3660
rect 11110 3608 11162 3660
rect 11174 3608 11226 3660
rect 20982 3608 21034 3660
rect 21046 3608 21098 3660
rect 21110 3608 21162 3660
rect 21174 3608 21226 3660
rect 24032 3370 24084 3422
rect 24124 3277 24176 3286
rect 24124 3243 24133 3277
rect 24133 3243 24167 3277
rect 24167 3243 24176 3277
rect 24124 3234 24176 3243
rect 5982 3064 6034 3116
rect 6046 3064 6098 3116
rect 6110 3064 6162 3116
rect 6174 3064 6226 3116
rect 15982 3064 16034 3116
rect 16046 3064 16098 3116
rect 16110 3064 16162 3116
rect 16174 3064 16226 3116
rect 25982 3064 26034 3116
rect 26046 3064 26098 3116
rect 26110 3064 26162 3116
rect 26174 3064 26226 3116
rect 24032 2962 24084 3014
rect 1400 2801 1452 2810
rect 1400 2767 1409 2801
rect 1409 2767 1443 2801
rect 1443 2767 1452 2801
rect 1400 2758 1452 2767
rect 23940 2801 23992 2810
rect 23940 2767 23949 2801
rect 23949 2767 23983 2801
rect 23983 2767 23992 2801
rect 23940 2758 23992 2767
rect 2688 2622 2740 2674
rect 24860 2622 24912 2674
rect 10982 2520 11034 2572
rect 11046 2520 11098 2572
rect 11110 2520 11162 2572
rect 11174 2520 11226 2572
rect 20982 2520 21034 2572
rect 21046 2520 21098 2572
rect 21110 2520 21162 2572
rect 21174 2520 21226 2572
rect 24216 2461 24268 2470
rect 24216 2427 24225 2461
rect 24225 2427 24259 2461
rect 24259 2427 24268 2461
rect 24216 2418 24268 2427
rect 2044 2325 2096 2334
rect 2044 2291 2053 2325
rect 2053 2291 2087 2325
rect 2087 2291 2096 2325
rect 2044 2282 2096 2291
rect 24032 2325 24084 2334
rect 24032 2291 24041 2325
rect 24041 2291 24075 2325
rect 24075 2291 24084 2325
rect 24032 2282 24084 2291
rect 25136 2325 25188 2334
rect 25136 2291 25145 2325
rect 25145 2291 25179 2325
rect 25179 2291 25188 2325
rect 25136 2282 25188 2291
rect 1584 2121 1636 2130
rect 1584 2087 1593 2121
rect 1593 2087 1627 2121
rect 1627 2087 1636 2121
rect 1584 2078 1636 2087
rect 25320 2121 25372 2130
rect 25320 2087 25329 2121
rect 25329 2087 25363 2121
rect 25363 2087 25372 2121
rect 25320 2078 25372 2087
rect 5982 1976 6034 2028
rect 6046 1976 6098 2028
rect 6110 1976 6162 2028
rect 6174 1976 6226 2028
rect 15982 1976 16034 2028
rect 16046 1976 16098 2028
rect 16110 1976 16162 2028
rect 16174 1976 16226 2028
rect 25982 1976 26034 2028
rect 26046 1976 26098 2028
rect 26110 1976 26162 2028
rect 26174 1976 26226 2028
<< metal2 >>
rect 3698 23346 3754 23826
rect 3882 23450 3938 23459
rect 3882 23385 3938 23394
rect 3054 22906 3110 22915
rect 3054 22841 3110 22850
rect 3068 18019 3096 22841
rect 3330 22226 3386 22235
rect 3330 22161 3386 22170
rect 3344 19107 3372 22161
rect 3422 21682 3478 21691
rect 3422 21617 3478 21626
rect 3436 20632 3464 21617
rect 3514 21138 3570 21147
rect 3514 21073 3570 21082
rect 3424 20626 3476 20632
rect 3424 20568 3476 20574
rect 3422 19234 3478 19243
rect 3422 19169 3478 19178
rect 3330 19098 3386 19107
rect 3330 19033 3386 19042
rect 3146 18690 3202 18699
rect 3146 18625 3202 18634
rect 3054 18010 3110 18019
rect 3054 17945 3110 17954
rect 2962 15698 3018 15707
rect 2962 15633 3018 15642
rect 1398 15154 1454 15163
rect 1398 15089 1454 15098
rect 1412 12608 1440 15089
rect 1674 13930 1730 13939
rect 1674 13865 1730 13874
rect 1490 13250 1546 13259
rect 1490 13185 1492 13194
rect 1544 13185 1546 13194
rect 1492 13156 1544 13162
rect 1504 12828 1532 13156
rect 1504 12800 1624 12828
rect 1400 12602 1452 12608
rect 1400 12544 1452 12550
rect 1492 12466 1544 12472
rect 1492 12408 1544 12414
rect 1398 9986 1454 9995
rect 1398 9921 1454 9930
rect 1412 8868 1440 9921
rect 1504 9564 1532 12408
rect 1596 12268 1624 12800
rect 1584 12262 1636 12268
rect 1584 12204 1636 12210
rect 1688 11520 1716 13865
rect 2136 13010 2188 13016
rect 2136 12952 2188 12958
rect 1858 12706 1914 12715
rect 1858 12641 1914 12650
rect 1676 11514 1728 11520
rect 1676 11456 1728 11462
rect 1768 10290 1820 10296
rect 1768 10232 1820 10238
rect 1584 9746 1636 9752
rect 1582 9714 1584 9723
rect 1636 9714 1638 9723
rect 1582 9649 1638 9658
rect 1504 9536 1624 9564
rect 1400 8862 1452 8868
rect 1400 8804 1452 8810
rect 1412 8460 1440 8804
rect 1492 8658 1544 8664
rect 1492 8600 1544 8606
rect 1400 8454 1452 8460
rect 1400 8396 1452 8402
rect 1400 8318 1452 8324
rect 1400 8260 1452 8266
rect 1412 2816 1440 8260
rect 1400 2810 1452 2816
rect 1400 2752 1452 2758
rect 1504 203 1532 8600
rect 1596 6692 1624 9536
rect 1676 9202 1728 9208
rect 1676 9144 1728 9150
rect 1584 6686 1636 6692
rect 1584 6628 1636 6634
rect 1584 2130 1636 2136
rect 1584 2072 1636 2078
rect 1596 747 1624 2072
rect 1688 1291 1716 9144
rect 1780 2515 1808 10232
rect 1872 8324 1900 12641
rect 2042 11074 2098 11083
rect 2042 11009 2044 11018
rect 2096 11009 2098 11018
rect 2044 10980 2096 10986
rect 1952 10902 2004 10908
rect 1952 10844 2004 10850
rect 1964 8748 1992 10844
rect 2056 10636 2084 10980
rect 2044 10630 2096 10636
rect 2044 10572 2096 10578
rect 2044 9950 2096 9956
rect 2044 9892 2096 9898
rect 2056 9859 2084 9892
rect 2042 9850 2098 9859
rect 2042 9785 2098 9794
rect 2056 9548 2084 9785
rect 2044 9542 2096 9548
rect 2044 9484 2096 9490
rect 1964 8720 2084 8748
rect 1860 8318 1912 8324
rect 1860 8260 1912 8266
rect 1860 6686 1912 6692
rect 1860 6628 1912 6634
rect 1872 2787 1900 6628
rect 2056 4124 2084 8720
rect 2148 6187 2176 12952
rect 2228 11378 2280 11384
rect 2228 11320 2280 11326
rect 2410 11346 2466 11355
rect 2134 6178 2190 6187
rect 2134 6113 2190 6122
rect 1964 4096 2084 4124
rect 1858 2778 1914 2787
rect 1858 2713 1914 2722
rect 1766 2506 1822 2515
rect 1766 2441 1822 2450
rect 1964 1971 1992 4096
rect 2042 2370 2098 2379
rect 2042 2305 2044 2314
rect 2096 2305 2098 2314
rect 2044 2276 2096 2282
rect 1950 1962 2006 1971
rect 1950 1897 2006 1906
rect 2240 1563 2268 11320
rect 2410 11281 2466 11290
rect 2424 10636 2452 11281
rect 2502 11210 2558 11219
rect 2502 11145 2558 11154
rect 2412 10630 2464 10636
rect 2412 10572 2464 10578
rect 2424 10432 2452 10572
rect 2412 10426 2464 10432
rect 2412 10368 2464 10374
rect 2516 9480 2544 11145
rect 2504 9474 2556 9480
rect 2504 9416 2556 9422
rect 2976 7932 3004 15633
rect 3160 13236 3188 18625
rect 3238 18146 3294 18155
rect 3238 18081 3294 18090
rect 3068 13208 3188 13236
rect 3068 8091 3096 13208
rect 3146 13114 3202 13123
rect 3146 13049 3202 13058
rect 3160 12035 3188 13049
rect 3252 12579 3280 18081
rect 3436 17860 3464 19169
rect 3528 18540 3556 21073
rect 3712 18699 3740 23346
rect 3790 19914 3846 19923
rect 3790 19849 3846 19858
rect 3698 18690 3754 18699
rect 3698 18625 3754 18634
rect 3528 18512 3740 18540
rect 3436 17832 3648 17860
rect 3330 17466 3386 17475
rect 3330 17401 3386 17410
rect 3238 12570 3294 12579
rect 3238 12505 3294 12514
rect 3146 12026 3202 12035
rect 3146 11961 3202 11970
rect 3344 9043 3372 17401
rect 3514 16922 3570 16931
rect 3514 16857 3570 16866
rect 3422 14474 3478 14483
rect 3422 14409 3478 14418
rect 3436 13123 3464 14409
rect 3422 13114 3478 13123
rect 3422 13049 3478 13058
rect 3422 11618 3478 11627
rect 3422 11553 3478 11562
rect 3436 10947 3464 11553
rect 3422 10938 3478 10947
rect 3422 10873 3478 10882
rect 3330 9034 3386 9043
rect 3330 8969 3386 8978
rect 3054 8082 3110 8091
rect 3054 8017 3110 8026
rect 2976 7904 3464 7932
rect 3436 3875 3464 7904
rect 3528 5099 3556 16857
rect 3620 12268 3648 17832
rect 3608 12262 3660 12268
rect 3608 12204 3660 12210
rect 3606 12162 3662 12171
rect 3606 12097 3662 12106
rect 3620 10131 3648 12097
rect 3606 10122 3662 10131
rect 3606 10057 3662 10066
rect 3712 9315 3740 18512
rect 3698 9306 3754 9315
rect 3698 9241 3754 9250
rect 3606 8082 3662 8091
rect 3606 8017 3662 8026
rect 3620 7683 3648 8017
rect 3698 7810 3754 7819
rect 3698 7745 3754 7754
rect 3606 7674 3662 7683
rect 3606 7609 3662 7618
rect 3712 7275 3740 7745
rect 3698 7266 3754 7275
rect 3698 7201 3754 7210
rect 3804 7139 3832 19849
rect 3896 18155 3924 23385
rect 11150 23346 11206 23826
rect 18694 23346 18750 23826
rect 25042 23450 25098 23459
rect 25042 23385 25098 23394
rect 5956 21614 6252 21634
rect 6012 21612 6036 21614
rect 6092 21612 6116 21614
rect 6172 21612 6196 21614
rect 6034 21560 6036 21612
rect 6098 21560 6110 21612
rect 6172 21560 6174 21612
rect 6012 21558 6036 21560
rect 6092 21558 6116 21560
rect 6172 21558 6196 21560
rect 5956 21538 6252 21558
rect 11164 21260 11192 23346
rect 15956 21614 16252 21634
rect 16012 21612 16036 21614
rect 16092 21612 16116 21614
rect 16172 21612 16196 21614
rect 16034 21560 16036 21612
rect 16098 21560 16110 21612
rect 16172 21560 16174 21612
rect 16012 21558 16036 21560
rect 16092 21558 16116 21560
rect 16172 21558 16196 21560
rect 15956 21538 16252 21558
rect 11164 21232 11376 21260
rect 10956 21070 11252 21090
rect 11012 21068 11036 21070
rect 11092 21068 11116 21070
rect 11172 21068 11196 21070
rect 11034 21016 11036 21068
rect 11098 21016 11110 21068
rect 11172 21016 11174 21068
rect 11012 21014 11036 21016
rect 11092 21014 11116 21016
rect 11172 21014 11196 21016
rect 10956 20994 11252 21014
rect 5956 20526 6252 20546
rect 6012 20524 6036 20526
rect 6092 20524 6116 20526
rect 6172 20524 6196 20526
rect 6034 20472 6036 20524
rect 6098 20472 6110 20524
rect 6172 20472 6174 20524
rect 6012 20470 6036 20472
rect 6092 20470 6116 20472
rect 6172 20470 6196 20472
rect 3974 20458 4030 20467
rect 5956 20450 6252 20470
rect 3974 20393 4030 20402
rect 3882 18146 3938 18155
rect 3882 18081 3938 18090
rect 3884 12262 3936 12268
rect 3884 12204 3936 12210
rect 3896 7275 3924 12204
rect 3988 8227 4016 20393
rect 10956 19982 11252 20002
rect 11012 19980 11036 19982
rect 11092 19980 11116 19982
rect 11172 19980 11196 19982
rect 11034 19928 11036 19980
rect 11098 19928 11110 19980
rect 11172 19928 11174 19980
rect 11012 19926 11036 19928
rect 11092 19926 11116 19928
rect 11172 19926 11196 19928
rect 10956 19906 11252 19926
rect 5956 19438 6252 19458
rect 6012 19436 6036 19438
rect 6092 19436 6116 19438
rect 6172 19436 6196 19438
rect 6034 19384 6036 19436
rect 6098 19384 6110 19436
rect 6172 19384 6174 19436
rect 6012 19382 6036 19384
rect 6092 19382 6116 19384
rect 6172 19382 6196 19384
rect 5956 19362 6252 19382
rect 11348 19243 11376 21232
rect 15956 20526 16252 20546
rect 16012 20524 16036 20526
rect 16092 20524 16116 20526
rect 16172 20524 16196 20526
rect 16034 20472 16036 20524
rect 16098 20472 16110 20524
rect 16172 20472 16174 20524
rect 16012 20470 16036 20472
rect 16092 20470 16116 20472
rect 16172 20470 16196 20472
rect 15956 20450 16252 20470
rect 15956 19438 16252 19458
rect 16012 19436 16036 19438
rect 16092 19436 16116 19438
rect 16172 19436 16196 19438
rect 16034 19384 16036 19436
rect 16098 19384 16110 19436
rect 16172 19384 16174 19436
rect 16012 19382 16036 19384
rect 16092 19382 16116 19384
rect 16172 19382 16196 19384
rect 15956 19362 16252 19382
rect 8850 19234 8906 19243
rect 8850 19169 8906 19178
rect 11334 19234 11390 19243
rect 11334 19169 11390 19178
rect 8864 18728 8892 19169
rect 10956 18894 11252 18914
rect 11012 18892 11036 18894
rect 11092 18892 11116 18894
rect 11172 18892 11196 18894
rect 11034 18840 11036 18892
rect 11098 18840 11110 18892
rect 11172 18840 11174 18892
rect 11012 18838 11036 18840
rect 11092 18838 11116 18840
rect 11172 18838 11196 18840
rect 10956 18818 11252 18838
rect 18708 18835 18736 23346
rect 24306 22906 24362 22915
rect 24306 22841 24362 22850
rect 20956 21070 21252 21090
rect 21012 21068 21036 21070
rect 21092 21068 21116 21070
rect 21172 21068 21196 21070
rect 21034 21016 21036 21068
rect 21098 21016 21110 21068
rect 21172 21016 21174 21068
rect 21012 21014 21036 21016
rect 21092 21014 21116 21016
rect 21172 21014 21196 21016
rect 20956 20994 21252 21014
rect 19800 20626 19852 20632
rect 19800 20568 19852 20574
rect 20168 20626 20220 20632
rect 20168 20568 20220 20574
rect 16670 18826 16726 18835
rect 16670 18761 16672 18770
rect 16724 18761 16726 18770
rect 18694 18826 18750 18835
rect 18694 18761 18750 18770
rect 16672 18732 16724 18738
rect 8852 18722 8904 18728
rect 7010 18690 7066 18699
rect 7010 18625 7066 18634
rect 8574 18690 8630 18699
rect 8852 18664 8904 18670
rect 12990 18690 13046 18699
rect 8574 18625 8576 18634
rect 5956 18350 6252 18370
rect 6012 18348 6036 18350
rect 6092 18348 6116 18350
rect 6172 18348 6196 18350
rect 6034 18296 6036 18348
rect 6098 18296 6110 18348
rect 6172 18296 6174 18348
rect 6012 18294 6036 18296
rect 6092 18294 6116 18296
rect 6172 18294 6196 18296
rect 5956 18274 6252 18294
rect 5956 17262 6252 17282
rect 6012 17260 6036 17262
rect 6092 17260 6116 17262
rect 6172 17260 6196 17262
rect 6034 17208 6036 17260
rect 6098 17208 6110 17260
rect 6172 17208 6174 17260
rect 6012 17206 6036 17208
rect 6092 17206 6116 17208
rect 6172 17206 6196 17208
rect 5956 17186 6252 17206
rect 4066 16242 4122 16251
rect 4066 16177 4122 16186
rect 3974 8218 4030 8227
rect 3974 8153 4030 8162
rect 3882 7266 3938 7275
rect 3882 7201 3938 7210
rect 3790 7130 3846 7139
rect 4080 7116 4108 16177
rect 5956 16174 6252 16194
rect 6012 16172 6036 16174
rect 6092 16172 6116 16174
rect 6172 16172 6196 16174
rect 6034 16120 6036 16172
rect 6098 16120 6110 16172
rect 6172 16120 6174 16172
rect 6012 16118 6036 16120
rect 6092 16118 6116 16120
rect 6172 16118 6196 16120
rect 5956 16098 6252 16118
rect 7024 16076 7052 18625
rect 8628 18625 8630 18634
rect 8576 18596 8628 18602
rect 8588 18184 8616 18596
rect 8864 18252 8892 18664
rect 15290 18690 15346 18699
rect 12990 18625 13046 18634
rect 15200 18654 15252 18660
rect 9956 18450 10008 18456
rect 9956 18392 10008 18398
rect 8852 18246 8904 18252
rect 8852 18188 8904 18194
rect 8576 18178 8628 18184
rect 8576 18120 8628 18126
rect 7012 16070 7064 16076
rect 7012 16012 7064 16018
rect 9968 15843 9996 18392
rect 10956 17806 11252 17826
rect 11012 17804 11036 17806
rect 11092 17804 11116 17806
rect 11172 17804 11196 17806
rect 11034 17752 11036 17804
rect 11098 17752 11110 17804
rect 11172 17752 11174 17804
rect 11012 17750 11036 17752
rect 11092 17750 11116 17752
rect 11172 17750 11196 17752
rect 10956 17730 11252 17750
rect 10956 16718 11252 16738
rect 11012 16716 11036 16718
rect 11092 16716 11116 16718
rect 11172 16716 11196 16718
rect 11034 16664 11036 16716
rect 11098 16664 11110 16716
rect 11172 16664 11174 16716
rect 11012 16662 11036 16664
rect 11092 16662 11116 16664
rect 11172 16662 11196 16664
rect 10956 16642 11252 16662
rect 13004 16484 13032 18625
rect 15290 18625 15346 18634
rect 15200 18596 15252 18602
rect 15212 17980 15240 18596
rect 15304 18592 15332 18625
rect 15292 18586 15344 18592
rect 15292 18528 15344 18534
rect 15304 18252 15332 18528
rect 15956 18350 16252 18370
rect 16012 18348 16036 18350
rect 16092 18348 16116 18350
rect 16172 18348 16196 18350
rect 16034 18296 16036 18348
rect 16098 18296 16110 18348
rect 16172 18296 16174 18348
rect 16012 18294 16036 18296
rect 16092 18294 16116 18296
rect 16172 18294 16196 18296
rect 15956 18274 16252 18294
rect 15292 18246 15344 18252
rect 15292 18188 15344 18194
rect 15200 17974 15252 17980
rect 15200 17916 15252 17922
rect 13542 16786 13598 16795
rect 13542 16721 13598 16730
rect 12992 16478 13044 16484
rect 12992 16420 13044 16426
rect 13004 16076 13032 16420
rect 12992 16070 13044 16076
rect 12992 16012 13044 16018
rect 7194 15834 7250 15843
rect 7194 15769 7196 15778
rect 7248 15769 7250 15778
rect 9954 15834 10010 15843
rect 9954 15769 10010 15778
rect 7196 15740 7248 15746
rect 7208 15532 7236 15740
rect 8576 15730 8628 15736
rect 8576 15672 8628 15678
rect 7196 15526 7248 15532
rect 7196 15468 7248 15474
rect 5956 15086 6252 15106
rect 6012 15084 6036 15086
rect 6092 15084 6116 15086
rect 6172 15084 6196 15086
rect 6034 15032 6036 15084
rect 6098 15032 6110 15084
rect 6172 15032 6174 15084
rect 6012 15030 6036 15032
rect 6092 15030 6116 15032
rect 6172 15030 6196 15032
rect 5956 15010 6252 15030
rect 5956 13998 6252 14018
rect 6012 13996 6036 13998
rect 6092 13996 6116 13998
rect 6172 13996 6196 13998
rect 6034 13944 6036 13996
rect 6098 13944 6110 13996
rect 6172 13944 6174 13996
rect 6012 13942 6036 13944
rect 6092 13942 6116 13944
rect 6172 13942 6196 13944
rect 5956 13922 6252 13942
rect 5956 12910 6252 12930
rect 6012 12908 6036 12910
rect 6092 12908 6116 12910
rect 6172 12908 6196 12910
rect 6034 12856 6036 12908
rect 6098 12856 6110 12908
rect 6172 12856 6174 12908
rect 6012 12854 6036 12856
rect 6092 12854 6116 12856
rect 6172 12854 6196 12856
rect 5956 12834 6252 12854
rect 5956 11822 6252 11842
rect 6012 11820 6036 11822
rect 6092 11820 6116 11822
rect 6172 11820 6196 11822
rect 6034 11768 6036 11820
rect 6098 11768 6110 11820
rect 6172 11768 6174 11820
rect 6012 11766 6036 11768
rect 6092 11766 6116 11768
rect 6172 11766 6196 11768
rect 5956 11746 6252 11766
rect 6642 11618 6698 11627
rect 6642 11553 6698 11562
rect 6656 11355 6684 11553
rect 6642 11346 6698 11355
rect 6642 11281 6698 11290
rect 7102 11210 7158 11219
rect 7102 11145 7158 11154
rect 5956 10734 6252 10754
rect 6012 10732 6036 10734
rect 6092 10732 6116 10734
rect 6172 10732 6196 10734
rect 6034 10680 6036 10732
rect 6098 10680 6110 10732
rect 6172 10680 6174 10732
rect 6012 10678 6036 10680
rect 6092 10678 6116 10680
rect 6172 10678 6196 10680
rect 5956 10658 6252 10678
rect 7116 10568 7144 11145
rect 7208 11112 7236 15468
rect 8588 12064 8616 15672
rect 10956 15630 11252 15650
rect 11012 15628 11036 15630
rect 11092 15628 11116 15630
rect 11172 15628 11196 15630
rect 11034 15576 11036 15628
rect 11098 15576 11110 15628
rect 11172 15576 11174 15628
rect 11012 15574 11036 15576
rect 11092 15574 11116 15576
rect 11172 15574 11196 15576
rect 10956 15554 11252 15574
rect 10956 14542 11252 14562
rect 11012 14540 11036 14542
rect 11092 14540 11116 14542
rect 11172 14540 11196 14542
rect 11034 14488 11036 14540
rect 11098 14488 11110 14540
rect 11172 14488 11174 14540
rect 11012 14486 11036 14488
rect 11092 14486 11116 14488
rect 11172 14486 11196 14488
rect 10956 14466 11252 14486
rect 10956 13454 11252 13474
rect 11012 13452 11036 13454
rect 11092 13452 11116 13454
rect 11172 13452 11196 13454
rect 11034 13400 11036 13452
rect 11098 13400 11110 13452
rect 11172 13400 11174 13452
rect 11012 13398 11036 13400
rect 11092 13398 11116 13400
rect 11172 13398 11196 13400
rect 10956 13378 11252 13398
rect 13556 13356 13584 16721
rect 15212 16620 15240 17916
rect 15956 17262 16252 17282
rect 16012 17260 16036 17262
rect 16092 17260 16116 17262
rect 16172 17260 16196 17262
rect 16034 17208 16036 17260
rect 16098 17208 16110 17260
rect 16172 17208 16174 17260
rect 16012 17206 16036 17208
rect 16092 17206 16116 17208
rect 16172 17206 16196 17208
rect 15956 17186 16252 17206
rect 18708 17028 18736 18761
rect 19340 17906 19392 17912
rect 19260 17854 19340 17860
rect 19260 17848 19392 17854
rect 19260 17832 19380 17848
rect 19260 17164 19288 17832
rect 19248 17158 19300 17164
rect 19248 17100 19300 17106
rect 18696 17022 18748 17028
rect 18696 16964 18748 16970
rect 17500 16818 17552 16824
rect 17498 16786 17500 16795
rect 18328 16818 18380 16824
rect 17552 16786 17554 16795
rect 18328 16760 18380 16766
rect 17498 16721 17554 16730
rect 18340 16620 18368 16760
rect 14188 16614 14240 16620
rect 14188 16556 14240 16562
rect 15200 16614 15252 16620
rect 15200 16556 15252 16562
rect 18328 16614 18380 16620
rect 18328 16556 18380 16562
rect 13728 16478 13780 16484
rect 13728 16420 13780 16426
rect 13740 15736 13768 16420
rect 13728 15730 13780 15736
rect 13728 15672 13780 15678
rect 13544 13350 13596 13356
rect 13544 13292 13596 13298
rect 11886 13114 11942 13123
rect 11886 13049 11942 13058
rect 10956 12366 11252 12386
rect 11012 12364 11036 12366
rect 11092 12364 11116 12366
rect 11172 12364 11196 12366
rect 11034 12312 11036 12364
rect 11098 12312 11110 12364
rect 11172 12312 11174 12364
rect 11012 12310 11036 12312
rect 11092 12310 11116 12312
rect 11172 12310 11196 12312
rect 10956 12290 11252 12310
rect 8668 12126 8720 12132
rect 8668 12068 8720 12074
rect 8576 12058 8628 12064
rect 7378 12026 7434 12035
rect 7378 11961 7434 11970
rect 7930 12026 7986 12035
rect 8576 12000 8628 12006
rect 7930 11961 7932 11970
rect 7196 11106 7248 11112
rect 7196 11048 7248 11054
rect 7392 10976 7420 11961
rect 7984 11961 7986 11970
rect 8300 11990 8352 11996
rect 7932 11932 7984 11938
rect 8300 11932 8352 11938
rect 8312 11384 8340 11932
rect 8390 11890 8446 11899
rect 8390 11825 8446 11834
rect 8300 11378 8352 11384
rect 8300 11320 8352 11326
rect 8312 11196 8340 11320
rect 8220 11168 8340 11196
rect 8116 11038 8168 11044
rect 8116 10980 8168 10986
rect 7380 10970 7432 10976
rect 8128 10947 8156 10980
rect 7380 10912 7432 10918
rect 8114 10938 8170 10947
rect 7104 10562 7156 10568
rect 7104 10504 7156 10510
rect 7392 10296 7420 10912
rect 8114 10873 8170 10882
rect 8128 10568 8156 10873
rect 8220 10636 8248 11168
rect 8404 10976 8432 11825
rect 8588 11724 8616 12000
rect 8576 11718 8628 11724
rect 8576 11660 8628 11666
rect 8680 11384 8708 12068
rect 11900 11724 11928 13049
rect 13084 13010 13136 13016
rect 13084 12952 13136 12958
rect 12900 12602 12952 12608
rect 12898 12570 12900 12579
rect 12952 12570 12954 12579
rect 12440 12534 12492 12540
rect 13096 12540 13124 12952
rect 13740 12676 13768 15672
rect 14200 14891 14228 16556
rect 15956 16174 16252 16194
rect 16012 16172 16036 16174
rect 16092 16172 16116 16174
rect 16172 16172 16196 16174
rect 16034 16120 16036 16172
rect 16098 16120 16110 16172
rect 16172 16120 16174 16172
rect 16012 16118 16036 16120
rect 16092 16118 16116 16120
rect 16172 16118 16196 16120
rect 15956 16098 16252 16118
rect 15956 15086 16252 15106
rect 16012 15084 16036 15086
rect 16092 15084 16116 15086
rect 16172 15084 16196 15086
rect 16034 15032 16036 15084
rect 16098 15032 16110 15084
rect 16172 15032 16174 15084
rect 16012 15030 16036 15032
rect 16092 15030 16116 15032
rect 16172 15030 16196 15032
rect 15956 15010 16252 15030
rect 18340 14988 18368 16556
rect 18604 15186 18656 15192
rect 18604 15128 18656 15134
rect 18328 14982 18380 14988
rect 18328 14924 18380 14930
rect 14186 14882 14242 14891
rect 14186 14817 14242 14826
rect 18326 14882 18382 14891
rect 18326 14817 18328 14826
rect 13912 13214 13964 13220
rect 13912 13156 13964 13162
rect 13820 13146 13872 13152
rect 13820 13088 13872 13094
rect 13728 12670 13780 12676
rect 13728 12612 13780 12618
rect 12898 12505 12954 12514
rect 13084 12534 13136 12540
rect 12440 12476 12492 12482
rect 13084 12476 13136 12482
rect 12452 12420 12480 12476
rect 12360 12392 12480 12420
rect 12072 11922 12124 11928
rect 12070 11890 12072 11899
rect 12124 11890 12126 11899
rect 12070 11825 12126 11834
rect 11888 11718 11940 11724
rect 11888 11660 11940 11666
rect 11518 11618 11574 11627
rect 11518 11553 11574 11562
rect 11532 11452 11560 11553
rect 11900 11520 11928 11660
rect 12084 11588 12112 11825
rect 12360 11724 12388 12392
rect 13740 12200 13768 12612
rect 13728 12194 13780 12200
rect 13726 12162 13728 12171
rect 13780 12162 13782 12171
rect 13726 12097 13782 12106
rect 13740 12071 13768 12097
rect 13832 12035 13860 13088
rect 13924 12744 13952 13156
rect 14200 13152 14228 14817
rect 18380 14817 18382 14826
rect 18328 14788 18380 14794
rect 18616 14716 18644 15128
rect 18604 14710 18656 14716
rect 18604 14652 18656 14658
rect 19248 14710 19300 14716
rect 19248 14652 19300 14658
rect 18972 14642 19024 14648
rect 18972 14584 19024 14590
rect 19260 14596 19288 14652
rect 18984 14444 19012 14584
rect 19260 14568 19380 14596
rect 18972 14438 19024 14444
rect 18972 14380 19024 14386
rect 15956 13998 16252 14018
rect 16012 13996 16036 13998
rect 16092 13996 16116 13998
rect 16172 13996 16196 13998
rect 16034 13944 16036 13996
rect 16098 13944 16110 13996
rect 16172 13944 16174 13996
rect 16012 13942 16036 13944
rect 16092 13942 16116 13944
rect 16172 13942 16196 13944
rect 15956 13922 16252 13942
rect 19064 13554 19116 13560
rect 19064 13496 19116 13502
rect 19076 13356 19104 13496
rect 19064 13350 19116 13356
rect 19064 13292 19116 13298
rect 14188 13146 14240 13152
rect 14188 13088 14240 13094
rect 14200 12812 14228 13088
rect 19352 13084 19380 14568
rect 19812 14308 19840 20568
rect 19890 18282 19946 18291
rect 19890 18217 19946 18226
rect 19616 14302 19668 14308
rect 19616 14244 19668 14250
rect 19800 14302 19852 14308
rect 19800 14244 19852 14250
rect 19628 13696 19656 14244
rect 19904 14240 19932 18217
rect 19892 14234 19944 14240
rect 19892 14176 19944 14182
rect 19904 13696 19932 14176
rect 19616 13690 19668 13696
rect 19616 13632 19668 13638
rect 19892 13690 19944 13696
rect 19892 13632 19944 13638
rect 19628 13123 19656 13632
rect 19904 13259 19932 13632
rect 20076 13350 20128 13356
rect 20076 13292 20128 13298
rect 19890 13250 19946 13259
rect 19708 13214 19760 13220
rect 19890 13185 19946 13194
rect 19708 13156 19760 13162
rect 19614 13114 19670 13123
rect 19340 13078 19392 13084
rect 19614 13049 19670 13058
rect 19340 13020 19392 13026
rect 15956 12910 16252 12930
rect 16012 12908 16036 12910
rect 16092 12908 16116 12910
rect 16172 12908 16196 12910
rect 16034 12856 16036 12908
rect 16098 12856 16110 12908
rect 16172 12856 16174 12908
rect 16012 12854 16036 12856
rect 16092 12854 16116 12856
rect 16172 12854 16196 12856
rect 15956 12834 16252 12854
rect 14188 12806 14240 12812
rect 14188 12748 14240 12754
rect 13912 12738 13964 12744
rect 13912 12680 13964 12686
rect 13924 12268 13952 12680
rect 14646 12570 14702 12579
rect 14646 12505 14702 12514
rect 13912 12262 13964 12268
rect 13912 12204 13964 12210
rect 13818 12026 13874 12035
rect 13740 11996 13818 12012
rect 13728 11990 13818 11996
rect 13780 11984 13818 11990
rect 13818 11961 13874 11970
rect 13728 11932 13780 11938
rect 12348 11718 12400 11724
rect 12348 11660 12400 11666
rect 12072 11582 12124 11588
rect 12072 11524 12124 11530
rect 11888 11514 11940 11520
rect 11888 11456 11940 11462
rect 12532 11514 12584 11520
rect 12532 11456 12584 11462
rect 13726 11482 13782 11491
rect 11520 11446 11572 11452
rect 11520 11388 11572 11394
rect 8668 11378 8720 11384
rect 8668 11320 8720 11326
rect 8680 11180 8708 11320
rect 10956 11278 11252 11298
rect 11012 11276 11036 11278
rect 11092 11276 11116 11278
rect 11172 11276 11196 11278
rect 11034 11224 11036 11276
rect 11098 11224 11110 11276
rect 11172 11224 11174 11276
rect 11012 11222 11036 11224
rect 11092 11222 11116 11224
rect 11172 11222 11196 11224
rect 10956 11202 11252 11222
rect 11532 11180 11560 11388
rect 12544 11384 12572 11456
rect 13726 11417 13728 11426
rect 13780 11417 13782 11426
rect 13728 11388 13780 11394
rect 12532 11378 12584 11384
rect 12532 11320 12584 11326
rect 12438 11210 12494 11219
rect 8668 11174 8720 11180
rect 8668 11116 8720 11122
rect 11520 11174 11572 11180
rect 12438 11145 12494 11154
rect 11520 11116 11572 11122
rect 8392 10970 8444 10976
rect 12452 10947 12480 11145
rect 8392 10912 8444 10918
rect 12438 10938 12494 10947
rect 8404 10636 8432 10912
rect 12438 10873 12494 10882
rect 8208 10630 8260 10636
rect 8208 10572 8260 10578
rect 8392 10630 8444 10636
rect 8392 10572 8444 10578
rect 8116 10562 8168 10568
rect 8116 10504 8168 10510
rect 8298 10394 8354 10403
rect 8404 10380 8432 10572
rect 8404 10352 8524 10380
rect 8298 10329 8300 10338
rect 8352 10329 8354 10338
rect 8300 10300 8352 10306
rect 7380 10290 7432 10296
rect 7380 10232 7432 10238
rect 7840 10290 7892 10296
rect 7840 10232 7892 10238
rect 5956 9646 6252 9666
rect 6012 9644 6036 9646
rect 6092 9644 6116 9646
rect 6172 9644 6196 9646
rect 6034 9592 6036 9644
rect 6098 9592 6110 9644
rect 6172 9592 6174 9644
rect 6012 9590 6036 9592
rect 6092 9590 6116 9592
rect 6172 9590 6196 9592
rect 5956 9570 6252 9590
rect 4802 9034 4858 9043
rect 4802 8969 4858 8978
rect 3790 7065 3846 7074
rect 3896 7088 4108 7116
rect 3514 5090 3570 5099
rect 3514 5025 3570 5034
rect 3896 4555 3924 7088
rect 4816 5604 4844 8969
rect 5956 8558 6252 8578
rect 6012 8556 6036 8558
rect 6092 8556 6116 8558
rect 6172 8556 6196 8558
rect 6034 8504 6036 8556
rect 6098 8504 6110 8556
rect 6172 8504 6174 8556
rect 6012 8502 6036 8504
rect 6092 8502 6116 8504
rect 6172 8502 6196 8504
rect 5956 8482 6252 8502
rect 5956 7470 6252 7490
rect 6012 7468 6036 7470
rect 6092 7468 6116 7470
rect 6172 7468 6196 7470
rect 6034 7416 6036 7468
rect 6098 7416 6110 7468
rect 6172 7416 6174 7468
rect 6012 7414 6036 7416
rect 6092 7414 6116 7416
rect 6172 7414 6196 7416
rect 5956 7394 6252 7414
rect 5956 6382 6252 6402
rect 6012 6380 6036 6382
rect 6092 6380 6116 6382
rect 6172 6380 6196 6382
rect 6034 6328 6036 6380
rect 6098 6328 6110 6380
rect 6172 6328 6174 6380
rect 6012 6326 6036 6328
rect 6092 6326 6116 6328
rect 6172 6326 6196 6328
rect 5956 6306 6252 6326
rect 4804 5598 4856 5604
rect 4804 5540 4856 5546
rect 4816 5196 4844 5540
rect 4986 5498 5042 5507
rect 4986 5433 4988 5442
rect 5040 5433 5042 5442
rect 4988 5404 5040 5410
rect 5956 5294 6252 5314
rect 6012 5292 6036 5294
rect 6092 5292 6116 5294
rect 6172 5292 6196 5294
rect 6034 5240 6036 5292
rect 6098 5240 6110 5292
rect 6172 5240 6174 5292
rect 6012 5238 6036 5240
rect 6092 5238 6116 5240
rect 6172 5238 6196 5240
rect 5956 5218 6252 5238
rect 4804 5190 4856 5196
rect 4804 5132 4856 5138
rect 3882 4546 3938 4555
rect 3882 4481 3938 4490
rect 5956 4206 6252 4226
rect 6012 4204 6036 4206
rect 6092 4204 6116 4206
rect 6172 4204 6196 4206
rect 6034 4152 6036 4204
rect 6098 4152 6110 4204
rect 6172 4152 6174 4204
rect 6012 4150 6036 4152
rect 6092 4150 6116 4152
rect 6172 4150 6196 4152
rect 5956 4130 6252 4150
rect 3422 3866 3478 3875
rect 3422 3801 3478 3810
rect 5956 3118 6252 3138
rect 6012 3116 6036 3118
rect 6092 3116 6116 3118
rect 6172 3116 6196 3118
rect 6034 3064 6036 3116
rect 6098 3064 6110 3116
rect 6172 3064 6174 3116
rect 6012 3062 6036 3064
rect 6092 3062 6116 3064
rect 6172 3062 6196 3064
rect 5956 3042 6252 3062
rect 7392 2923 7420 10232
rect 7852 10131 7880 10232
rect 7838 10122 7894 10131
rect 8312 10092 8340 10300
rect 8392 10290 8444 10296
rect 8392 10232 8444 10238
rect 7838 10057 7894 10066
rect 8300 10086 8352 10092
rect 8300 10028 8352 10034
rect 8312 9995 8340 10028
rect 8298 9986 8354 9995
rect 8298 9921 8354 9930
rect 7378 2914 7434 2923
rect 7378 2849 7434 2858
rect 2688 2674 2740 2680
rect 2688 2616 2740 2622
rect 2226 1554 2282 1563
rect 2226 1489 2282 1498
rect 1674 1282 1730 1291
rect 1674 1217 1730 1226
rect 1582 738 1638 747
rect 1582 673 1638 682
rect 2700 203 2728 2616
rect 5956 2030 6252 2050
rect 6012 2028 6036 2030
rect 6092 2028 6116 2030
rect 6172 2028 6196 2030
rect 6034 1976 6036 2028
rect 6098 1976 6110 2028
rect 6172 1976 6174 2028
rect 6012 1974 6036 1976
rect 6092 1974 6116 1976
rect 6172 1974 6196 1976
rect 5956 1954 6252 1974
rect 8404 1835 8432 10232
rect 8496 10092 8524 10352
rect 10956 10190 11252 10210
rect 11012 10188 11036 10190
rect 11092 10188 11116 10190
rect 11172 10188 11196 10190
rect 11034 10136 11036 10188
rect 11098 10136 11110 10188
rect 11172 10136 11174 10188
rect 11012 10134 11036 10136
rect 11092 10134 11116 10136
rect 11172 10134 11196 10136
rect 10956 10114 11252 10134
rect 8484 10086 8536 10092
rect 8484 10028 8536 10034
rect 10956 9102 11252 9122
rect 11012 9100 11036 9102
rect 11092 9100 11116 9102
rect 11172 9100 11196 9102
rect 11034 9048 11036 9100
rect 11098 9048 11110 9100
rect 11172 9048 11174 9100
rect 11012 9046 11036 9048
rect 11092 9046 11116 9048
rect 11172 9046 11196 9048
rect 10956 9026 11252 9046
rect 10784 8114 10836 8120
rect 10782 8082 10784 8091
rect 11336 8114 11388 8120
rect 10836 8082 10838 8091
rect 11334 8082 11336 8091
rect 11388 8082 11390 8091
rect 10782 8017 10838 8026
rect 10956 8014 11252 8034
rect 11334 8017 11390 8026
rect 11012 8012 11036 8014
rect 11092 8012 11116 8014
rect 11172 8012 11196 8014
rect 11034 7960 11036 8012
rect 11098 7960 11110 8012
rect 11172 7960 11174 8012
rect 11012 7958 11036 7960
rect 11092 7958 11116 7960
rect 11172 7958 11196 7960
rect 10956 7938 11252 7958
rect 10874 7674 10930 7683
rect 10874 7609 10930 7618
rect 10888 6692 10916 7609
rect 10956 6926 11252 6946
rect 11012 6924 11036 6926
rect 11092 6924 11116 6926
rect 11172 6924 11196 6926
rect 11034 6872 11036 6924
rect 11098 6872 11110 6924
rect 11172 6872 11174 6924
rect 11012 6870 11036 6872
rect 11092 6870 11116 6872
rect 11172 6870 11196 6872
rect 10956 6850 11252 6870
rect 10876 6686 10928 6692
rect 10876 6628 10928 6634
rect 10888 6284 10916 6628
rect 11060 6482 11112 6488
rect 11060 6424 11112 6430
rect 10876 6278 10928 6284
rect 10876 6220 10928 6226
rect 11072 6187 11100 6424
rect 11058 6178 11114 6187
rect 11058 6113 11114 6122
rect 10956 5838 11252 5858
rect 11012 5836 11036 5838
rect 11092 5836 11116 5838
rect 11172 5836 11196 5838
rect 11034 5784 11036 5836
rect 11098 5784 11110 5836
rect 11172 5784 11174 5836
rect 11012 5782 11036 5784
rect 11092 5782 11116 5784
rect 11172 5782 11196 5784
rect 10956 5762 11252 5782
rect 10956 4750 11252 4770
rect 11012 4748 11036 4750
rect 11092 4748 11116 4750
rect 11172 4748 11196 4750
rect 11034 4696 11036 4748
rect 11098 4696 11110 4748
rect 11172 4696 11174 4748
rect 11012 4694 11036 4696
rect 11092 4694 11116 4696
rect 11172 4694 11196 4696
rect 10956 4674 11252 4694
rect 10956 3662 11252 3682
rect 11012 3660 11036 3662
rect 11092 3660 11116 3662
rect 11172 3660 11196 3662
rect 11034 3608 11036 3660
rect 11098 3608 11110 3660
rect 11172 3608 11174 3660
rect 11012 3606 11036 3608
rect 11092 3606 11116 3608
rect 11172 3606 11196 3608
rect 10956 3586 11252 3606
rect 10956 2574 11252 2594
rect 11012 2572 11036 2574
rect 11092 2572 11116 2574
rect 11172 2572 11196 2574
rect 11034 2520 11036 2572
rect 11098 2520 11110 2572
rect 11172 2520 11174 2572
rect 11012 2518 11036 2520
rect 11092 2518 11116 2520
rect 11172 2518 11196 2520
rect 10956 2498 11252 2518
rect 12544 2243 12572 11320
rect 14660 6692 14688 12505
rect 19720 12472 19748 13156
rect 20088 12812 20116 13292
rect 20180 13220 20208 20568
rect 20956 19982 21252 20002
rect 21012 19980 21036 19982
rect 21092 19980 21116 19982
rect 21172 19980 21196 19982
rect 21034 19928 21036 19980
rect 21098 19928 21110 19980
rect 21172 19928 21174 19980
rect 21012 19926 21036 19928
rect 21092 19926 21116 19928
rect 21172 19926 21196 19928
rect 20956 19906 21252 19926
rect 20626 19642 20682 19651
rect 20626 19577 20682 19586
rect 20640 18796 20668 19577
rect 23940 19130 23992 19136
rect 23938 19098 23940 19107
rect 23992 19098 23994 19107
rect 23938 19033 23994 19042
rect 20956 18894 21252 18914
rect 21012 18892 21036 18894
rect 21092 18892 21116 18894
rect 21172 18892 21196 18894
rect 21034 18840 21036 18892
rect 21098 18840 21110 18892
rect 21172 18840 21174 18892
rect 21012 18838 21036 18840
rect 21092 18838 21116 18840
rect 21172 18838 21196 18840
rect 20956 18818 21252 18838
rect 20628 18790 20680 18796
rect 20628 18732 20680 18738
rect 20444 18654 20496 18660
rect 20444 18596 20496 18602
rect 23756 18654 23808 18660
rect 23756 18596 23808 18602
rect 20456 17912 20484 18596
rect 23768 18184 23796 18596
rect 24124 18450 24176 18456
rect 24124 18392 24176 18398
rect 23756 18178 23808 18184
rect 23754 18146 23756 18155
rect 23808 18146 23810 18155
rect 23754 18081 23810 18090
rect 23940 18042 23992 18048
rect 23938 18010 23940 18019
rect 23992 18010 23994 18019
rect 23938 17945 23994 17954
rect 20444 17906 20496 17912
rect 20444 17848 20496 17854
rect 20956 17806 21252 17826
rect 21012 17804 21036 17806
rect 21092 17804 21116 17806
rect 21172 17804 21196 17806
rect 21034 17752 21036 17804
rect 21098 17752 21110 17804
rect 21172 17752 21174 17804
rect 21012 17750 21036 17752
rect 21092 17750 21116 17752
rect 21172 17750 21196 17752
rect 20956 17730 21252 17750
rect 23480 17362 23532 17368
rect 23480 17304 23532 17310
rect 20956 16718 21252 16738
rect 21012 16716 21036 16718
rect 21092 16716 21116 16718
rect 21172 16716 21196 16718
rect 21034 16664 21036 16716
rect 21098 16664 21110 16716
rect 21172 16664 21174 16716
rect 21012 16662 21036 16664
rect 21092 16662 21116 16664
rect 21172 16662 21196 16664
rect 20956 16642 21252 16662
rect 20956 15630 21252 15650
rect 21012 15628 21036 15630
rect 21092 15628 21116 15630
rect 21172 15628 21196 15630
rect 21034 15576 21036 15628
rect 21098 15576 21110 15628
rect 21172 15576 21174 15628
rect 21012 15574 21036 15576
rect 21092 15574 21116 15576
rect 21172 15574 21196 15576
rect 20956 15554 21252 15574
rect 20956 14542 21252 14562
rect 21012 14540 21036 14542
rect 21092 14540 21116 14542
rect 21172 14540 21196 14542
rect 21034 14488 21036 14540
rect 21098 14488 21110 14540
rect 21172 14488 21174 14540
rect 21012 14486 21036 14488
rect 21092 14486 21116 14488
rect 21172 14486 21196 14488
rect 20956 14466 21252 14486
rect 20444 14234 20496 14240
rect 20444 14176 20496 14182
rect 20456 13560 20484 14176
rect 23110 13658 23166 13667
rect 23110 13593 23166 13602
rect 20444 13554 20496 13560
rect 20444 13496 20496 13502
rect 20168 13214 20220 13220
rect 20168 13156 20220 13162
rect 20456 13152 20484 13496
rect 20956 13454 21252 13474
rect 21012 13452 21036 13454
rect 21092 13452 21116 13454
rect 21172 13452 21196 13454
rect 21034 13400 21036 13452
rect 21098 13400 21110 13452
rect 21172 13400 21174 13452
rect 21012 13398 21036 13400
rect 21092 13398 21116 13400
rect 21172 13398 21196 13400
rect 20956 13378 21252 13398
rect 20444 13146 20496 13152
rect 20444 13088 20496 13094
rect 20076 12806 20128 12812
rect 20076 12748 20128 12754
rect 20456 12472 20484 13088
rect 19708 12466 19760 12472
rect 19708 12408 19760 12414
rect 20444 12466 20496 12472
rect 20444 12408 20496 12414
rect 17222 12026 17278 12035
rect 17222 11961 17278 11970
rect 15956 11822 16252 11842
rect 16012 11820 16036 11822
rect 16092 11820 16116 11822
rect 16172 11820 16196 11822
rect 16034 11768 16036 11820
rect 16098 11768 16110 11820
rect 16172 11768 16174 11820
rect 16012 11766 16036 11768
rect 16092 11766 16116 11768
rect 16172 11766 16196 11768
rect 15956 11746 16252 11766
rect 17236 11355 17264 11961
rect 17498 11618 17554 11627
rect 17498 11553 17554 11562
rect 17222 11346 17278 11355
rect 17222 11281 17278 11290
rect 17512 11083 17540 11553
rect 17498 11074 17554 11083
rect 17498 11009 17554 11018
rect 15956 10734 16252 10754
rect 16012 10732 16036 10734
rect 16092 10732 16116 10734
rect 16172 10732 16196 10734
rect 16034 10680 16036 10732
rect 16098 10680 16110 10732
rect 16172 10680 16174 10732
rect 16012 10678 16036 10680
rect 16092 10678 16116 10680
rect 16172 10678 16196 10680
rect 15956 10658 16252 10678
rect 19720 9859 19748 12408
rect 20456 12171 20484 12408
rect 20956 12366 21252 12386
rect 21012 12364 21036 12366
rect 21092 12364 21116 12366
rect 21172 12364 21196 12366
rect 21034 12312 21036 12364
rect 21098 12312 21110 12364
rect 21172 12312 21174 12364
rect 21012 12310 21036 12312
rect 21092 12310 21116 12312
rect 21172 12310 21196 12312
rect 20956 12290 21252 12310
rect 20442 12162 20498 12171
rect 20442 12097 20498 12106
rect 20956 11278 21252 11298
rect 21012 11276 21036 11278
rect 21092 11276 21116 11278
rect 21172 11276 21196 11278
rect 21034 11224 21036 11276
rect 21098 11224 21110 11276
rect 21172 11224 21174 11276
rect 21012 11222 21036 11224
rect 21092 11222 21116 11224
rect 21172 11222 21196 11224
rect 20956 11202 21252 11222
rect 20956 10190 21252 10210
rect 21012 10188 21036 10190
rect 21092 10188 21116 10190
rect 21172 10188 21196 10190
rect 21034 10136 21036 10188
rect 21098 10136 21110 10188
rect 21172 10136 21174 10188
rect 21012 10134 21036 10136
rect 21092 10134 21116 10136
rect 21172 10134 21196 10136
rect 20956 10114 21252 10134
rect 19706 9850 19762 9859
rect 19706 9785 19762 9794
rect 15956 9646 16252 9666
rect 16012 9644 16036 9646
rect 16092 9644 16116 9646
rect 16172 9644 16196 9646
rect 16034 9592 16036 9644
rect 16098 9592 16110 9644
rect 16172 9592 16174 9644
rect 16012 9590 16036 9592
rect 16092 9590 16116 9592
rect 16172 9590 16196 9592
rect 15956 9570 16252 9590
rect 20956 9102 21252 9122
rect 21012 9100 21036 9102
rect 21092 9100 21116 9102
rect 21172 9100 21196 9102
rect 21034 9048 21036 9100
rect 21098 9048 21110 9100
rect 21172 9048 21174 9100
rect 21012 9046 21036 9048
rect 21092 9046 21116 9048
rect 21172 9046 21196 9048
rect 20956 9026 21252 9046
rect 15956 8558 16252 8578
rect 16012 8556 16036 8558
rect 16092 8556 16116 8558
rect 16172 8556 16196 8558
rect 16034 8504 16036 8556
rect 16098 8504 16110 8556
rect 16172 8504 16174 8556
rect 16012 8502 16036 8504
rect 16092 8502 16116 8504
rect 16172 8502 16196 8504
rect 15956 8482 16252 8502
rect 20956 8014 21252 8034
rect 21012 8012 21036 8014
rect 21092 8012 21116 8014
rect 21172 8012 21196 8014
rect 21034 7960 21036 8012
rect 21098 7960 21110 8012
rect 21172 7960 21174 8012
rect 21012 7958 21036 7960
rect 21092 7958 21116 7960
rect 21172 7958 21196 7960
rect 20956 7938 21252 7958
rect 22650 7538 22706 7547
rect 15956 7470 16252 7490
rect 22650 7473 22706 7482
rect 16012 7468 16036 7470
rect 16092 7468 16116 7470
rect 16172 7468 16196 7470
rect 16034 7416 16036 7468
rect 16098 7416 16110 7468
rect 16172 7416 16174 7468
rect 16012 7414 16036 7416
rect 16092 7414 16116 7416
rect 16172 7414 16196 7416
rect 15956 7394 16252 7414
rect 22664 7372 22692 7473
rect 23124 7372 23152 13593
rect 23492 13236 23520 17304
rect 23570 16922 23626 16931
rect 23570 16857 23626 16866
rect 23400 13208 23520 13236
rect 23400 11899 23428 13208
rect 23478 13114 23534 13123
rect 23478 13049 23534 13058
rect 23386 11890 23442 11899
rect 23386 11825 23442 11834
rect 23492 11520 23520 13049
rect 23480 11514 23532 11520
rect 23480 11456 23532 11462
rect 23480 8386 23532 8392
rect 23480 8328 23532 8334
rect 23492 7819 23520 8328
rect 23478 7810 23534 7819
rect 23478 7745 23534 7754
rect 22652 7366 22704 7372
rect 22652 7308 22704 7314
rect 23112 7366 23164 7372
rect 23112 7308 23164 7314
rect 18880 7298 18932 7304
rect 18694 7266 18750 7275
rect 18694 7201 18750 7210
rect 18878 7266 18880 7275
rect 18932 7266 18934 7275
rect 18878 7201 18934 7210
rect 18708 7168 18736 7201
rect 23124 7168 23152 7308
rect 18696 7162 18748 7168
rect 18696 7104 18748 7110
rect 23112 7162 23164 7168
rect 23112 7104 23164 7110
rect 20956 6926 21252 6946
rect 21012 6924 21036 6926
rect 21092 6924 21116 6926
rect 21172 6924 21196 6926
rect 21034 6872 21036 6924
rect 21098 6872 21110 6924
rect 21172 6872 21174 6924
rect 21012 6870 21036 6872
rect 21092 6870 21116 6872
rect 21172 6870 21196 6872
rect 20956 6850 21252 6870
rect 14648 6686 14700 6692
rect 14648 6628 14700 6634
rect 14660 6284 14688 6628
rect 14832 6482 14884 6488
rect 14832 6424 14884 6430
rect 17222 6450 17278 6459
rect 14648 6278 14700 6284
rect 14648 6220 14700 6226
rect 14844 6187 14872 6424
rect 15956 6382 16252 6402
rect 17222 6385 17278 6394
rect 16012 6380 16036 6382
rect 16092 6380 16116 6382
rect 16172 6380 16196 6382
rect 16034 6328 16036 6380
rect 16098 6328 16110 6380
rect 16172 6328 16174 6380
rect 16012 6326 16036 6328
rect 16092 6326 16116 6328
rect 16172 6326 16196 6328
rect 15956 6306 16252 6326
rect 14830 6178 14886 6187
rect 14830 6113 14886 6122
rect 17236 6051 17264 6385
rect 12806 6042 12862 6051
rect 12806 5977 12862 5986
rect 17222 6042 17278 6051
rect 17222 5977 17278 5986
rect 12820 5740 12848 5977
rect 20956 5838 21252 5858
rect 21012 5836 21036 5838
rect 21092 5836 21116 5838
rect 21172 5836 21196 5838
rect 21034 5784 21036 5836
rect 21098 5784 21110 5836
rect 21172 5784 21174 5836
rect 21012 5782 21036 5784
rect 21092 5782 21116 5784
rect 21172 5782 21196 5784
rect 20956 5762 21252 5782
rect 12808 5734 12860 5740
rect 12808 5676 12860 5682
rect 12622 5634 12678 5643
rect 12622 5569 12624 5578
rect 12676 5569 12678 5578
rect 12624 5540 12676 5546
rect 12636 5196 12664 5540
rect 15956 5294 16252 5314
rect 16012 5292 16036 5294
rect 16092 5292 16116 5294
rect 16172 5292 16196 5294
rect 16034 5240 16036 5292
rect 16098 5240 16110 5292
rect 16172 5240 16174 5292
rect 16012 5238 16036 5240
rect 16092 5238 16116 5240
rect 16172 5238 16196 5240
rect 15956 5218 16252 5238
rect 16394 5226 16450 5235
rect 12624 5190 12676 5196
rect 16394 5161 16396 5170
rect 12624 5132 12676 5138
rect 16448 5161 16450 5170
rect 16396 5132 16448 5138
rect 13726 5090 13782 5099
rect 13726 5025 13782 5034
rect 13740 4992 13768 5025
rect 23584 4992 23612 16857
rect 23664 15730 23716 15736
rect 23664 15672 23716 15678
rect 23676 9451 23704 15672
rect 24032 15390 24084 15396
rect 24032 15332 24084 15338
rect 23938 15290 23994 15299
rect 23938 15225 23994 15234
rect 23756 15186 23808 15192
rect 23756 15128 23808 15134
rect 23662 9442 23718 9451
rect 23662 9377 23718 9386
rect 23768 8907 23796 15128
rect 23952 10516 23980 15225
rect 24044 14988 24072 15332
rect 24032 14982 24084 14988
rect 24032 14924 24084 14930
rect 24136 11491 24164 18392
rect 24216 17906 24268 17912
rect 24216 17848 24268 17854
rect 24228 13696 24256 17848
rect 24320 17572 24348 22841
rect 24398 22226 24454 22235
rect 24398 22161 24454 22170
rect 24308 17566 24360 17572
rect 24308 17508 24360 17514
rect 24320 17164 24348 17508
rect 24308 17158 24360 17164
rect 24308 17100 24360 17106
rect 24216 13690 24268 13696
rect 24216 13632 24268 13638
rect 24122 11482 24178 11491
rect 24122 11417 24178 11426
rect 24412 11044 24440 22161
rect 24858 21410 24914 21419
rect 24858 21345 24914 21354
rect 24490 21138 24546 21147
rect 24490 21073 24546 21082
rect 24504 16076 24532 21073
rect 24872 20632 24900 21345
rect 24860 20626 24912 20632
rect 24860 20568 24912 20574
rect 24858 20322 24914 20331
rect 24858 20257 24914 20266
rect 24676 18994 24728 19000
rect 24676 18936 24728 18942
rect 24582 17738 24638 17747
rect 24582 17673 24638 17682
rect 24492 16070 24544 16076
rect 24492 16012 24544 16018
rect 24504 15872 24532 16012
rect 24492 15866 24544 15872
rect 24492 15808 24544 15814
rect 24490 12298 24546 12307
rect 24490 12233 24546 12242
rect 24032 11038 24084 11044
rect 24032 10980 24084 10986
rect 24400 11038 24452 11044
rect 24400 10980 24452 10986
rect 24044 10636 24072 10980
rect 24124 10902 24176 10908
rect 24124 10844 24176 10850
rect 24032 10630 24084 10636
rect 24032 10572 24084 10578
rect 24136 10539 24164 10844
rect 24122 10530 24178 10539
rect 23952 10488 24072 10516
rect 23940 9338 23992 9344
rect 23938 9306 23940 9315
rect 23992 9306 23994 9315
rect 23938 9241 23994 9250
rect 23754 8898 23810 8907
rect 23754 8833 23810 8842
rect 23940 7774 23992 7780
rect 23940 7716 23992 7722
rect 23952 7168 23980 7716
rect 23940 7162 23992 7168
rect 23938 7130 23940 7139
rect 23992 7130 23994 7139
rect 23938 7065 23994 7074
rect 23940 6686 23992 6692
rect 23940 6628 23992 6634
rect 23952 6284 23980 6628
rect 23940 6278 23992 6284
rect 23940 6220 23992 6226
rect 13728 4986 13780 4992
rect 13728 4928 13780 4934
rect 23572 4986 23624 4992
rect 23572 4928 23624 4934
rect 20956 4750 21252 4770
rect 21012 4748 21036 4750
rect 21092 4748 21116 4750
rect 21172 4748 21196 4750
rect 21034 4696 21036 4748
rect 21098 4696 21110 4748
rect 21172 4696 21174 4748
rect 21012 4694 21036 4696
rect 21092 4694 21116 4696
rect 21172 4694 21196 4696
rect 20956 4674 21252 4694
rect 20718 4546 20774 4555
rect 16396 4510 16448 4516
rect 20718 4481 20720 4490
rect 16396 4452 16448 4458
rect 20772 4481 20774 4490
rect 20720 4452 20772 4458
rect 15956 4206 16252 4226
rect 16012 4204 16036 4206
rect 16092 4204 16116 4206
rect 16172 4204 16196 4206
rect 16034 4152 16036 4204
rect 16098 4152 16110 4204
rect 16172 4152 16174 4204
rect 16012 4150 16036 4152
rect 16092 4150 16116 4152
rect 16172 4150 16196 4152
rect 15956 4130 16252 4150
rect 16408 4040 16436 4452
rect 16486 4410 16542 4419
rect 16486 4345 16488 4354
rect 16540 4345 16542 4354
rect 16488 4316 16540 4322
rect 20732 4108 20760 4452
rect 20902 4410 20958 4419
rect 20902 4345 20904 4354
rect 20956 4345 20958 4354
rect 20904 4316 20956 4322
rect 20720 4102 20772 4108
rect 20720 4044 20772 4050
rect 16396 4034 16448 4040
rect 16394 4002 16396 4011
rect 16448 4002 16450 4011
rect 16394 3937 16450 3946
rect 23940 3898 23992 3904
rect 23938 3866 23940 3875
rect 23992 3866 23994 3875
rect 23938 3801 23994 3810
rect 21640 3762 21692 3768
rect 21640 3704 21692 3710
rect 22100 3762 22152 3768
rect 22100 3704 22152 3710
rect 20956 3662 21252 3682
rect 21012 3660 21036 3662
rect 21092 3660 21116 3662
rect 21172 3660 21196 3662
rect 21034 3608 21036 3660
rect 21098 3608 21110 3660
rect 21172 3608 21174 3660
rect 21012 3606 21036 3608
rect 21092 3606 21116 3608
rect 21172 3606 21196 3608
rect 20956 3586 21252 3606
rect 21652 3467 21680 3704
rect 22112 3603 22140 3704
rect 22098 3594 22154 3603
rect 22098 3529 22154 3538
rect 21638 3458 21694 3467
rect 24044 3428 24072 10488
rect 24122 10465 24178 10474
rect 24124 9202 24176 9208
rect 24122 9170 24124 9179
rect 24176 9170 24178 9179
rect 24122 9105 24178 9114
rect 24504 9020 24532 12233
rect 24320 8992 24532 9020
rect 24124 8658 24176 8664
rect 24124 8600 24176 8606
rect 24136 8363 24164 8600
rect 24122 8354 24178 8363
rect 24122 8289 24178 8298
rect 24122 7946 24178 7955
rect 24122 7881 24124 7890
rect 24176 7881 24178 7890
rect 24124 7852 24176 7858
rect 24320 7796 24348 8992
rect 24492 8862 24544 8868
rect 24492 8804 24544 8810
rect 24504 8256 24532 8804
rect 24596 8460 24624 17673
rect 24688 11899 24716 18936
rect 24872 18404 24900 20257
rect 24950 19914 25006 19923
rect 24950 19849 25006 19858
rect 24780 18376 24900 18404
rect 24780 15396 24808 18376
rect 24964 17747 24992 19849
rect 25056 18660 25084 23385
rect 26146 23346 26202 23826
rect 26160 21804 26188 23346
rect 25884 21776 26188 21804
rect 25884 19651 25912 21776
rect 25956 21614 26252 21634
rect 26012 21612 26036 21614
rect 26092 21612 26116 21614
rect 26172 21612 26196 21614
rect 26034 21560 26036 21612
rect 26098 21560 26110 21612
rect 26172 21560 26174 21612
rect 26012 21558 26036 21560
rect 26092 21558 26116 21560
rect 26172 21558 26196 21560
rect 25956 21538 26252 21558
rect 25956 20526 26252 20546
rect 26012 20524 26036 20526
rect 26092 20524 26116 20526
rect 26172 20524 26196 20526
rect 26034 20472 26036 20524
rect 26098 20472 26110 20524
rect 26172 20472 26174 20524
rect 26012 20470 26036 20472
rect 26092 20470 26116 20472
rect 26172 20470 26196 20472
rect 25956 20450 26252 20470
rect 25870 19642 25926 19651
rect 25870 19577 25926 19586
rect 25956 19438 26252 19458
rect 26012 19436 26036 19438
rect 26092 19436 26116 19438
rect 26172 19436 26196 19438
rect 26034 19384 26036 19436
rect 26098 19384 26110 19436
rect 26172 19384 26174 19436
rect 26012 19382 26036 19384
rect 26092 19382 26116 19384
rect 26172 19382 26196 19384
rect 25956 19362 26252 19382
rect 25594 19234 25650 19243
rect 25594 19169 25650 19178
rect 25226 18690 25282 18699
rect 25044 18654 25096 18660
rect 25226 18625 25282 18634
rect 25044 18596 25096 18602
rect 25056 18252 25084 18596
rect 25044 18246 25096 18252
rect 25044 18188 25096 18194
rect 24950 17738 25006 17747
rect 24950 17673 25006 17682
rect 24768 15390 24820 15396
rect 24768 15332 24820 15338
rect 24860 13894 24912 13900
rect 24860 13836 24912 13842
rect 24768 13690 24820 13696
rect 24768 13632 24820 13638
rect 24674 11890 24730 11899
rect 24674 11825 24730 11834
rect 24780 10947 24808 13632
rect 24872 12035 24900 13836
rect 25134 13250 25190 13259
rect 25134 13185 25190 13194
rect 24950 12162 25006 12171
rect 24950 12097 25006 12106
rect 24858 12026 24914 12035
rect 24858 11961 24914 11970
rect 24860 11650 24912 11656
rect 24860 11592 24912 11598
rect 24766 10938 24822 10947
rect 24766 10873 24822 10882
rect 24872 9859 24900 11592
rect 24964 10403 24992 12097
rect 25042 11890 25098 11899
rect 25042 11825 25098 11834
rect 24950 10394 25006 10403
rect 24950 10329 25006 10338
rect 25056 10267 25084 11825
rect 25148 11083 25176 13185
rect 25240 12307 25268 18625
rect 25320 18450 25372 18456
rect 25320 18392 25372 18398
rect 25332 13900 25360 18392
rect 25502 15698 25558 15707
rect 25502 15633 25558 15642
rect 25410 14474 25466 14483
rect 25410 14409 25466 14418
rect 25320 13894 25372 13900
rect 25320 13836 25372 13842
rect 25318 13794 25374 13803
rect 25318 13729 25374 13738
rect 25226 12298 25282 12307
rect 25226 12233 25282 12242
rect 25332 11627 25360 13729
rect 25424 11763 25452 14409
rect 25410 11754 25466 11763
rect 25410 11689 25466 11698
rect 25318 11618 25374 11627
rect 25318 11553 25374 11562
rect 25134 11074 25190 11083
rect 25134 11009 25190 11018
rect 25042 10258 25098 10267
rect 25042 10193 25098 10202
rect 24858 9850 24914 9859
rect 24858 9785 24914 9794
rect 24584 8454 24636 8460
rect 24584 8396 24636 8402
rect 24492 8250 24544 8256
rect 24490 8218 24492 8227
rect 24544 8218 24546 8227
rect 24490 8153 24546 8162
rect 24136 7768 24348 7796
rect 24136 6692 24164 7768
rect 24124 6686 24176 6692
rect 24124 6628 24176 6634
rect 24122 6586 24178 6595
rect 24122 6521 24124 6530
rect 24176 6521 24178 6530
rect 24124 6492 24176 6498
rect 24122 4954 24178 4963
rect 24122 4889 24178 4898
rect 24136 4856 24164 4889
rect 24124 4850 24176 4856
rect 24124 4792 24176 4798
rect 24124 3762 24176 3768
rect 24122 3730 24124 3739
rect 24176 3730 24178 3739
rect 24122 3665 24178 3674
rect 25516 3603 25544 15633
rect 25608 13667 25636 19169
rect 25956 18350 26252 18370
rect 26012 18348 26036 18350
rect 26092 18348 26116 18350
rect 26172 18348 26196 18350
rect 26034 18296 26036 18348
rect 26098 18296 26110 18348
rect 26172 18296 26174 18348
rect 26012 18294 26036 18296
rect 26092 18294 26116 18296
rect 26172 18294 26196 18296
rect 25956 18274 26252 18294
rect 25778 17466 25834 17475
rect 25778 17401 25834 17410
rect 25686 15970 25742 15979
rect 25686 15905 25742 15914
rect 25594 13658 25650 13667
rect 25594 13593 25650 13602
rect 25594 12706 25650 12715
rect 25594 12641 25650 12650
rect 25502 3594 25558 3603
rect 25502 3529 25558 3538
rect 21638 3393 21694 3402
rect 24032 3422 24084 3428
rect 24032 3364 24084 3370
rect 15956 3118 16252 3138
rect 16012 3116 16036 3118
rect 16092 3116 16116 3118
rect 16172 3116 16196 3118
rect 16034 3064 16036 3116
rect 16098 3064 16110 3116
rect 16172 3064 16174 3116
rect 16012 3062 16036 3064
rect 16092 3062 16116 3064
rect 16172 3062 16196 3064
rect 15956 3042 16252 3062
rect 24044 3020 24072 3364
rect 24122 3322 24178 3331
rect 24122 3257 24124 3266
rect 24176 3257 24178 3266
rect 24124 3228 24176 3234
rect 24032 3014 24084 3020
rect 24032 2956 24084 2962
rect 23938 2914 23994 2923
rect 23938 2849 23994 2858
rect 23952 2816 23980 2849
rect 23940 2810 23992 2816
rect 23940 2752 23992 2758
rect 24860 2674 24912 2680
rect 24860 2616 24912 2622
rect 20956 2574 21252 2594
rect 21012 2572 21036 2574
rect 21092 2572 21116 2574
rect 21172 2572 21196 2574
rect 21034 2520 21036 2572
rect 21098 2520 21110 2572
rect 21172 2520 21174 2572
rect 21012 2518 21036 2520
rect 21092 2518 21116 2520
rect 21172 2518 21196 2520
rect 20956 2498 21252 2518
rect 24214 2506 24270 2515
rect 24214 2441 24216 2450
rect 24268 2441 24270 2450
rect 24216 2412 24268 2418
rect 24032 2334 24084 2340
rect 24032 2276 24084 2282
rect 24044 2243 24072 2276
rect 12530 2234 12586 2243
rect 12530 2169 12586 2178
rect 24030 2234 24086 2243
rect 24030 2169 24086 2178
rect 15956 2030 16252 2050
rect 16012 2028 16036 2030
rect 16092 2028 16116 2030
rect 16172 2028 16196 2030
rect 16034 1976 16036 2028
rect 16098 1976 16110 2028
rect 16172 1976 16174 2028
rect 16012 1974 16036 1976
rect 16092 1974 16116 1976
rect 16172 1974 16196 1976
rect 15956 1954 16252 1974
rect 8390 1826 8446 1835
rect 8390 1761 8446 1770
rect 24872 1427 24900 2616
rect 25608 2379 25636 12641
rect 25700 4011 25728 15905
rect 25792 5643 25820 17401
rect 25956 17262 26252 17282
rect 26012 17260 26036 17262
rect 26092 17260 26116 17262
rect 26172 17260 26196 17262
rect 26034 17208 26036 17260
rect 26098 17208 26110 17260
rect 26172 17208 26174 17260
rect 26012 17206 26036 17208
rect 26092 17206 26116 17208
rect 26172 17206 26196 17208
rect 25956 17186 26252 17206
rect 25956 16174 26252 16194
rect 26012 16172 26036 16174
rect 26092 16172 26116 16174
rect 26172 16172 26196 16174
rect 26034 16120 26036 16172
rect 26098 16120 26110 16172
rect 26172 16120 26174 16172
rect 26012 16118 26036 16120
rect 26092 16118 26116 16120
rect 26172 16118 26196 16120
rect 25956 16098 26252 16118
rect 25956 15086 26252 15106
rect 26012 15084 26036 15086
rect 26092 15084 26116 15086
rect 26172 15084 26196 15086
rect 26034 15032 26036 15084
rect 26098 15032 26110 15084
rect 26172 15032 26174 15084
rect 26012 15030 26036 15032
rect 26092 15030 26116 15032
rect 26172 15030 26196 15032
rect 25956 15010 26252 15030
rect 25956 13998 26252 14018
rect 26012 13996 26036 13998
rect 26092 13996 26116 13998
rect 26172 13996 26196 13998
rect 26034 13944 26036 13996
rect 26098 13944 26110 13996
rect 26172 13944 26174 13996
rect 26012 13942 26036 13944
rect 26092 13942 26116 13944
rect 26172 13942 26196 13944
rect 25956 13922 26252 13942
rect 25956 12910 26252 12930
rect 26012 12908 26036 12910
rect 26092 12908 26116 12910
rect 26172 12908 26196 12910
rect 26034 12856 26036 12908
rect 26098 12856 26110 12908
rect 26172 12856 26174 12908
rect 26012 12854 26036 12856
rect 26092 12854 26116 12856
rect 26172 12854 26196 12856
rect 25956 12834 26252 12854
rect 25956 11822 26252 11842
rect 26012 11820 26036 11822
rect 26092 11820 26116 11822
rect 26172 11820 26196 11822
rect 26034 11768 26036 11820
rect 26098 11768 26110 11820
rect 26172 11768 26174 11820
rect 26012 11766 26036 11768
rect 26092 11766 26116 11768
rect 26172 11766 26196 11768
rect 25956 11746 26252 11766
rect 25956 10734 26252 10754
rect 26012 10732 26036 10734
rect 26092 10732 26116 10734
rect 26172 10732 26196 10734
rect 26034 10680 26036 10732
rect 26098 10680 26110 10732
rect 26172 10680 26174 10732
rect 26012 10678 26036 10680
rect 26092 10678 26116 10680
rect 26172 10678 26196 10680
rect 25956 10658 26252 10678
rect 25956 9646 26252 9666
rect 26012 9644 26036 9646
rect 26092 9644 26116 9646
rect 26172 9644 26196 9646
rect 26034 9592 26036 9644
rect 26098 9592 26110 9644
rect 26172 9592 26174 9644
rect 26012 9590 26036 9592
rect 26092 9590 26116 9592
rect 26172 9590 26196 9592
rect 25956 9570 26252 9590
rect 25956 8558 26252 8578
rect 26012 8556 26036 8558
rect 26092 8556 26116 8558
rect 26172 8556 26196 8558
rect 26034 8504 26036 8556
rect 26098 8504 26110 8556
rect 26172 8504 26174 8556
rect 26012 8502 26036 8504
rect 26092 8502 26116 8504
rect 26172 8502 26196 8504
rect 25956 8482 26252 8502
rect 25956 7470 26252 7490
rect 26012 7468 26036 7470
rect 26092 7468 26116 7470
rect 26172 7468 26196 7470
rect 26034 7416 26036 7468
rect 26098 7416 26110 7468
rect 26172 7416 26174 7468
rect 26012 7414 26036 7416
rect 26092 7414 26116 7416
rect 26172 7414 26196 7416
rect 25956 7394 26252 7414
rect 25956 6382 26252 6402
rect 26012 6380 26036 6382
rect 26092 6380 26116 6382
rect 26172 6380 26196 6382
rect 26034 6328 26036 6380
rect 26098 6328 26110 6380
rect 26172 6328 26174 6380
rect 26012 6326 26036 6328
rect 26092 6326 26116 6328
rect 26172 6326 26196 6328
rect 25956 6306 26252 6326
rect 25778 5634 25834 5643
rect 25778 5569 25834 5578
rect 25956 5294 26252 5314
rect 26012 5292 26036 5294
rect 26092 5292 26116 5294
rect 26172 5292 26196 5294
rect 26034 5240 26036 5292
rect 26098 5240 26110 5292
rect 26172 5240 26174 5292
rect 26012 5238 26036 5240
rect 26092 5238 26116 5240
rect 26172 5238 26196 5240
rect 25956 5218 26252 5238
rect 25956 4206 26252 4226
rect 26012 4204 26036 4206
rect 26092 4204 26116 4206
rect 26172 4204 26196 4206
rect 26034 4152 26036 4204
rect 26098 4152 26110 4204
rect 26172 4152 26174 4204
rect 26012 4150 26036 4152
rect 26092 4150 26116 4152
rect 26172 4150 26196 4152
rect 25956 4130 26252 4150
rect 25686 4002 25742 4011
rect 25686 3937 25742 3946
rect 25956 3118 26252 3138
rect 26012 3116 26036 3118
rect 26092 3116 26116 3118
rect 26172 3116 26196 3118
rect 26034 3064 26036 3116
rect 26098 3064 26110 3116
rect 26172 3064 26174 3116
rect 26012 3062 26036 3064
rect 26092 3062 26116 3064
rect 26172 3062 26196 3064
rect 25956 3042 26252 3062
rect 25594 2370 25650 2379
rect 25136 2334 25188 2340
rect 25594 2305 25650 2314
rect 25136 2276 25188 2282
rect 25148 1835 25176 2276
rect 25320 2130 25372 2136
rect 25320 2072 25372 2078
rect 25134 1826 25190 1835
rect 25134 1761 25190 1770
rect 24858 1418 24914 1427
rect 24858 1353 24914 1362
rect 25332 203 25360 2072
rect 25956 2030 26252 2050
rect 26012 2028 26036 2030
rect 26092 2028 26116 2030
rect 26172 2028 26196 2030
rect 26034 1976 26036 2028
rect 26098 1976 26110 2028
rect 26172 1976 26174 2028
rect 26012 1974 26036 1976
rect 26092 1974 26116 1976
rect 26172 1974 26196 1976
rect 25956 1954 26252 1974
rect 1490 194 1546 203
rect 1490 129 1546 138
rect 2686 194 2742 203
rect 2686 129 2742 138
rect 25318 194 25374 203
rect 25318 129 25374 138
<< via2 >>
rect 3882 23394 3938 23450
rect 3054 22850 3110 22906
rect 3330 22170 3386 22226
rect 3422 21626 3478 21682
rect 3514 21082 3570 21138
rect 3422 19178 3478 19234
rect 3330 19042 3386 19098
rect 3146 18634 3202 18690
rect 3054 17954 3110 18010
rect 2962 15642 3018 15698
rect 1398 15098 1454 15154
rect 1674 13874 1730 13930
rect 1490 13214 1546 13250
rect 1490 13194 1492 13214
rect 1492 13194 1544 13214
rect 1544 13194 1546 13214
rect 1398 9930 1454 9986
rect 1858 12650 1914 12706
rect 1582 9694 1584 9714
rect 1584 9694 1636 9714
rect 1636 9694 1638 9714
rect 1582 9658 1638 9694
rect 2042 11038 2098 11074
rect 2042 11018 2044 11038
rect 2044 11018 2096 11038
rect 2096 11018 2098 11038
rect 2042 9794 2098 9850
rect 2134 6122 2190 6178
rect 1858 2722 1914 2778
rect 1766 2450 1822 2506
rect 2042 2334 2098 2370
rect 2042 2314 2044 2334
rect 2044 2314 2096 2334
rect 2096 2314 2098 2334
rect 1950 1906 2006 1962
rect 2410 11290 2466 11346
rect 2502 11154 2558 11210
rect 3238 18090 3294 18146
rect 3146 13058 3202 13114
rect 3790 19858 3846 19914
rect 3698 18634 3754 18690
rect 3330 17410 3386 17466
rect 3238 12514 3294 12570
rect 3146 11970 3202 12026
rect 3514 16866 3570 16922
rect 3422 14418 3478 14474
rect 3422 13058 3478 13114
rect 3422 11562 3478 11618
rect 3422 10882 3478 10938
rect 3330 8978 3386 9034
rect 3054 8026 3110 8082
rect 3606 12106 3662 12162
rect 3606 10066 3662 10122
rect 3698 9250 3754 9306
rect 3606 8026 3662 8082
rect 3698 7754 3754 7810
rect 3606 7618 3662 7674
rect 3698 7210 3754 7266
rect 25042 23394 25098 23450
rect 5956 21612 6012 21614
rect 6036 21612 6092 21614
rect 6116 21612 6172 21614
rect 6196 21612 6252 21614
rect 5956 21560 5982 21612
rect 5982 21560 6012 21612
rect 6036 21560 6046 21612
rect 6046 21560 6092 21612
rect 6116 21560 6162 21612
rect 6162 21560 6172 21612
rect 6196 21560 6226 21612
rect 6226 21560 6252 21612
rect 5956 21558 6012 21560
rect 6036 21558 6092 21560
rect 6116 21558 6172 21560
rect 6196 21558 6252 21560
rect 15956 21612 16012 21614
rect 16036 21612 16092 21614
rect 16116 21612 16172 21614
rect 16196 21612 16252 21614
rect 15956 21560 15982 21612
rect 15982 21560 16012 21612
rect 16036 21560 16046 21612
rect 16046 21560 16092 21612
rect 16116 21560 16162 21612
rect 16162 21560 16172 21612
rect 16196 21560 16226 21612
rect 16226 21560 16252 21612
rect 15956 21558 16012 21560
rect 16036 21558 16092 21560
rect 16116 21558 16172 21560
rect 16196 21558 16252 21560
rect 10956 21068 11012 21070
rect 11036 21068 11092 21070
rect 11116 21068 11172 21070
rect 11196 21068 11252 21070
rect 10956 21016 10982 21068
rect 10982 21016 11012 21068
rect 11036 21016 11046 21068
rect 11046 21016 11092 21068
rect 11116 21016 11162 21068
rect 11162 21016 11172 21068
rect 11196 21016 11226 21068
rect 11226 21016 11252 21068
rect 10956 21014 11012 21016
rect 11036 21014 11092 21016
rect 11116 21014 11172 21016
rect 11196 21014 11252 21016
rect 5956 20524 6012 20526
rect 6036 20524 6092 20526
rect 6116 20524 6172 20526
rect 6196 20524 6252 20526
rect 5956 20472 5982 20524
rect 5982 20472 6012 20524
rect 6036 20472 6046 20524
rect 6046 20472 6092 20524
rect 6116 20472 6162 20524
rect 6162 20472 6172 20524
rect 6196 20472 6226 20524
rect 6226 20472 6252 20524
rect 5956 20470 6012 20472
rect 6036 20470 6092 20472
rect 6116 20470 6172 20472
rect 6196 20470 6252 20472
rect 3974 20402 4030 20458
rect 3882 18090 3938 18146
rect 10956 19980 11012 19982
rect 11036 19980 11092 19982
rect 11116 19980 11172 19982
rect 11196 19980 11252 19982
rect 10956 19928 10982 19980
rect 10982 19928 11012 19980
rect 11036 19928 11046 19980
rect 11046 19928 11092 19980
rect 11116 19928 11162 19980
rect 11162 19928 11172 19980
rect 11196 19928 11226 19980
rect 11226 19928 11252 19980
rect 10956 19926 11012 19928
rect 11036 19926 11092 19928
rect 11116 19926 11172 19928
rect 11196 19926 11252 19928
rect 5956 19436 6012 19438
rect 6036 19436 6092 19438
rect 6116 19436 6172 19438
rect 6196 19436 6252 19438
rect 5956 19384 5982 19436
rect 5982 19384 6012 19436
rect 6036 19384 6046 19436
rect 6046 19384 6092 19436
rect 6116 19384 6162 19436
rect 6162 19384 6172 19436
rect 6196 19384 6226 19436
rect 6226 19384 6252 19436
rect 5956 19382 6012 19384
rect 6036 19382 6092 19384
rect 6116 19382 6172 19384
rect 6196 19382 6252 19384
rect 15956 20524 16012 20526
rect 16036 20524 16092 20526
rect 16116 20524 16172 20526
rect 16196 20524 16252 20526
rect 15956 20472 15982 20524
rect 15982 20472 16012 20524
rect 16036 20472 16046 20524
rect 16046 20472 16092 20524
rect 16116 20472 16162 20524
rect 16162 20472 16172 20524
rect 16196 20472 16226 20524
rect 16226 20472 16252 20524
rect 15956 20470 16012 20472
rect 16036 20470 16092 20472
rect 16116 20470 16172 20472
rect 16196 20470 16252 20472
rect 15956 19436 16012 19438
rect 16036 19436 16092 19438
rect 16116 19436 16172 19438
rect 16196 19436 16252 19438
rect 15956 19384 15982 19436
rect 15982 19384 16012 19436
rect 16036 19384 16046 19436
rect 16046 19384 16092 19436
rect 16116 19384 16162 19436
rect 16162 19384 16172 19436
rect 16196 19384 16226 19436
rect 16226 19384 16252 19436
rect 15956 19382 16012 19384
rect 16036 19382 16092 19384
rect 16116 19382 16172 19384
rect 16196 19382 16252 19384
rect 8850 19178 8906 19234
rect 11334 19178 11390 19234
rect 10956 18892 11012 18894
rect 11036 18892 11092 18894
rect 11116 18892 11172 18894
rect 11196 18892 11252 18894
rect 10956 18840 10982 18892
rect 10982 18840 11012 18892
rect 11036 18840 11046 18892
rect 11046 18840 11092 18892
rect 11116 18840 11162 18892
rect 11162 18840 11172 18892
rect 11196 18840 11226 18892
rect 11226 18840 11252 18892
rect 10956 18838 11012 18840
rect 11036 18838 11092 18840
rect 11116 18838 11172 18840
rect 11196 18838 11252 18840
rect 24306 22850 24362 22906
rect 20956 21068 21012 21070
rect 21036 21068 21092 21070
rect 21116 21068 21172 21070
rect 21196 21068 21252 21070
rect 20956 21016 20982 21068
rect 20982 21016 21012 21068
rect 21036 21016 21046 21068
rect 21046 21016 21092 21068
rect 21116 21016 21162 21068
rect 21162 21016 21172 21068
rect 21196 21016 21226 21068
rect 21226 21016 21252 21068
rect 20956 21014 21012 21016
rect 21036 21014 21092 21016
rect 21116 21014 21172 21016
rect 21196 21014 21252 21016
rect 16670 18790 16726 18826
rect 16670 18770 16672 18790
rect 16672 18770 16724 18790
rect 16724 18770 16726 18790
rect 18694 18770 18750 18826
rect 7010 18634 7066 18690
rect 8574 18654 8630 18690
rect 8574 18634 8576 18654
rect 8576 18634 8628 18654
rect 8628 18634 8630 18654
rect 5956 18348 6012 18350
rect 6036 18348 6092 18350
rect 6116 18348 6172 18350
rect 6196 18348 6252 18350
rect 5956 18296 5982 18348
rect 5982 18296 6012 18348
rect 6036 18296 6046 18348
rect 6046 18296 6092 18348
rect 6116 18296 6162 18348
rect 6162 18296 6172 18348
rect 6196 18296 6226 18348
rect 6226 18296 6252 18348
rect 5956 18294 6012 18296
rect 6036 18294 6092 18296
rect 6116 18294 6172 18296
rect 6196 18294 6252 18296
rect 5956 17260 6012 17262
rect 6036 17260 6092 17262
rect 6116 17260 6172 17262
rect 6196 17260 6252 17262
rect 5956 17208 5982 17260
rect 5982 17208 6012 17260
rect 6036 17208 6046 17260
rect 6046 17208 6092 17260
rect 6116 17208 6162 17260
rect 6162 17208 6172 17260
rect 6196 17208 6226 17260
rect 6226 17208 6252 17260
rect 5956 17206 6012 17208
rect 6036 17206 6092 17208
rect 6116 17206 6172 17208
rect 6196 17206 6252 17208
rect 4066 16186 4122 16242
rect 3974 8162 4030 8218
rect 3882 7210 3938 7266
rect 3790 7074 3846 7130
rect 5956 16172 6012 16174
rect 6036 16172 6092 16174
rect 6116 16172 6172 16174
rect 6196 16172 6252 16174
rect 5956 16120 5982 16172
rect 5982 16120 6012 16172
rect 6036 16120 6046 16172
rect 6046 16120 6092 16172
rect 6116 16120 6162 16172
rect 6162 16120 6172 16172
rect 6196 16120 6226 16172
rect 6226 16120 6252 16172
rect 5956 16118 6012 16120
rect 6036 16118 6092 16120
rect 6116 16118 6172 16120
rect 6196 16118 6252 16120
rect 12990 18634 13046 18690
rect 10956 17804 11012 17806
rect 11036 17804 11092 17806
rect 11116 17804 11172 17806
rect 11196 17804 11252 17806
rect 10956 17752 10982 17804
rect 10982 17752 11012 17804
rect 11036 17752 11046 17804
rect 11046 17752 11092 17804
rect 11116 17752 11162 17804
rect 11162 17752 11172 17804
rect 11196 17752 11226 17804
rect 11226 17752 11252 17804
rect 10956 17750 11012 17752
rect 11036 17750 11092 17752
rect 11116 17750 11172 17752
rect 11196 17750 11252 17752
rect 10956 16716 11012 16718
rect 11036 16716 11092 16718
rect 11116 16716 11172 16718
rect 11196 16716 11252 16718
rect 10956 16664 10982 16716
rect 10982 16664 11012 16716
rect 11036 16664 11046 16716
rect 11046 16664 11092 16716
rect 11116 16664 11162 16716
rect 11162 16664 11172 16716
rect 11196 16664 11226 16716
rect 11226 16664 11252 16716
rect 10956 16662 11012 16664
rect 11036 16662 11092 16664
rect 11116 16662 11172 16664
rect 11196 16662 11252 16664
rect 15290 18634 15346 18690
rect 15956 18348 16012 18350
rect 16036 18348 16092 18350
rect 16116 18348 16172 18350
rect 16196 18348 16252 18350
rect 15956 18296 15982 18348
rect 15982 18296 16012 18348
rect 16036 18296 16046 18348
rect 16046 18296 16092 18348
rect 16116 18296 16162 18348
rect 16162 18296 16172 18348
rect 16196 18296 16226 18348
rect 16226 18296 16252 18348
rect 15956 18294 16012 18296
rect 16036 18294 16092 18296
rect 16116 18294 16172 18296
rect 16196 18294 16252 18296
rect 13542 16730 13598 16786
rect 7194 15798 7250 15834
rect 7194 15778 7196 15798
rect 7196 15778 7248 15798
rect 7248 15778 7250 15798
rect 9954 15778 10010 15834
rect 5956 15084 6012 15086
rect 6036 15084 6092 15086
rect 6116 15084 6172 15086
rect 6196 15084 6252 15086
rect 5956 15032 5982 15084
rect 5982 15032 6012 15084
rect 6036 15032 6046 15084
rect 6046 15032 6092 15084
rect 6116 15032 6162 15084
rect 6162 15032 6172 15084
rect 6196 15032 6226 15084
rect 6226 15032 6252 15084
rect 5956 15030 6012 15032
rect 6036 15030 6092 15032
rect 6116 15030 6172 15032
rect 6196 15030 6252 15032
rect 5956 13996 6012 13998
rect 6036 13996 6092 13998
rect 6116 13996 6172 13998
rect 6196 13996 6252 13998
rect 5956 13944 5982 13996
rect 5982 13944 6012 13996
rect 6036 13944 6046 13996
rect 6046 13944 6092 13996
rect 6116 13944 6162 13996
rect 6162 13944 6172 13996
rect 6196 13944 6226 13996
rect 6226 13944 6252 13996
rect 5956 13942 6012 13944
rect 6036 13942 6092 13944
rect 6116 13942 6172 13944
rect 6196 13942 6252 13944
rect 5956 12908 6012 12910
rect 6036 12908 6092 12910
rect 6116 12908 6172 12910
rect 6196 12908 6252 12910
rect 5956 12856 5982 12908
rect 5982 12856 6012 12908
rect 6036 12856 6046 12908
rect 6046 12856 6092 12908
rect 6116 12856 6162 12908
rect 6162 12856 6172 12908
rect 6196 12856 6226 12908
rect 6226 12856 6252 12908
rect 5956 12854 6012 12856
rect 6036 12854 6092 12856
rect 6116 12854 6172 12856
rect 6196 12854 6252 12856
rect 5956 11820 6012 11822
rect 6036 11820 6092 11822
rect 6116 11820 6172 11822
rect 6196 11820 6252 11822
rect 5956 11768 5982 11820
rect 5982 11768 6012 11820
rect 6036 11768 6046 11820
rect 6046 11768 6092 11820
rect 6116 11768 6162 11820
rect 6162 11768 6172 11820
rect 6196 11768 6226 11820
rect 6226 11768 6252 11820
rect 5956 11766 6012 11768
rect 6036 11766 6092 11768
rect 6116 11766 6172 11768
rect 6196 11766 6252 11768
rect 6642 11562 6698 11618
rect 6642 11290 6698 11346
rect 7102 11154 7158 11210
rect 5956 10732 6012 10734
rect 6036 10732 6092 10734
rect 6116 10732 6172 10734
rect 6196 10732 6252 10734
rect 5956 10680 5982 10732
rect 5982 10680 6012 10732
rect 6036 10680 6046 10732
rect 6046 10680 6092 10732
rect 6116 10680 6162 10732
rect 6162 10680 6172 10732
rect 6196 10680 6226 10732
rect 6226 10680 6252 10732
rect 5956 10678 6012 10680
rect 6036 10678 6092 10680
rect 6116 10678 6172 10680
rect 6196 10678 6252 10680
rect 10956 15628 11012 15630
rect 11036 15628 11092 15630
rect 11116 15628 11172 15630
rect 11196 15628 11252 15630
rect 10956 15576 10982 15628
rect 10982 15576 11012 15628
rect 11036 15576 11046 15628
rect 11046 15576 11092 15628
rect 11116 15576 11162 15628
rect 11162 15576 11172 15628
rect 11196 15576 11226 15628
rect 11226 15576 11252 15628
rect 10956 15574 11012 15576
rect 11036 15574 11092 15576
rect 11116 15574 11172 15576
rect 11196 15574 11252 15576
rect 10956 14540 11012 14542
rect 11036 14540 11092 14542
rect 11116 14540 11172 14542
rect 11196 14540 11252 14542
rect 10956 14488 10982 14540
rect 10982 14488 11012 14540
rect 11036 14488 11046 14540
rect 11046 14488 11092 14540
rect 11116 14488 11162 14540
rect 11162 14488 11172 14540
rect 11196 14488 11226 14540
rect 11226 14488 11252 14540
rect 10956 14486 11012 14488
rect 11036 14486 11092 14488
rect 11116 14486 11172 14488
rect 11196 14486 11252 14488
rect 10956 13452 11012 13454
rect 11036 13452 11092 13454
rect 11116 13452 11172 13454
rect 11196 13452 11252 13454
rect 10956 13400 10982 13452
rect 10982 13400 11012 13452
rect 11036 13400 11046 13452
rect 11046 13400 11092 13452
rect 11116 13400 11162 13452
rect 11162 13400 11172 13452
rect 11196 13400 11226 13452
rect 11226 13400 11252 13452
rect 10956 13398 11012 13400
rect 11036 13398 11092 13400
rect 11116 13398 11172 13400
rect 11196 13398 11252 13400
rect 15956 17260 16012 17262
rect 16036 17260 16092 17262
rect 16116 17260 16172 17262
rect 16196 17260 16252 17262
rect 15956 17208 15982 17260
rect 15982 17208 16012 17260
rect 16036 17208 16046 17260
rect 16046 17208 16092 17260
rect 16116 17208 16162 17260
rect 16162 17208 16172 17260
rect 16196 17208 16226 17260
rect 16226 17208 16252 17260
rect 15956 17206 16012 17208
rect 16036 17206 16092 17208
rect 16116 17206 16172 17208
rect 16196 17206 16252 17208
rect 17498 16766 17500 16786
rect 17500 16766 17552 16786
rect 17552 16766 17554 16786
rect 17498 16730 17554 16766
rect 11886 13058 11942 13114
rect 10956 12364 11012 12366
rect 11036 12364 11092 12366
rect 11116 12364 11172 12366
rect 11196 12364 11252 12366
rect 10956 12312 10982 12364
rect 10982 12312 11012 12364
rect 11036 12312 11046 12364
rect 11046 12312 11092 12364
rect 11116 12312 11162 12364
rect 11162 12312 11172 12364
rect 11196 12312 11226 12364
rect 11226 12312 11252 12364
rect 10956 12310 11012 12312
rect 11036 12310 11092 12312
rect 11116 12310 11172 12312
rect 11196 12310 11252 12312
rect 7378 11970 7434 12026
rect 7930 11990 7986 12026
rect 7930 11970 7932 11990
rect 7932 11970 7984 11990
rect 7984 11970 7986 11990
rect 8390 11834 8446 11890
rect 8114 10882 8170 10938
rect 12898 12550 12900 12570
rect 12900 12550 12952 12570
rect 12952 12550 12954 12570
rect 12898 12514 12954 12550
rect 15956 16172 16012 16174
rect 16036 16172 16092 16174
rect 16116 16172 16172 16174
rect 16196 16172 16252 16174
rect 15956 16120 15982 16172
rect 15982 16120 16012 16172
rect 16036 16120 16046 16172
rect 16046 16120 16092 16172
rect 16116 16120 16162 16172
rect 16162 16120 16172 16172
rect 16196 16120 16226 16172
rect 16226 16120 16252 16172
rect 15956 16118 16012 16120
rect 16036 16118 16092 16120
rect 16116 16118 16172 16120
rect 16196 16118 16252 16120
rect 15956 15084 16012 15086
rect 16036 15084 16092 15086
rect 16116 15084 16172 15086
rect 16196 15084 16252 15086
rect 15956 15032 15982 15084
rect 15982 15032 16012 15084
rect 16036 15032 16046 15084
rect 16046 15032 16092 15084
rect 16116 15032 16162 15084
rect 16162 15032 16172 15084
rect 16196 15032 16226 15084
rect 16226 15032 16252 15084
rect 15956 15030 16012 15032
rect 16036 15030 16092 15032
rect 16116 15030 16172 15032
rect 16196 15030 16252 15032
rect 14186 14826 14242 14882
rect 18326 14846 18382 14882
rect 18326 14826 18328 14846
rect 18328 14826 18380 14846
rect 18380 14826 18382 14846
rect 12070 11870 12072 11890
rect 12072 11870 12124 11890
rect 12124 11870 12126 11890
rect 12070 11834 12126 11870
rect 11518 11562 11574 11618
rect 13726 12142 13728 12162
rect 13728 12142 13780 12162
rect 13780 12142 13782 12162
rect 13726 12106 13782 12142
rect 15956 13996 16012 13998
rect 16036 13996 16092 13998
rect 16116 13996 16172 13998
rect 16196 13996 16252 13998
rect 15956 13944 15982 13996
rect 15982 13944 16012 13996
rect 16036 13944 16046 13996
rect 16046 13944 16092 13996
rect 16116 13944 16162 13996
rect 16162 13944 16172 13996
rect 16196 13944 16226 13996
rect 16226 13944 16252 13996
rect 15956 13942 16012 13944
rect 16036 13942 16092 13944
rect 16116 13942 16172 13944
rect 16196 13942 16252 13944
rect 19890 18226 19946 18282
rect 19890 13194 19946 13250
rect 19614 13058 19670 13114
rect 15956 12908 16012 12910
rect 16036 12908 16092 12910
rect 16116 12908 16172 12910
rect 16196 12908 16252 12910
rect 15956 12856 15982 12908
rect 15982 12856 16012 12908
rect 16036 12856 16046 12908
rect 16046 12856 16092 12908
rect 16116 12856 16162 12908
rect 16162 12856 16172 12908
rect 16196 12856 16226 12908
rect 16226 12856 16252 12908
rect 15956 12854 16012 12856
rect 16036 12854 16092 12856
rect 16116 12854 16172 12856
rect 16196 12854 16252 12856
rect 14646 12514 14702 12570
rect 13818 11970 13874 12026
rect 10956 11276 11012 11278
rect 11036 11276 11092 11278
rect 11116 11276 11172 11278
rect 11196 11276 11252 11278
rect 10956 11224 10982 11276
rect 10982 11224 11012 11276
rect 11036 11224 11046 11276
rect 11046 11224 11092 11276
rect 11116 11224 11162 11276
rect 11162 11224 11172 11276
rect 11196 11224 11226 11276
rect 11226 11224 11252 11276
rect 10956 11222 11012 11224
rect 11036 11222 11092 11224
rect 11116 11222 11172 11224
rect 11196 11222 11252 11224
rect 13726 11446 13782 11482
rect 13726 11426 13728 11446
rect 13728 11426 13780 11446
rect 13780 11426 13782 11446
rect 12438 11154 12494 11210
rect 12438 10882 12494 10938
rect 8298 10358 8354 10394
rect 8298 10338 8300 10358
rect 8300 10338 8352 10358
rect 8352 10338 8354 10358
rect 5956 9644 6012 9646
rect 6036 9644 6092 9646
rect 6116 9644 6172 9646
rect 6196 9644 6252 9646
rect 5956 9592 5982 9644
rect 5982 9592 6012 9644
rect 6036 9592 6046 9644
rect 6046 9592 6092 9644
rect 6116 9592 6162 9644
rect 6162 9592 6172 9644
rect 6196 9592 6226 9644
rect 6226 9592 6252 9644
rect 5956 9590 6012 9592
rect 6036 9590 6092 9592
rect 6116 9590 6172 9592
rect 6196 9590 6252 9592
rect 4802 8978 4858 9034
rect 3514 5034 3570 5090
rect 5956 8556 6012 8558
rect 6036 8556 6092 8558
rect 6116 8556 6172 8558
rect 6196 8556 6252 8558
rect 5956 8504 5982 8556
rect 5982 8504 6012 8556
rect 6036 8504 6046 8556
rect 6046 8504 6092 8556
rect 6116 8504 6162 8556
rect 6162 8504 6172 8556
rect 6196 8504 6226 8556
rect 6226 8504 6252 8556
rect 5956 8502 6012 8504
rect 6036 8502 6092 8504
rect 6116 8502 6172 8504
rect 6196 8502 6252 8504
rect 5956 7468 6012 7470
rect 6036 7468 6092 7470
rect 6116 7468 6172 7470
rect 6196 7468 6252 7470
rect 5956 7416 5982 7468
rect 5982 7416 6012 7468
rect 6036 7416 6046 7468
rect 6046 7416 6092 7468
rect 6116 7416 6162 7468
rect 6162 7416 6172 7468
rect 6196 7416 6226 7468
rect 6226 7416 6252 7468
rect 5956 7414 6012 7416
rect 6036 7414 6092 7416
rect 6116 7414 6172 7416
rect 6196 7414 6252 7416
rect 5956 6380 6012 6382
rect 6036 6380 6092 6382
rect 6116 6380 6172 6382
rect 6196 6380 6252 6382
rect 5956 6328 5982 6380
rect 5982 6328 6012 6380
rect 6036 6328 6046 6380
rect 6046 6328 6092 6380
rect 6116 6328 6162 6380
rect 6162 6328 6172 6380
rect 6196 6328 6226 6380
rect 6226 6328 6252 6380
rect 5956 6326 6012 6328
rect 6036 6326 6092 6328
rect 6116 6326 6172 6328
rect 6196 6326 6252 6328
rect 4986 5462 5042 5498
rect 4986 5442 4988 5462
rect 4988 5442 5040 5462
rect 5040 5442 5042 5462
rect 5956 5292 6012 5294
rect 6036 5292 6092 5294
rect 6116 5292 6172 5294
rect 6196 5292 6252 5294
rect 5956 5240 5982 5292
rect 5982 5240 6012 5292
rect 6036 5240 6046 5292
rect 6046 5240 6092 5292
rect 6116 5240 6162 5292
rect 6162 5240 6172 5292
rect 6196 5240 6226 5292
rect 6226 5240 6252 5292
rect 5956 5238 6012 5240
rect 6036 5238 6092 5240
rect 6116 5238 6172 5240
rect 6196 5238 6252 5240
rect 3882 4490 3938 4546
rect 5956 4204 6012 4206
rect 6036 4204 6092 4206
rect 6116 4204 6172 4206
rect 6196 4204 6252 4206
rect 5956 4152 5982 4204
rect 5982 4152 6012 4204
rect 6036 4152 6046 4204
rect 6046 4152 6092 4204
rect 6116 4152 6162 4204
rect 6162 4152 6172 4204
rect 6196 4152 6226 4204
rect 6226 4152 6252 4204
rect 5956 4150 6012 4152
rect 6036 4150 6092 4152
rect 6116 4150 6172 4152
rect 6196 4150 6252 4152
rect 3422 3810 3478 3866
rect 5956 3116 6012 3118
rect 6036 3116 6092 3118
rect 6116 3116 6172 3118
rect 6196 3116 6252 3118
rect 5956 3064 5982 3116
rect 5982 3064 6012 3116
rect 6036 3064 6046 3116
rect 6046 3064 6092 3116
rect 6116 3064 6162 3116
rect 6162 3064 6172 3116
rect 6196 3064 6226 3116
rect 6226 3064 6252 3116
rect 5956 3062 6012 3064
rect 6036 3062 6092 3064
rect 6116 3062 6172 3064
rect 6196 3062 6252 3064
rect 7838 10066 7894 10122
rect 8298 9930 8354 9986
rect 7378 2858 7434 2914
rect 2226 1498 2282 1554
rect 1674 1226 1730 1282
rect 1582 682 1638 738
rect 5956 2028 6012 2030
rect 6036 2028 6092 2030
rect 6116 2028 6172 2030
rect 6196 2028 6252 2030
rect 5956 1976 5982 2028
rect 5982 1976 6012 2028
rect 6036 1976 6046 2028
rect 6046 1976 6092 2028
rect 6116 1976 6162 2028
rect 6162 1976 6172 2028
rect 6196 1976 6226 2028
rect 6226 1976 6252 2028
rect 5956 1974 6012 1976
rect 6036 1974 6092 1976
rect 6116 1974 6172 1976
rect 6196 1974 6252 1976
rect 10956 10188 11012 10190
rect 11036 10188 11092 10190
rect 11116 10188 11172 10190
rect 11196 10188 11252 10190
rect 10956 10136 10982 10188
rect 10982 10136 11012 10188
rect 11036 10136 11046 10188
rect 11046 10136 11092 10188
rect 11116 10136 11162 10188
rect 11162 10136 11172 10188
rect 11196 10136 11226 10188
rect 11226 10136 11252 10188
rect 10956 10134 11012 10136
rect 11036 10134 11092 10136
rect 11116 10134 11172 10136
rect 11196 10134 11252 10136
rect 10956 9100 11012 9102
rect 11036 9100 11092 9102
rect 11116 9100 11172 9102
rect 11196 9100 11252 9102
rect 10956 9048 10982 9100
rect 10982 9048 11012 9100
rect 11036 9048 11046 9100
rect 11046 9048 11092 9100
rect 11116 9048 11162 9100
rect 11162 9048 11172 9100
rect 11196 9048 11226 9100
rect 11226 9048 11252 9100
rect 10956 9046 11012 9048
rect 11036 9046 11092 9048
rect 11116 9046 11172 9048
rect 11196 9046 11252 9048
rect 10782 8062 10784 8082
rect 10784 8062 10836 8082
rect 10836 8062 10838 8082
rect 10782 8026 10838 8062
rect 11334 8062 11336 8082
rect 11336 8062 11388 8082
rect 11388 8062 11390 8082
rect 11334 8026 11390 8062
rect 10956 8012 11012 8014
rect 11036 8012 11092 8014
rect 11116 8012 11172 8014
rect 11196 8012 11252 8014
rect 10956 7960 10982 8012
rect 10982 7960 11012 8012
rect 11036 7960 11046 8012
rect 11046 7960 11092 8012
rect 11116 7960 11162 8012
rect 11162 7960 11172 8012
rect 11196 7960 11226 8012
rect 11226 7960 11252 8012
rect 10956 7958 11012 7960
rect 11036 7958 11092 7960
rect 11116 7958 11172 7960
rect 11196 7958 11252 7960
rect 10874 7618 10930 7674
rect 10956 6924 11012 6926
rect 11036 6924 11092 6926
rect 11116 6924 11172 6926
rect 11196 6924 11252 6926
rect 10956 6872 10982 6924
rect 10982 6872 11012 6924
rect 11036 6872 11046 6924
rect 11046 6872 11092 6924
rect 11116 6872 11162 6924
rect 11162 6872 11172 6924
rect 11196 6872 11226 6924
rect 11226 6872 11252 6924
rect 10956 6870 11012 6872
rect 11036 6870 11092 6872
rect 11116 6870 11172 6872
rect 11196 6870 11252 6872
rect 11058 6122 11114 6178
rect 10956 5836 11012 5838
rect 11036 5836 11092 5838
rect 11116 5836 11172 5838
rect 11196 5836 11252 5838
rect 10956 5784 10982 5836
rect 10982 5784 11012 5836
rect 11036 5784 11046 5836
rect 11046 5784 11092 5836
rect 11116 5784 11162 5836
rect 11162 5784 11172 5836
rect 11196 5784 11226 5836
rect 11226 5784 11252 5836
rect 10956 5782 11012 5784
rect 11036 5782 11092 5784
rect 11116 5782 11172 5784
rect 11196 5782 11252 5784
rect 10956 4748 11012 4750
rect 11036 4748 11092 4750
rect 11116 4748 11172 4750
rect 11196 4748 11252 4750
rect 10956 4696 10982 4748
rect 10982 4696 11012 4748
rect 11036 4696 11046 4748
rect 11046 4696 11092 4748
rect 11116 4696 11162 4748
rect 11162 4696 11172 4748
rect 11196 4696 11226 4748
rect 11226 4696 11252 4748
rect 10956 4694 11012 4696
rect 11036 4694 11092 4696
rect 11116 4694 11172 4696
rect 11196 4694 11252 4696
rect 10956 3660 11012 3662
rect 11036 3660 11092 3662
rect 11116 3660 11172 3662
rect 11196 3660 11252 3662
rect 10956 3608 10982 3660
rect 10982 3608 11012 3660
rect 11036 3608 11046 3660
rect 11046 3608 11092 3660
rect 11116 3608 11162 3660
rect 11162 3608 11172 3660
rect 11196 3608 11226 3660
rect 11226 3608 11252 3660
rect 10956 3606 11012 3608
rect 11036 3606 11092 3608
rect 11116 3606 11172 3608
rect 11196 3606 11252 3608
rect 10956 2572 11012 2574
rect 11036 2572 11092 2574
rect 11116 2572 11172 2574
rect 11196 2572 11252 2574
rect 10956 2520 10982 2572
rect 10982 2520 11012 2572
rect 11036 2520 11046 2572
rect 11046 2520 11092 2572
rect 11116 2520 11162 2572
rect 11162 2520 11172 2572
rect 11196 2520 11226 2572
rect 11226 2520 11252 2572
rect 10956 2518 11012 2520
rect 11036 2518 11092 2520
rect 11116 2518 11172 2520
rect 11196 2518 11252 2520
rect 20956 19980 21012 19982
rect 21036 19980 21092 19982
rect 21116 19980 21172 19982
rect 21196 19980 21252 19982
rect 20956 19928 20982 19980
rect 20982 19928 21012 19980
rect 21036 19928 21046 19980
rect 21046 19928 21092 19980
rect 21116 19928 21162 19980
rect 21162 19928 21172 19980
rect 21196 19928 21226 19980
rect 21226 19928 21252 19980
rect 20956 19926 21012 19928
rect 21036 19926 21092 19928
rect 21116 19926 21172 19928
rect 21196 19926 21252 19928
rect 20626 19586 20682 19642
rect 23938 19078 23940 19098
rect 23940 19078 23992 19098
rect 23992 19078 23994 19098
rect 23938 19042 23994 19078
rect 20956 18892 21012 18894
rect 21036 18892 21092 18894
rect 21116 18892 21172 18894
rect 21196 18892 21252 18894
rect 20956 18840 20982 18892
rect 20982 18840 21012 18892
rect 21036 18840 21046 18892
rect 21046 18840 21092 18892
rect 21116 18840 21162 18892
rect 21162 18840 21172 18892
rect 21196 18840 21226 18892
rect 21226 18840 21252 18892
rect 20956 18838 21012 18840
rect 21036 18838 21092 18840
rect 21116 18838 21172 18840
rect 21196 18838 21252 18840
rect 23754 18126 23756 18146
rect 23756 18126 23808 18146
rect 23808 18126 23810 18146
rect 23754 18090 23810 18126
rect 23938 17990 23940 18010
rect 23940 17990 23992 18010
rect 23992 17990 23994 18010
rect 23938 17954 23994 17990
rect 20956 17804 21012 17806
rect 21036 17804 21092 17806
rect 21116 17804 21172 17806
rect 21196 17804 21252 17806
rect 20956 17752 20982 17804
rect 20982 17752 21012 17804
rect 21036 17752 21046 17804
rect 21046 17752 21092 17804
rect 21116 17752 21162 17804
rect 21162 17752 21172 17804
rect 21196 17752 21226 17804
rect 21226 17752 21252 17804
rect 20956 17750 21012 17752
rect 21036 17750 21092 17752
rect 21116 17750 21172 17752
rect 21196 17750 21252 17752
rect 20956 16716 21012 16718
rect 21036 16716 21092 16718
rect 21116 16716 21172 16718
rect 21196 16716 21252 16718
rect 20956 16664 20982 16716
rect 20982 16664 21012 16716
rect 21036 16664 21046 16716
rect 21046 16664 21092 16716
rect 21116 16664 21162 16716
rect 21162 16664 21172 16716
rect 21196 16664 21226 16716
rect 21226 16664 21252 16716
rect 20956 16662 21012 16664
rect 21036 16662 21092 16664
rect 21116 16662 21172 16664
rect 21196 16662 21252 16664
rect 20956 15628 21012 15630
rect 21036 15628 21092 15630
rect 21116 15628 21172 15630
rect 21196 15628 21252 15630
rect 20956 15576 20982 15628
rect 20982 15576 21012 15628
rect 21036 15576 21046 15628
rect 21046 15576 21092 15628
rect 21116 15576 21162 15628
rect 21162 15576 21172 15628
rect 21196 15576 21226 15628
rect 21226 15576 21252 15628
rect 20956 15574 21012 15576
rect 21036 15574 21092 15576
rect 21116 15574 21172 15576
rect 21196 15574 21252 15576
rect 20956 14540 21012 14542
rect 21036 14540 21092 14542
rect 21116 14540 21172 14542
rect 21196 14540 21252 14542
rect 20956 14488 20982 14540
rect 20982 14488 21012 14540
rect 21036 14488 21046 14540
rect 21046 14488 21092 14540
rect 21116 14488 21162 14540
rect 21162 14488 21172 14540
rect 21196 14488 21226 14540
rect 21226 14488 21252 14540
rect 20956 14486 21012 14488
rect 21036 14486 21092 14488
rect 21116 14486 21172 14488
rect 21196 14486 21252 14488
rect 23110 13602 23166 13658
rect 20956 13452 21012 13454
rect 21036 13452 21092 13454
rect 21116 13452 21172 13454
rect 21196 13452 21252 13454
rect 20956 13400 20982 13452
rect 20982 13400 21012 13452
rect 21036 13400 21046 13452
rect 21046 13400 21092 13452
rect 21116 13400 21162 13452
rect 21162 13400 21172 13452
rect 21196 13400 21226 13452
rect 21226 13400 21252 13452
rect 20956 13398 21012 13400
rect 21036 13398 21092 13400
rect 21116 13398 21172 13400
rect 21196 13398 21252 13400
rect 17222 11970 17278 12026
rect 15956 11820 16012 11822
rect 16036 11820 16092 11822
rect 16116 11820 16172 11822
rect 16196 11820 16252 11822
rect 15956 11768 15982 11820
rect 15982 11768 16012 11820
rect 16036 11768 16046 11820
rect 16046 11768 16092 11820
rect 16116 11768 16162 11820
rect 16162 11768 16172 11820
rect 16196 11768 16226 11820
rect 16226 11768 16252 11820
rect 15956 11766 16012 11768
rect 16036 11766 16092 11768
rect 16116 11766 16172 11768
rect 16196 11766 16252 11768
rect 17498 11562 17554 11618
rect 17222 11290 17278 11346
rect 17498 11018 17554 11074
rect 15956 10732 16012 10734
rect 16036 10732 16092 10734
rect 16116 10732 16172 10734
rect 16196 10732 16252 10734
rect 15956 10680 15982 10732
rect 15982 10680 16012 10732
rect 16036 10680 16046 10732
rect 16046 10680 16092 10732
rect 16116 10680 16162 10732
rect 16162 10680 16172 10732
rect 16196 10680 16226 10732
rect 16226 10680 16252 10732
rect 15956 10678 16012 10680
rect 16036 10678 16092 10680
rect 16116 10678 16172 10680
rect 16196 10678 16252 10680
rect 20956 12364 21012 12366
rect 21036 12364 21092 12366
rect 21116 12364 21172 12366
rect 21196 12364 21252 12366
rect 20956 12312 20982 12364
rect 20982 12312 21012 12364
rect 21036 12312 21046 12364
rect 21046 12312 21092 12364
rect 21116 12312 21162 12364
rect 21162 12312 21172 12364
rect 21196 12312 21226 12364
rect 21226 12312 21252 12364
rect 20956 12310 21012 12312
rect 21036 12310 21092 12312
rect 21116 12310 21172 12312
rect 21196 12310 21252 12312
rect 20442 12106 20498 12162
rect 20956 11276 21012 11278
rect 21036 11276 21092 11278
rect 21116 11276 21172 11278
rect 21196 11276 21252 11278
rect 20956 11224 20982 11276
rect 20982 11224 21012 11276
rect 21036 11224 21046 11276
rect 21046 11224 21092 11276
rect 21116 11224 21162 11276
rect 21162 11224 21172 11276
rect 21196 11224 21226 11276
rect 21226 11224 21252 11276
rect 20956 11222 21012 11224
rect 21036 11222 21092 11224
rect 21116 11222 21172 11224
rect 21196 11222 21252 11224
rect 20956 10188 21012 10190
rect 21036 10188 21092 10190
rect 21116 10188 21172 10190
rect 21196 10188 21252 10190
rect 20956 10136 20982 10188
rect 20982 10136 21012 10188
rect 21036 10136 21046 10188
rect 21046 10136 21092 10188
rect 21116 10136 21162 10188
rect 21162 10136 21172 10188
rect 21196 10136 21226 10188
rect 21226 10136 21252 10188
rect 20956 10134 21012 10136
rect 21036 10134 21092 10136
rect 21116 10134 21172 10136
rect 21196 10134 21252 10136
rect 19706 9794 19762 9850
rect 15956 9644 16012 9646
rect 16036 9644 16092 9646
rect 16116 9644 16172 9646
rect 16196 9644 16252 9646
rect 15956 9592 15982 9644
rect 15982 9592 16012 9644
rect 16036 9592 16046 9644
rect 16046 9592 16092 9644
rect 16116 9592 16162 9644
rect 16162 9592 16172 9644
rect 16196 9592 16226 9644
rect 16226 9592 16252 9644
rect 15956 9590 16012 9592
rect 16036 9590 16092 9592
rect 16116 9590 16172 9592
rect 16196 9590 16252 9592
rect 20956 9100 21012 9102
rect 21036 9100 21092 9102
rect 21116 9100 21172 9102
rect 21196 9100 21252 9102
rect 20956 9048 20982 9100
rect 20982 9048 21012 9100
rect 21036 9048 21046 9100
rect 21046 9048 21092 9100
rect 21116 9048 21162 9100
rect 21162 9048 21172 9100
rect 21196 9048 21226 9100
rect 21226 9048 21252 9100
rect 20956 9046 21012 9048
rect 21036 9046 21092 9048
rect 21116 9046 21172 9048
rect 21196 9046 21252 9048
rect 15956 8556 16012 8558
rect 16036 8556 16092 8558
rect 16116 8556 16172 8558
rect 16196 8556 16252 8558
rect 15956 8504 15982 8556
rect 15982 8504 16012 8556
rect 16036 8504 16046 8556
rect 16046 8504 16092 8556
rect 16116 8504 16162 8556
rect 16162 8504 16172 8556
rect 16196 8504 16226 8556
rect 16226 8504 16252 8556
rect 15956 8502 16012 8504
rect 16036 8502 16092 8504
rect 16116 8502 16172 8504
rect 16196 8502 16252 8504
rect 20956 8012 21012 8014
rect 21036 8012 21092 8014
rect 21116 8012 21172 8014
rect 21196 8012 21252 8014
rect 20956 7960 20982 8012
rect 20982 7960 21012 8012
rect 21036 7960 21046 8012
rect 21046 7960 21092 8012
rect 21116 7960 21162 8012
rect 21162 7960 21172 8012
rect 21196 7960 21226 8012
rect 21226 7960 21252 8012
rect 20956 7958 21012 7960
rect 21036 7958 21092 7960
rect 21116 7958 21172 7960
rect 21196 7958 21252 7960
rect 22650 7482 22706 7538
rect 15956 7468 16012 7470
rect 16036 7468 16092 7470
rect 16116 7468 16172 7470
rect 16196 7468 16252 7470
rect 15956 7416 15982 7468
rect 15982 7416 16012 7468
rect 16036 7416 16046 7468
rect 16046 7416 16092 7468
rect 16116 7416 16162 7468
rect 16162 7416 16172 7468
rect 16196 7416 16226 7468
rect 16226 7416 16252 7468
rect 15956 7414 16012 7416
rect 16036 7414 16092 7416
rect 16116 7414 16172 7416
rect 16196 7414 16252 7416
rect 23570 16866 23626 16922
rect 23478 13058 23534 13114
rect 23386 11834 23442 11890
rect 23478 7754 23534 7810
rect 18694 7210 18750 7266
rect 18878 7246 18880 7266
rect 18880 7246 18932 7266
rect 18932 7246 18934 7266
rect 18878 7210 18934 7246
rect 20956 6924 21012 6926
rect 21036 6924 21092 6926
rect 21116 6924 21172 6926
rect 21196 6924 21252 6926
rect 20956 6872 20982 6924
rect 20982 6872 21012 6924
rect 21036 6872 21046 6924
rect 21046 6872 21092 6924
rect 21116 6872 21162 6924
rect 21162 6872 21172 6924
rect 21196 6872 21226 6924
rect 21226 6872 21252 6924
rect 20956 6870 21012 6872
rect 21036 6870 21092 6872
rect 21116 6870 21172 6872
rect 21196 6870 21252 6872
rect 17222 6394 17278 6450
rect 15956 6380 16012 6382
rect 16036 6380 16092 6382
rect 16116 6380 16172 6382
rect 16196 6380 16252 6382
rect 15956 6328 15982 6380
rect 15982 6328 16012 6380
rect 16036 6328 16046 6380
rect 16046 6328 16092 6380
rect 16116 6328 16162 6380
rect 16162 6328 16172 6380
rect 16196 6328 16226 6380
rect 16226 6328 16252 6380
rect 15956 6326 16012 6328
rect 16036 6326 16092 6328
rect 16116 6326 16172 6328
rect 16196 6326 16252 6328
rect 14830 6122 14886 6178
rect 12806 5986 12862 6042
rect 17222 5986 17278 6042
rect 20956 5836 21012 5838
rect 21036 5836 21092 5838
rect 21116 5836 21172 5838
rect 21196 5836 21252 5838
rect 20956 5784 20982 5836
rect 20982 5784 21012 5836
rect 21036 5784 21046 5836
rect 21046 5784 21092 5836
rect 21116 5784 21162 5836
rect 21162 5784 21172 5836
rect 21196 5784 21226 5836
rect 21226 5784 21252 5836
rect 20956 5782 21012 5784
rect 21036 5782 21092 5784
rect 21116 5782 21172 5784
rect 21196 5782 21252 5784
rect 12622 5598 12678 5634
rect 12622 5578 12624 5598
rect 12624 5578 12676 5598
rect 12676 5578 12678 5598
rect 15956 5292 16012 5294
rect 16036 5292 16092 5294
rect 16116 5292 16172 5294
rect 16196 5292 16252 5294
rect 15956 5240 15982 5292
rect 15982 5240 16012 5292
rect 16036 5240 16046 5292
rect 16046 5240 16092 5292
rect 16116 5240 16162 5292
rect 16162 5240 16172 5292
rect 16196 5240 16226 5292
rect 16226 5240 16252 5292
rect 15956 5238 16012 5240
rect 16036 5238 16092 5240
rect 16116 5238 16172 5240
rect 16196 5238 16252 5240
rect 16394 5190 16450 5226
rect 16394 5170 16396 5190
rect 16396 5170 16448 5190
rect 16448 5170 16450 5190
rect 13726 5034 13782 5090
rect 23938 15234 23994 15290
rect 23662 9386 23718 9442
rect 24398 22170 24454 22226
rect 24122 11426 24178 11482
rect 24858 21354 24914 21410
rect 24490 21082 24546 21138
rect 24858 20266 24914 20322
rect 24582 17682 24638 17738
rect 24490 12242 24546 12298
rect 23938 9286 23940 9306
rect 23940 9286 23992 9306
rect 23992 9286 23994 9306
rect 23938 9250 23994 9286
rect 23754 8842 23810 8898
rect 23938 7110 23940 7130
rect 23940 7110 23992 7130
rect 23992 7110 23994 7130
rect 23938 7074 23994 7110
rect 20956 4748 21012 4750
rect 21036 4748 21092 4750
rect 21116 4748 21172 4750
rect 21196 4748 21252 4750
rect 20956 4696 20982 4748
rect 20982 4696 21012 4748
rect 21036 4696 21046 4748
rect 21046 4696 21092 4748
rect 21116 4696 21162 4748
rect 21162 4696 21172 4748
rect 21196 4696 21226 4748
rect 21226 4696 21252 4748
rect 20956 4694 21012 4696
rect 21036 4694 21092 4696
rect 21116 4694 21172 4696
rect 21196 4694 21252 4696
rect 20718 4510 20774 4546
rect 20718 4490 20720 4510
rect 20720 4490 20772 4510
rect 20772 4490 20774 4510
rect 15956 4204 16012 4206
rect 16036 4204 16092 4206
rect 16116 4204 16172 4206
rect 16196 4204 16252 4206
rect 15956 4152 15982 4204
rect 15982 4152 16012 4204
rect 16036 4152 16046 4204
rect 16046 4152 16092 4204
rect 16116 4152 16162 4204
rect 16162 4152 16172 4204
rect 16196 4152 16226 4204
rect 16226 4152 16252 4204
rect 15956 4150 16012 4152
rect 16036 4150 16092 4152
rect 16116 4150 16172 4152
rect 16196 4150 16252 4152
rect 16486 4374 16542 4410
rect 16486 4354 16488 4374
rect 16488 4354 16540 4374
rect 16540 4354 16542 4374
rect 20902 4374 20958 4410
rect 20902 4354 20904 4374
rect 20904 4354 20956 4374
rect 20956 4354 20958 4374
rect 16394 3982 16396 4002
rect 16396 3982 16448 4002
rect 16448 3982 16450 4002
rect 16394 3946 16450 3982
rect 23938 3846 23940 3866
rect 23940 3846 23992 3866
rect 23992 3846 23994 3866
rect 23938 3810 23994 3846
rect 20956 3660 21012 3662
rect 21036 3660 21092 3662
rect 21116 3660 21172 3662
rect 21196 3660 21252 3662
rect 20956 3608 20982 3660
rect 20982 3608 21012 3660
rect 21036 3608 21046 3660
rect 21046 3608 21092 3660
rect 21116 3608 21162 3660
rect 21162 3608 21172 3660
rect 21196 3608 21226 3660
rect 21226 3608 21252 3660
rect 20956 3606 21012 3608
rect 21036 3606 21092 3608
rect 21116 3606 21172 3608
rect 21196 3606 21252 3608
rect 22098 3538 22154 3594
rect 21638 3402 21694 3458
rect 24122 10474 24178 10530
rect 24122 9150 24124 9170
rect 24124 9150 24176 9170
rect 24176 9150 24178 9170
rect 24122 9114 24178 9150
rect 24122 8298 24178 8354
rect 24122 7910 24178 7946
rect 24122 7890 24124 7910
rect 24124 7890 24176 7910
rect 24176 7890 24178 7910
rect 24950 19858 25006 19914
rect 25956 21612 26012 21614
rect 26036 21612 26092 21614
rect 26116 21612 26172 21614
rect 26196 21612 26252 21614
rect 25956 21560 25982 21612
rect 25982 21560 26012 21612
rect 26036 21560 26046 21612
rect 26046 21560 26092 21612
rect 26116 21560 26162 21612
rect 26162 21560 26172 21612
rect 26196 21560 26226 21612
rect 26226 21560 26252 21612
rect 25956 21558 26012 21560
rect 26036 21558 26092 21560
rect 26116 21558 26172 21560
rect 26196 21558 26252 21560
rect 25956 20524 26012 20526
rect 26036 20524 26092 20526
rect 26116 20524 26172 20526
rect 26196 20524 26252 20526
rect 25956 20472 25982 20524
rect 25982 20472 26012 20524
rect 26036 20472 26046 20524
rect 26046 20472 26092 20524
rect 26116 20472 26162 20524
rect 26162 20472 26172 20524
rect 26196 20472 26226 20524
rect 26226 20472 26252 20524
rect 25956 20470 26012 20472
rect 26036 20470 26092 20472
rect 26116 20470 26172 20472
rect 26196 20470 26252 20472
rect 25870 19586 25926 19642
rect 25956 19436 26012 19438
rect 26036 19436 26092 19438
rect 26116 19436 26172 19438
rect 26196 19436 26252 19438
rect 25956 19384 25982 19436
rect 25982 19384 26012 19436
rect 26036 19384 26046 19436
rect 26046 19384 26092 19436
rect 26116 19384 26162 19436
rect 26162 19384 26172 19436
rect 26196 19384 26226 19436
rect 26226 19384 26252 19436
rect 25956 19382 26012 19384
rect 26036 19382 26092 19384
rect 26116 19382 26172 19384
rect 26196 19382 26252 19384
rect 25594 19178 25650 19234
rect 25226 18634 25282 18690
rect 24950 17682 25006 17738
rect 24674 11834 24730 11890
rect 25134 13194 25190 13250
rect 24950 12106 25006 12162
rect 24858 11970 24914 12026
rect 24766 10882 24822 10938
rect 25042 11834 25098 11890
rect 24950 10338 25006 10394
rect 25502 15642 25558 15698
rect 25410 14418 25466 14474
rect 25318 13738 25374 13794
rect 25226 12242 25282 12298
rect 25410 11698 25466 11754
rect 25318 11562 25374 11618
rect 25134 11018 25190 11074
rect 25042 10202 25098 10258
rect 24858 9794 24914 9850
rect 24490 8198 24492 8218
rect 24492 8198 24544 8218
rect 24544 8198 24546 8218
rect 24490 8162 24546 8198
rect 24122 6550 24178 6586
rect 24122 6530 24124 6550
rect 24124 6530 24176 6550
rect 24176 6530 24178 6550
rect 24122 4898 24178 4954
rect 24122 3710 24124 3730
rect 24124 3710 24176 3730
rect 24176 3710 24178 3730
rect 24122 3674 24178 3710
rect 25956 18348 26012 18350
rect 26036 18348 26092 18350
rect 26116 18348 26172 18350
rect 26196 18348 26252 18350
rect 25956 18296 25982 18348
rect 25982 18296 26012 18348
rect 26036 18296 26046 18348
rect 26046 18296 26092 18348
rect 26116 18296 26162 18348
rect 26162 18296 26172 18348
rect 26196 18296 26226 18348
rect 26226 18296 26252 18348
rect 25956 18294 26012 18296
rect 26036 18294 26092 18296
rect 26116 18294 26172 18296
rect 26196 18294 26252 18296
rect 25778 17410 25834 17466
rect 25686 15914 25742 15970
rect 25594 13602 25650 13658
rect 25594 12650 25650 12706
rect 25502 3538 25558 3594
rect 15956 3116 16012 3118
rect 16036 3116 16092 3118
rect 16116 3116 16172 3118
rect 16196 3116 16252 3118
rect 15956 3064 15982 3116
rect 15982 3064 16012 3116
rect 16036 3064 16046 3116
rect 16046 3064 16092 3116
rect 16116 3064 16162 3116
rect 16162 3064 16172 3116
rect 16196 3064 16226 3116
rect 16226 3064 16252 3116
rect 15956 3062 16012 3064
rect 16036 3062 16092 3064
rect 16116 3062 16172 3064
rect 16196 3062 16252 3064
rect 24122 3286 24178 3322
rect 24122 3266 24124 3286
rect 24124 3266 24176 3286
rect 24176 3266 24178 3286
rect 23938 2858 23994 2914
rect 20956 2572 21012 2574
rect 21036 2572 21092 2574
rect 21116 2572 21172 2574
rect 21196 2572 21252 2574
rect 20956 2520 20982 2572
rect 20982 2520 21012 2572
rect 21036 2520 21046 2572
rect 21046 2520 21092 2572
rect 21116 2520 21162 2572
rect 21162 2520 21172 2572
rect 21196 2520 21226 2572
rect 21226 2520 21252 2572
rect 20956 2518 21012 2520
rect 21036 2518 21092 2520
rect 21116 2518 21172 2520
rect 21196 2518 21252 2520
rect 24214 2470 24270 2506
rect 24214 2450 24216 2470
rect 24216 2450 24268 2470
rect 24268 2450 24270 2470
rect 12530 2178 12586 2234
rect 24030 2178 24086 2234
rect 15956 2028 16012 2030
rect 16036 2028 16092 2030
rect 16116 2028 16172 2030
rect 16196 2028 16252 2030
rect 15956 1976 15982 2028
rect 15982 1976 16012 2028
rect 16036 1976 16046 2028
rect 16046 1976 16092 2028
rect 16116 1976 16162 2028
rect 16162 1976 16172 2028
rect 16196 1976 16226 2028
rect 16226 1976 16252 2028
rect 15956 1974 16012 1976
rect 16036 1974 16092 1976
rect 16116 1974 16172 1976
rect 16196 1974 16252 1976
rect 8390 1770 8446 1826
rect 25956 17260 26012 17262
rect 26036 17260 26092 17262
rect 26116 17260 26172 17262
rect 26196 17260 26252 17262
rect 25956 17208 25982 17260
rect 25982 17208 26012 17260
rect 26036 17208 26046 17260
rect 26046 17208 26092 17260
rect 26116 17208 26162 17260
rect 26162 17208 26172 17260
rect 26196 17208 26226 17260
rect 26226 17208 26252 17260
rect 25956 17206 26012 17208
rect 26036 17206 26092 17208
rect 26116 17206 26172 17208
rect 26196 17206 26252 17208
rect 25956 16172 26012 16174
rect 26036 16172 26092 16174
rect 26116 16172 26172 16174
rect 26196 16172 26252 16174
rect 25956 16120 25982 16172
rect 25982 16120 26012 16172
rect 26036 16120 26046 16172
rect 26046 16120 26092 16172
rect 26116 16120 26162 16172
rect 26162 16120 26172 16172
rect 26196 16120 26226 16172
rect 26226 16120 26252 16172
rect 25956 16118 26012 16120
rect 26036 16118 26092 16120
rect 26116 16118 26172 16120
rect 26196 16118 26252 16120
rect 25956 15084 26012 15086
rect 26036 15084 26092 15086
rect 26116 15084 26172 15086
rect 26196 15084 26252 15086
rect 25956 15032 25982 15084
rect 25982 15032 26012 15084
rect 26036 15032 26046 15084
rect 26046 15032 26092 15084
rect 26116 15032 26162 15084
rect 26162 15032 26172 15084
rect 26196 15032 26226 15084
rect 26226 15032 26252 15084
rect 25956 15030 26012 15032
rect 26036 15030 26092 15032
rect 26116 15030 26172 15032
rect 26196 15030 26252 15032
rect 25956 13996 26012 13998
rect 26036 13996 26092 13998
rect 26116 13996 26172 13998
rect 26196 13996 26252 13998
rect 25956 13944 25982 13996
rect 25982 13944 26012 13996
rect 26036 13944 26046 13996
rect 26046 13944 26092 13996
rect 26116 13944 26162 13996
rect 26162 13944 26172 13996
rect 26196 13944 26226 13996
rect 26226 13944 26252 13996
rect 25956 13942 26012 13944
rect 26036 13942 26092 13944
rect 26116 13942 26172 13944
rect 26196 13942 26252 13944
rect 25956 12908 26012 12910
rect 26036 12908 26092 12910
rect 26116 12908 26172 12910
rect 26196 12908 26252 12910
rect 25956 12856 25982 12908
rect 25982 12856 26012 12908
rect 26036 12856 26046 12908
rect 26046 12856 26092 12908
rect 26116 12856 26162 12908
rect 26162 12856 26172 12908
rect 26196 12856 26226 12908
rect 26226 12856 26252 12908
rect 25956 12854 26012 12856
rect 26036 12854 26092 12856
rect 26116 12854 26172 12856
rect 26196 12854 26252 12856
rect 25956 11820 26012 11822
rect 26036 11820 26092 11822
rect 26116 11820 26172 11822
rect 26196 11820 26252 11822
rect 25956 11768 25982 11820
rect 25982 11768 26012 11820
rect 26036 11768 26046 11820
rect 26046 11768 26092 11820
rect 26116 11768 26162 11820
rect 26162 11768 26172 11820
rect 26196 11768 26226 11820
rect 26226 11768 26252 11820
rect 25956 11766 26012 11768
rect 26036 11766 26092 11768
rect 26116 11766 26172 11768
rect 26196 11766 26252 11768
rect 25956 10732 26012 10734
rect 26036 10732 26092 10734
rect 26116 10732 26172 10734
rect 26196 10732 26252 10734
rect 25956 10680 25982 10732
rect 25982 10680 26012 10732
rect 26036 10680 26046 10732
rect 26046 10680 26092 10732
rect 26116 10680 26162 10732
rect 26162 10680 26172 10732
rect 26196 10680 26226 10732
rect 26226 10680 26252 10732
rect 25956 10678 26012 10680
rect 26036 10678 26092 10680
rect 26116 10678 26172 10680
rect 26196 10678 26252 10680
rect 25956 9644 26012 9646
rect 26036 9644 26092 9646
rect 26116 9644 26172 9646
rect 26196 9644 26252 9646
rect 25956 9592 25982 9644
rect 25982 9592 26012 9644
rect 26036 9592 26046 9644
rect 26046 9592 26092 9644
rect 26116 9592 26162 9644
rect 26162 9592 26172 9644
rect 26196 9592 26226 9644
rect 26226 9592 26252 9644
rect 25956 9590 26012 9592
rect 26036 9590 26092 9592
rect 26116 9590 26172 9592
rect 26196 9590 26252 9592
rect 25956 8556 26012 8558
rect 26036 8556 26092 8558
rect 26116 8556 26172 8558
rect 26196 8556 26252 8558
rect 25956 8504 25982 8556
rect 25982 8504 26012 8556
rect 26036 8504 26046 8556
rect 26046 8504 26092 8556
rect 26116 8504 26162 8556
rect 26162 8504 26172 8556
rect 26196 8504 26226 8556
rect 26226 8504 26252 8556
rect 25956 8502 26012 8504
rect 26036 8502 26092 8504
rect 26116 8502 26172 8504
rect 26196 8502 26252 8504
rect 25956 7468 26012 7470
rect 26036 7468 26092 7470
rect 26116 7468 26172 7470
rect 26196 7468 26252 7470
rect 25956 7416 25982 7468
rect 25982 7416 26012 7468
rect 26036 7416 26046 7468
rect 26046 7416 26092 7468
rect 26116 7416 26162 7468
rect 26162 7416 26172 7468
rect 26196 7416 26226 7468
rect 26226 7416 26252 7468
rect 25956 7414 26012 7416
rect 26036 7414 26092 7416
rect 26116 7414 26172 7416
rect 26196 7414 26252 7416
rect 25956 6380 26012 6382
rect 26036 6380 26092 6382
rect 26116 6380 26172 6382
rect 26196 6380 26252 6382
rect 25956 6328 25982 6380
rect 25982 6328 26012 6380
rect 26036 6328 26046 6380
rect 26046 6328 26092 6380
rect 26116 6328 26162 6380
rect 26162 6328 26172 6380
rect 26196 6328 26226 6380
rect 26226 6328 26252 6380
rect 25956 6326 26012 6328
rect 26036 6326 26092 6328
rect 26116 6326 26172 6328
rect 26196 6326 26252 6328
rect 25778 5578 25834 5634
rect 25956 5292 26012 5294
rect 26036 5292 26092 5294
rect 26116 5292 26172 5294
rect 26196 5292 26252 5294
rect 25956 5240 25982 5292
rect 25982 5240 26012 5292
rect 26036 5240 26046 5292
rect 26046 5240 26092 5292
rect 26116 5240 26162 5292
rect 26162 5240 26172 5292
rect 26196 5240 26226 5292
rect 26226 5240 26252 5292
rect 25956 5238 26012 5240
rect 26036 5238 26092 5240
rect 26116 5238 26172 5240
rect 26196 5238 26252 5240
rect 25956 4204 26012 4206
rect 26036 4204 26092 4206
rect 26116 4204 26172 4206
rect 26196 4204 26252 4206
rect 25956 4152 25982 4204
rect 25982 4152 26012 4204
rect 26036 4152 26046 4204
rect 26046 4152 26092 4204
rect 26116 4152 26162 4204
rect 26162 4152 26172 4204
rect 26196 4152 26226 4204
rect 26226 4152 26252 4204
rect 25956 4150 26012 4152
rect 26036 4150 26092 4152
rect 26116 4150 26172 4152
rect 26196 4150 26252 4152
rect 25686 3946 25742 4002
rect 25956 3116 26012 3118
rect 26036 3116 26092 3118
rect 26116 3116 26172 3118
rect 26196 3116 26252 3118
rect 25956 3064 25982 3116
rect 25982 3064 26012 3116
rect 26036 3064 26046 3116
rect 26046 3064 26092 3116
rect 26116 3064 26162 3116
rect 26162 3064 26172 3116
rect 26196 3064 26226 3116
rect 26226 3064 26252 3116
rect 25956 3062 26012 3064
rect 26036 3062 26092 3064
rect 26116 3062 26172 3064
rect 26196 3062 26252 3064
rect 25594 2314 25650 2370
rect 25134 1770 25190 1826
rect 24858 1362 24914 1418
rect 25956 2028 26012 2030
rect 26036 2028 26092 2030
rect 26116 2028 26172 2030
rect 26196 2028 26252 2030
rect 25956 1976 25982 2028
rect 25982 1976 26012 2028
rect 26036 1976 26046 2028
rect 26046 1976 26092 2028
rect 26116 1976 26162 2028
rect 26162 1976 26172 2028
rect 26196 1976 26226 2028
rect 26226 1976 26252 2028
rect 25956 1974 26012 1976
rect 26036 1974 26092 1976
rect 26116 1974 26172 1976
rect 26196 1974 26252 1976
rect 1490 138 1546 194
rect 2686 138 2742 194
rect 25318 138 25374 194
<< metal3 >>
rect 0 23452 480 23482
rect 3877 23452 3943 23455
rect 0 23450 3943 23452
rect 0 23394 3882 23450
rect 3938 23394 3943 23450
rect 0 23392 3943 23394
rect 0 23362 480 23392
rect 3877 23389 3943 23392
rect 25037 23452 25103 23455
rect 29520 23452 30000 23482
rect 25037 23450 30000 23452
rect 25037 23394 25042 23450
rect 25098 23394 30000 23450
rect 25037 23392 30000 23394
rect 25037 23389 25103 23392
rect 29520 23362 30000 23392
rect 0 22908 480 22938
rect 3049 22908 3115 22911
rect 0 22906 3115 22908
rect 0 22850 3054 22906
rect 3110 22850 3115 22906
rect 0 22848 3115 22850
rect 0 22818 480 22848
rect 3049 22845 3115 22848
rect 24301 22908 24367 22911
rect 29520 22908 30000 22938
rect 24301 22906 30000 22908
rect 24301 22850 24306 22906
rect 24362 22850 30000 22906
rect 24301 22848 30000 22850
rect 24301 22845 24367 22848
rect 29520 22818 30000 22848
rect 0 22228 480 22258
rect 3325 22228 3391 22231
rect 0 22226 3391 22228
rect 0 22170 3330 22226
rect 3386 22170 3391 22226
rect 0 22168 3391 22170
rect 0 22138 480 22168
rect 3325 22165 3391 22168
rect 24393 22228 24459 22231
rect 29520 22228 30000 22258
rect 24393 22226 30000 22228
rect 24393 22170 24398 22226
rect 24454 22170 30000 22226
rect 24393 22168 30000 22170
rect 24393 22165 24459 22168
rect 29520 22138 30000 22168
rect 0 21684 480 21714
rect 3417 21684 3483 21687
rect 29520 21684 30000 21714
rect 0 21682 3483 21684
rect 0 21626 3422 21682
rect 3478 21626 3483 21682
rect 0 21624 3483 21626
rect 0 21594 480 21624
rect 3417 21621 3483 21624
rect 27846 21624 30000 21684
rect 5944 21618 6264 21619
rect 5944 21554 5952 21618
rect 6016 21554 6032 21618
rect 6096 21554 6112 21618
rect 6176 21554 6192 21618
rect 6256 21554 6264 21618
rect 5944 21553 6264 21554
rect 15944 21618 16264 21619
rect 15944 21554 15952 21618
rect 16016 21554 16032 21618
rect 16096 21554 16112 21618
rect 16176 21554 16192 21618
rect 16256 21554 16264 21618
rect 15944 21553 16264 21554
rect 25944 21618 26264 21619
rect 25944 21554 25952 21618
rect 26016 21554 26032 21618
rect 26096 21554 26112 21618
rect 26176 21554 26192 21618
rect 26256 21554 26264 21618
rect 25944 21553 26264 21554
rect 24853 21412 24919 21415
rect 27846 21412 27906 21624
rect 29520 21594 30000 21624
rect 24853 21410 27906 21412
rect 24853 21354 24858 21410
rect 24914 21354 27906 21410
rect 24853 21352 27906 21354
rect 24853 21349 24919 21352
rect 0 21140 480 21170
rect 3509 21140 3575 21143
rect 0 21138 3575 21140
rect 0 21082 3514 21138
rect 3570 21082 3575 21138
rect 0 21080 3575 21082
rect 0 21050 480 21080
rect 3509 21077 3575 21080
rect 24485 21140 24551 21143
rect 29520 21140 30000 21170
rect 24485 21138 30000 21140
rect 24485 21082 24490 21138
rect 24546 21082 30000 21138
rect 24485 21080 30000 21082
rect 24485 21077 24551 21080
rect 10944 21074 11264 21075
rect 10944 21010 10952 21074
rect 11016 21010 11032 21074
rect 11096 21010 11112 21074
rect 11176 21010 11192 21074
rect 11256 21010 11264 21074
rect 10944 21009 11264 21010
rect 20944 21074 21264 21075
rect 20944 21010 20952 21074
rect 21016 21010 21032 21074
rect 21096 21010 21112 21074
rect 21176 21010 21192 21074
rect 21256 21010 21264 21074
rect 29520 21050 30000 21080
rect 20944 21009 21264 21010
rect 5944 20530 6264 20531
rect 0 20460 480 20490
rect 5944 20466 5952 20530
rect 6016 20466 6032 20530
rect 6096 20466 6112 20530
rect 6176 20466 6192 20530
rect 6256 20466 6264 20530
rect 5944 20465 6264 20466
rect 15944 20530 16264 20531
rect 15944 20466 15952 20530
rect 16016 20466 16032 20530
rect 16096 20466 16112 20530
rect 16176 20466 16192 20530
rect 16256 20466 16264 20530
rect 15944 20465 16264 20466
rect 25944 20530 26264 20531
rect 25944 20466 25952 20530
rect 26016 20466 26032 20530
rect 26096 20466 26112 20530
rect 26176 20466 26192 20530
rect 26256 20466 26264 20530
rect 25944 20465 26264 20466
rect 3969 20460 4035 20463
rect 29520 20460 30000 20490
rect 0 20458 4035 20460
rect 0 20402 3974 20458
rect 4030 20402 4035 20458
rect 0 20400 4035 20402
rect 0 20370 480 20400
rect 3969 20397 4035 20400
rect 27846 20400 30000 20460
rect 24853 20324 24919 20327
rect 27846 20324 27906 20400
rect 29520 20370 30000 20400
rect 24853 20322 27906 20324
rect 24853 20266 24858 20322
rect 24914 20266 27906 20322
rect 24853 20264 27906 20266
rect 24853 20261 24919 20264
rect 10944 19986 11264 19987
rect 0 19916 480 19946
rect 10944 19922 10952 19986
rect 11016 19922 11032 19986
rect 11096 19922 11112 19986
rect 11176 19922 11192 19986
rect 11256 19922 11264 19986
rect 10944 19921 11264 19922
rect 20944 19986 21264 19987
rect 20944 19922 20952 19986
rect 21016 19922 21032 19986
rect 21096 19922 21112 19986
rect 21176 19922 21192 19986
rect 21256 19922 21264 19986
rect 20944 19921 21264 19922
rect 3785 19916 3851 19919
rect 0 19914 3851 19916
rect 0 19858 3790 19914
rect 3846 19858 3851 19914
rect 0 19856 3851 19858
rect 0 19826 480 19856
rect 3785 19853 3851 19856
rect 24945 19916 25011 19919
rect 29520 19916 30000 19946
rect 24945 19914 30000 19916
rect 24945 19858 24950 19914
rect 25006 19858 30000 19914
rect 24945 19856 30000 19858
rect 24945 19853 25011 19856
rect 29520 19826 30000 19856
rect 20621 19644 20687 19647
rect 25865 19644 25931 19647
rect 20621 19642 25931 19644
rect 20621 19586 20626 19642
rect 20682 19586 25870 19642
rect 25926 19586 25931 19642
rect 20621 19584 25931 19586
rect 20621 19581 20687 19584
rect 25865 19581 25931 19584
rect 5944 19442 6264 19443
rect 5944 19378 5952 19442
rect 6016 19378 6032 19442
rect 6096 19378 6112 19442
rect 6176 19378 6192 19442
rect 6256 19378 6264 19442
rect 5944 19377 6264 19378
rect 15944 19442 16264 19443
rect 15944 19378 15952 19442
rect 16016 19378 16032 19442
rect 16096 19378 16112 19442
rect 16176 19378 16192 19442
rect 16256 19378 16264 19442
rect 15944 19377 16264 19378
rect 25944 19442 26264 19443
rect 25944 19378 25952 19442
rect 26016 19378 26032 19442
rect 26096 19378 26112 19442
rect 26176 19378 26192 19442
rect 26256 19378 26264 19442
rect 25944 19377 26264 19378
rect 0 19236 480 19266
rect 3417 19236 3483 19239
rect 0 19234 3483 19236
rect 0 19178 3422 19234
rect 3478 19178 3483 19234
rect 0 19176 3483 19178
rect 0 19146 480 19176
rect 3417 19173 3483 19176
rect 8845 19236 8911 19239
rect 11329 19236 11395 19239
rect 8845 19234 11395 19236
rect 8845 19178 8850 19234
rect 8906 19178 11334 19234
rect 11390 19178 11395 19234
rect 8845 19176 11395 19178
rect 8845 19173 8911 19176
rect 11329 19173 11395 19176
rect 25589 19236 25655 19239
rect 29520 19236 30000 19266
rect 25589 19234 30000 19236
rect 25589 19178 25594 19234
rect 25650 19178 30000 19234
rect 25589 19176 30000 19178
rect 25589 19173 25655 19176
rect 29520 19146 30000 19176
rect 3325 19100 3391 19103
rect 23933 19100 23999 19103
rect 3325 19098 23999 19100
rect 3325 19042 3330 19098
rect 3386 19042 23938 19098
rect 23994 19042 23999 19098
rect 3325 19040 23999 19042
rect 3325 19037 3391 19040
rect 23933 19037 23999 19040
rect 10944 18898 11264 18899
rect 10944 18834 10952 18898
rect 11016 18834 11032 18898
rect 11096 18834 11112 18898
rect 11176 18834 11192 18898
rect 11256 18834 11264 18898
rect 10944 18833 11264 18834
rect 20944 18898 21264 18899
rect 20944 18834 20952 18898
rect 21016 18834 21032 18898
rect 21096 18834 21112 18898
rect 21176 18834 21192 18898
rect 21256 18834 21264 18898
rect 20944 18833 21264 18834
rect 16665 18828 16731 18831
rect 18689 18828 18755 18831
rect 16665 18826 18755 18828
rect 16665 18770 16670 18826
rect 16726 18770 18694 18826
rect 18750 18770 18755 18826
rect 16665 18768 18755 18770
rect 16665 18765 16731 18768
rect 18689 18765 18755 18768
rect 0 18692 480 18722
rect 3141 18692 3207 18695
rect 0 18690 3207 18692
rect 0 18634 3146 18690
rect 3202 18634 3207 18690
rect 0 18632 3207 18634
rect 0 18602 480 18632
rect 3141 18629 3207 18632
rect 3693 18692 3759 18695
rect 7005 18692 7071 18695
rect 8569 18692 8635 18695
rect 12985 18692 13051 18695
rect 15285 18692 15351 18695
rect 3693 18690 15351 18692
rect 3693 18634 3698 18690
rect 3754 18634 7010 18690
rect 7066 18634 8574 18690
rect 8630 18634 12990 18690
rect 13046 18634 15290 18690
rect 15346 18634 15351 18690
rect 3693 18632 15351 18634
rect 3693 18629 3759 18632
rect 7005 18629 7071 18632
rect 8569 18629 8635 18632
rect 12985 18629 13051 18632
rect 15285 18629 15351 18632
rect 25221 18692 25287 18695
rect 29520 18692 30000 18722
rect 25221 18690 30000 18692
rect 25221 18634 25226 18690
rect 25282 18634 30000 18690
rect 25221 18632 30000 18634
rect 25221 18629 25287 18632
rect 29520 18602 30000 18632
rect 5944 18354 6264 18355
rect 5944 18290 5952 18354
rect 6016 18290 6032 18354
rect 6096 18290 6112 18354
rect 6176 18290 6192 18354
rect 6256 18290 6264 18354
rect 5944 18289 6264 18290
rect 15944 18354 16264 18355
rect 15944 18290 15952 18354
rect 16016 18290 16032 18354
rect 16096 18290 16112 18354
rect 16176 18290 16192 18354
rect 16256 18290 16264 18354
rect 15944 18289 16264 18290
rect 25944 18354 26264 18355
rect 25944 18290 25952 18354
rect 26016 18290 26032 18354
rect 26096 18290 26112 18354
rect 26176 18290 26192 18354
rect 26256 18290 26264 18354
rect 25944 18289 26264 18290
rect 19885 18284 19951 18287
rect 19885 18282 24042 18284
rect 19885 18226 19890 18282
rect 19946 18226 24042 18282
rect 19885 18224 24042 18226
rect 19885 18221 19951 18224
rect 0 18148 480 18178
rect 3233 18148 3299 18151
rect 0 18146 3299 18148
rect 0 18090 3238 18146
rect 3294 18090 3299 18146
rect 0 18088 3299 18090
rect 0 18058 480 18088
rect 3233 18085 3299 18088
rect 3877 18148 3943 18151
rect 23749 18148 23815 18151
rect 3877 18146 23815 18148
rect 3877 18090 3882 18146
rect 3938 18090 23754 18146
rect 23810 18090 23815 18146
rect 3877 18088 23815 18090
rect 23982 18148 24042 18224
rect 29520 18148 30000 18178
rect 23982 18088 30000 18148
rect 3877 18085 3943 18088
rect 23749 18085 23815 18088
rect 29520 18058 30000 18088
rect 3049 18012 3115 18015
rect 23933 18012 23999 18015
rect 3049 18010 23999 18012
rect 3049 17954 3054 18010
rect 3110 17954 23938 18010
rect 23994 17954 23999 18010
rect 3049 17952 23999 17954
rect 3049 17949 3115 17952
rect 23933 17949 23999 17952
rect 10944 17810 11264 17811
rect 10944 17746 10952 17810
rect 11016 17746 11032 17810
rect 11096 17746 11112 17810
rect 11176 17746 11192 17810
rect 11256 17746 11264 17810
rect 10944 17745 11264 17746
rect 20944 17810 21264 17811
rect 20944 17746 20952 17810
rect 21016 17746 21032 17810
rect 21096 17746 21112 17810
rect 21176 17746 21192 17810
rect 21256 17746 21264 17810
rect 20944 17745 21264 17746
rect 24577 17740 24643 17743
rect 24945 17740 25011 17743
rect 24577 17738 25011 17740
rect 24577 17682 24582 17738
rect 24638 17682 24950 17738
rect 25006 17682 25011 17738
rect 24577 17680 25011 17682
rect 24577 17677 24643 17680
rect 24945 17677 25011 17680
rect 0 17468 480 17498
rect 3325 17468 3391 17471
rect 0 17466 3391 17468
rect 0 17410 3330 17466
rect 3386 17410 3391 17466
rect 0 17408 3391 17410
rect 0 17378 480 17408
rect 3325 17405 3391 17408
rect 25773 17468 25839 17471
rect 29520 17468 30000 17498
rect 25773 17466 30000 17468
rect 25773 17410 25778 17466
rect 25834 17410 30000 17466
rect 25773 17408 30000 17410
rect 25773 17405 25839 17408
rect 29520 17378 30000 17408
rect 5944 17266 6264 17267
rect 5944 17202 5952 17266
rect 6016 17202 6032 17266
rect 6096 17202 6112 17266
rect 6176 17202 6192 17266
rect 6256 17202 6264 17266
rect 5944 17201 6264 17202
rect 15944 17266 16264 17267
rect 15944 17202 15952 17266
rect 16016 17202 16032 17266
rect 16096 17202 16112 17266
rect 16176 17202 16192 17266
rect 16256 17202 16264 17266
rect 15944 17201 16264 17202
rect 25944 17266 26264 17267
rect 25944 17202 25952 17266
rect 26016 17202 26032 17266
rect 26096 17202 26112 17266
rect 26176 17202 26192 17266
rect 26256 17202 26264 17266
rect 25944 17201 26264 17202
rect 0 16924 480 16954
rect 3509 16924 3575 16927
rect 0 16922 3575 16924
rect 0 16866 3514 16922
rect 3570 16866 3575 16922
rect 0 16864 3575 16866
rect 0 16834 480 16864
rect 3509 16861 3575 16864
rect 23565 16924 23631 16927
rect 29520 16924 30000 16954
rect 23565 16922 30000 16924
rect 23565 16866 23570 16922
rect 23626 16866 30000 16922
rect 23565 16864 30000 16866
rect 23565 16861 23631 16864
rect 29520 16834 30000 16864
rect 13537 16788 13603 16791
rect 17493 16788 17559 16791
rect 13537 16786 17559 16788
rect 13537 16730 13542 16786
rect 13598 16730 17498 16786
rect 17554 16730 17559 16786
rect 13537 16728 17559 16730
rect 13537 16725 13603 16728
rect 17493 16725 17559 16728
rect 10944 16722 11264 16723
rect 10944 16658 10952 16722
rect 11016 16658 11032 16722
rect 11096 16658 11112 16722
rect 11176 16658 11192 16722
rect 11256 16658 11264 16722
rect 10944 16657 11264 16658
rect 20944 16722 21264 16723
rect 20944 16658 20952 16722
rect 21016 16658 21032 16722
rect 21096 16658 21112 16722
rect 21176 16658 21192 16722
rect 21256 16658 21264 16722
rect 20944 16657 21264 16658
rect 0 16244 480 16274
rect 4061 16244 4127 16247
rect 29520 16244 30000 16274
rect 0 16242 4127 16244
rect 0 16186 4066 16242
rect 4122 16186 4127 16242
rect 0 16184 4127 16186
rect 0 16154 480 16184
rect 4061 16181 4127 16184
rect 27846 16184 30000 16244
rect 5944 16178 6264 16179
rect 5944 16114 5952 16178
rect 6016 16114 6032 16178
rect 6096 16114 6112 16178
rect 6176 16114 6192 16178
rect 6256 16114 6264 16178
rect 5944 16113 6264 16114
rect 15944 16178 16264 16179
rect 15944 16114 15952 16178
rect 16016 16114 16032 16178
rect 16096 16114 16112 16178
rect 16176 16114 16192 16178
rect 16256 16114 16264 16178
rect 15944 16113 16264 16114
rect 25944 16178 26264 16179
rect 25944 16114 25952 16178
rect 26016 16114 26032 16178
rect 26096 16114 26112 16178
rect 26176 16114 26192 16178
rect 26256 16114 26264 16178
rect 25944 16113 26264 16114
rect 25681 15972 25747 15975
rect 27846 15972 27906 16184
rect 29520 16154 30000 16184
rect 25681 15970 27906 15972
rect 25681 15914 25686 15970
rect 25742 15914 27906 15970
rect 25681 15912 27906 15914
rect 25681 15909 25747 15912
rect 7189 15836 7255 15839
rect 9949 15836 10015 15839
rect 7189 15834 10015 15836
rect 7189 15778 7194 15834
rect 7250 15778 9954 15834
rect 10010 15778 10015 15834
rect 7189 15776 10015 15778
rect 7189 15773 7255 15776
rect 9949 15773 10015 15776
rect 0 15700 480 15730
rect 2957 15700 3023 15703
rect 0 15698 3023 15700
rect 0 15642 2962 15698
rect 3018 15642 3023 15698
rect 0 15640 3023 15642
rect 0 15610 480 15640
rect 2957 15637 3023 15640
rect 25497 15700 25563 15703
rect 29520 15700 30000 15730
rect 25497 15698 30000 15700
rect 25497 15642 25502 15698
rect 25558 15642 30000 15698
rect 25497 15640 30000 15642
rect 25497 15637 25563 15640
rect 10944 15634 11264 15635
rect 10944 15570 10952 15634
rect 11016 15570 11032 15634
rect 11096 15570 11112 15634
rect 11176 15570 11192 15634
rect 11256 15570 11264 15634
rect 10944 15569 11264 15570
rect 20944 15634 21264 15635
rect 20944 15570 20952 15634
rect 21016 15570 21032 15634
rect 21096 15570 21112 15634
rect 21176 15570 21192 15634
rect 21256 15570 21264 15634
rect 29520 15610 30000 15640
rect 20944 15569 21264 15570
rect 23933 15292 23999 15295
rect 23933 15290 27906 15292
rect 23933 15234 23938 15290
rect 23994 15234 27906 15290
rect 23933 15232 27906 15234
rect 23933 15229 23999 15232
rect 0 15156 480 15186
rect 1393 15156 1459 15159
rect 0 15154 1459 15156
rect 0 15098 1398 15154
rect 1454 15098 1459 15154
rect 0 15096 1459 15098
rect 27846 15156 27906 15232
rect 29520 15156 30000 15186
rect 27846 15096 30000 15156
rect 0 15066 480 15096
rect 1393 15093 1459 15096
rect 5944 15090 6264 15091
rect 5944 15026 5952 15090
rect 6016 15026 6032 15090
rect 6096 15026 6112 15090
rect 6176 15026 6192 15090
rect 6256 15026 6264 15090
rect 5944 15025 6264 15026
rect 15944 15090 16264 15091
rect 15944 15026 15952 15090
rect 16016 15026 16032 15090
rect 16096 15026 16112 15090
rect 16176 15026 16192 15090
rect 16256 15026 16264 15090
rect 15944 15025 16264 15026
rect 25944 15090 26264 15091
rect 25944 15026 25952 15090
rect 26016 15026 26032 15090
rect 26096 15026 26112 15090
rect 26176 15026 26192 15090
rect 26256 15026 26264 15090
rect 29520 15066 30000 15096
rect 25944 15025 26264 15026
rect 14181 14884 14247 14887
rect 18321 14884 18387 14887
rect 14181 14882 18387 14884
rect 14181 14826 14186 14882
rect 14242 14826 18326 14882
rect 18382 14826 18387 14882
rect 14181 14824 18387 14826
rect 14181 14821 14247 14824
rect 18321 14821 18387 14824
rect 10944 14546 11264 14547
rect 0 14476 480 14506
rect 10944 14482 10952 14546
rect 11016 14482 11032 14546
rect 11096 14482 11112 14546
rect 11176 14482 11192 14546
rect 11256 14482 11264 14546
rect 10944 14481 11264 14482
rect 20944 14546 21264 14547
rect 20944 14482 20952 14546
rect 21016 14482 21032 14546
rect 21096 14482 21112 14546
rect 21176 14482 21192 14546
rect 21256 14482 21264 14546
rect 20944 14481 21264 14482
rect 3417 14476 3483 14479
rect 0 14474 3483 14476
rect 0 14418 3422 14474
rect 3478 14418 3483 14474
rect 0 14416 3483 14418
rect 0 14386 480 14416
rect 3417 14413 3483 14416
rect 25405 14476 25471 14479
rect 29520 14476 30000 14506
rect 25405 14474 30000 14476
rect 25405 14418 25410 14474
rect 25466 14418 30000 14474
rect 25405 14416 30000 14418
rect 25405 14413 25471 14416
rect 29520 14386 30000 14416
rect 5944 14002 6264 14003
rect 0 13932 480 13962
rect 5944 13938 5952 14002
rect 6016 13938 6032 14002
rect 6096 13938 6112 14002
rect 6176 13938 6192 14002
rect 6256 13938 6264 14002
rect 5944 13937 6264 13938
rect 15944 14002 16264 14003
rect 15944 13938 15952 14002
rect 16016 13938 16032 14002
rect 16096 13938 16112 14002
rect 16176 13938 16192 14002
rect 16256 13938 16264 14002
rect 15944 13937 16264 13938
rect 25944 14002 26264 14003
rect 25944 13938 25952 14002
rect 26016 13938 26032 14002
rect 26096 13938 26112 14002
rect 26176 13938 26192 14002
rect 26256 13938 26264 14002
rect 25944 13937 26264 13938
rect 1669 13932 1735 13935
rect 29520 13932 30000 13962
rect 0 13930 1735 13932
rect 0 13874 1674 13930
rect 1730 13874 1735 13930
rect 0 13872 1735 13874
rect 0 13842 480 13872
rect 1669 13869 1735 13872
rect 27846 13872 30000 13932
rect 25313 13796 25379 13799
rect 27846 13796 27906 13872
rect 29520 13842 30000 13872
rect 25313 13794 27906 13796
rect 25313 13738 25318 13794
rect 25374 13738 27906 13794
rect 25313 13736 27906 13738
rect 25313 13733 25379 13736
rect 23105 13660 23171 13663
rect 25589 13660 25655 13663
rect 23105 13658 25655 13660
rect 23105 13602 23110 13658
rect 23166 13602 25594 13658
rect 25650 13602 25655 13658
rect 23105 13600 25655 13602
rect 23105 13597 23171 13600
rect 25589 13597 25655 13600
rect 10944 13458 11264 13459
rect 10944 13394 10952 13458
rect 11016 13394 11032 13458
rect 11096 13394 11112 13458
rect 11176 13394 11192 13458
rect 11256 13394 11264 13458
rect 10944 13393 11264 13394
rect 20944 13458 21264 13459
rect 20944 13394 20952 13458
rect 21016 13394 21032 13458
rect 21096 13394 21112 13458
rect 21176 13394 21192 13458
rect 21256 13394 21264 13458
rect 20944 13393 21264 13394
rect 0 13252 480 13282
rect 1485 13252 1551 13255
rect 19885 13252 19951 13255
rect 0 13192 1410 13252
rect 0 13162 480 13192
rect 1350 13116 1410 13192
rect 1485 13250 19951 13252
rect 1485 13194 1490 13250
rect 1546 13194 19890 13250
rect 19946 13194 19951 13250
rect 1485 13192 19951 13194
rect 1485 13189 1551 13192
rect 19885 13189 19951 13192
rect 25129 13252 25195 13255
rect 29520 13252 30000 13282
rect 25129 13250 30000 13252
rect 25129 13194 25134 13250
rect 25190 13194 30000 13250
rect 25129 13192 30000 13194
rect 25129 13189 25195 13192
rect 29520 13162 30000 13192
rect 3141 13116 3207 13119
rect 1350 13114 3207 13116
rect 1350 13058 3146 13114
rect 3202 13058 3207 13114
rect 1350 13056 3207 13058
rect 3141 13053 3207 13056
rect 3417 13116 3483 13119
rect 11881 13116 11947 13119
rect 3417 13114 11947 13116
rect 3417 13058 3422 13114
rect 3478 13058 11886 13114
rect 11942 13058 11947 13114
rect 3417 13056 11947 13058
rect 3417 13053 3483 13056
rect 11881 13053 11947 13056
rect 19609 13116 19675 13119
rect 23473 13116 23539 13119
rect 19609 13114 23539 13116
rect 19609 13058 19614 13114
rect 19670 13058 23478 13114
rect 23534 13058 23539 13114
rect 19609 13056 23539 13058
rect 19609 13053 19675 13056
rect 23473 13053 23539 13056
rect 5944 12914 6264 12915
rect 5944 12850 5952 12914
rect 6016 12850 6032 12914
rect 6096 12850 6112 12914
rect 6176 12850 6192 12914
rect 6256 12850 6264 12914
rect 5944 12849 6264 12850
rect 15944 12914 16264 12915
rect 15944 12850 15952 12914
rect 16016 12850 16032 12914
rect 16096 12850 16112 12914
rect 16176 12850 16192 12914
rect 16256 12850 16264 12914
rect 15944 12849 16264 12850
rect 25944 12914 26264 12915
rect 25944 12850 25952 12914
rect 26016 12850 26032 12914
rect 26096 12850 26112 12914
rect 26176 12850 26192 12914
rect 26256 12850 26264 12914
rect 25944 12849 26264 12850
rect 0 12708 480 12738
rect 1853 12708 1919 12711
rect 0 12706 1919 12708
rect 0 12650 1858 12706
rect 1914 12650 1919 12706
rect 0 12648 1919 12650
rect 0 12618 480 12648
rect 1853 12645 1919 12648
rect 25589 12708 25655 12711
rect 29520 12708 30000 12738
rect 25589 12706 30000 12708
rect 25589 12650 25594 12706
rect 25650 12650 30000 12706
rect 25589 12648 30000 12650
rect 25589 12645 25655 12648
rect 29520 12618 30000 12648
rect 3233 12572 3299 12575
rect 12893 12572 12959 12575
rect 14641 12572 14707 12575
rect 3233 12570 14707 12572
rect 3233 12514 3238 12570
rect 3294 12514 12898 12570
rect 12954 12514 14646 12570
rect 14702 12514 14707 12570
rect 3233 12512 14707 12514
rect 3233 12509 3299 12512
rect 12893 12509 12959 12512
rect 14641 12509 14707 12512
rect 10944 12370 11264 12371
rect 10944 12306 10952 12370
rect 11016 12306 11032 12370
rect 11096 12306 11112 12370
rect 11176 12306 11192 12370
rect 11256 12306 11264 12370
rect 10944 12305 11264 12306
rect 20944 12370 21264 12371
rect 20944 12306 20952 12370
rect 21016 12306 21032 12370
rect 21096 12306 21112 12370
rect 21176 12306 21192 12370
rect 21256 12306 21264 12370
rect 20944 12305 21264 12306
rect 24485 12300 24551 12303
rect 25221 12300 25287 12303
rect 24485 12298 25287 12300
rect 24485 12242 24490 12298
rect 24546 12242 25226 12298
rect 25282 12242 25287 12298
rect 24485 12240 25287 12242
rect 24485 12237 24551 12240
rect 25221 12237 25287 12240
rect 0 12164 480 12194
rect 3601 12164 3667 12167
rect 0 12162 3667 12164
rect 0 12106 3606 12162
rect 3662 12106 3667 12162
rect 0 12104 3667 12106
rect 0 12074 480 12104
rect 3601 12101 3667 12104
rect 13721 12164 13787 12167
rect 20437 12164 20503 12167
rect 13721 12162 20503 12164
rect 13721 12106 13726 12162
rect 13782 12106 20442 12162
rect 20498 12106 20503 12162
rect 13721 12104 20503 12106
rect 13721 12101 13787 12104
rect 20437 12101 20503 12104
rect 24945 12164 25011 12167
rect 29520 12164 30000 12194
rect 24945 12162 30000 12164
rect 24945 12106 24950 12162
rect 25006 12106 30000 12162
rect 24945 12104 30000 12106
rect 24945 12101 25011 12104
rect 29520 12074 30000 12104
rect 3141 12028 3207 12031
rect 7373 12028 7439 12031
rect 3141 12026 7439 12028
rect 3141 11970 3146 12026
rect 3202 11970 7378 12026
rect 7434 11970 7439 12026
rect 3141 11968 7439 11970
rect 3141 11965 3207 11968
rect 7373 11965 7439 11968
rect 7925 12028 7991 12031
rect 13813 12028 13879 12031
rect 17217 12028 17283 12031
rect 24853 12028 24919 12031
rect 7925 12026 13879 12028
rect 7925 11970 7930 12026
rect 7986 11970 13818 12026
rect 13874 11970 13879 12026
rect 7925 11968 13879 11970
rect 7925 11965 7991 11968
rect 13813 11965 13879 11968
rect 15702 11968 16498 12028
rect 8385 11892 8451 11895
rect 12065 11892 12131 11895
rect 8385 11890 12131 11892
rect 8385 11834 8390 11890
rect 8446 11834 12070 11890
rect 12126 11834 12131 11890
rect 8385 11832 12131 11834
rect 8385 11829 8451 11832
rect 12065 11829 12131 11832
rect 5944 11826 6264 11827
rect 5944 11762 5952 11826
rect 6016 11762 6032 11826
rect 6096 11762 6112 11826
rect 6176 11762 6192 11826
rect 6256 11762 6264 11826
rect 5944 11761 6264 11762
rect 15702 11756 15762 11968
rect 16438 11892 16498 11968
rect 17217 12026 24919 12028
rect 17217 11970 17222 12026
rect 17278 11970 24858 12026
rect 24914 11970 24919 12026
rect 17217 11968 24919 11970
rect 17217 11965 17283 11968
rect 24853 11965 24919 11968
rect 23381 11892 23447 11895
rect 16438 11890 23447 11892
rect 16438 11834 23386 11890
rect 23442 11834 23447 11890
rect 16438 11832 23447 11834
rect 23381 11829 23447 11832
rect 24669 11892 24735 11895
rect 25037 11892 25103 11895
rect 24669 11890 25103 11892
rect 24669 11834 24674 11890
rect 24730 11834 25042 11890
rect 25098 11834 25103 11890
rect 24669 11832 25103 11834
rect 24669 11829 24735 11832
rect 25037 11829 25103 11832
rect 15944 11826 16264 11827
rect 15944 11762 15952 11826
rect 16016 11762 16032 11826
rect 16096 11762 16112 11826
rect 16176 11762 16192 11826
rect 16256 11762 16264 11826
rect 15944 11761 16264 11762
rect 25944 11826 26264 11827
rect 25944 11762 25952 11826
rect 26016 11762 26032 11826
rect 26096 11762 26112 11826
rect 26176 11762 26192 11826
rect 26256 11762 26264 11826
rect 25944 11761 26264 11762
rect 25405 11756 25471 11759
rect 6502 11696 15762 11756
rect 17358 11754 25471 11756
rect 17358 11698 25410 11754
rect 25466 11698 25471 11754
rect 17358 11696 25471 11698
rect 3417 11620 3483 11623
rect 6502 11620 6562 11696
rect 3417 11618 6562 11620
rect 3417 11562 3422 11618
rect 3478 11562 6562 11618
rect 3417 11560 6562 11562
rect 6637 11620 6703 11623
rect 11513 11620 11579 11623
rect 6637 11618 11579 11620
rect 6637 11562 6642 11618
rect 6698 11562 11518 11618
rect 11574 11562 11579 11618
rect 6637 11560 11579 11562
rect 3417 11557 3483 11560
rect 6637 11557 6703 11560
rect 11513 11557 11579 11560
rect 0 11484 480 11514
rect 13721 11484 13787 11487
rect 17358 11484 17418 11696
rect 25405 11693 25471 11696
rect 17493 11620 17559 11623
rect 25313 11620 25379 11623
rect 17493 11618 25379 11620
rect 17493 11562 17498 11618
rect 17554 11562 25318 11618
rect 25374 11562 25379 11618
rect 17493 11560 25379 11562
rect 17493 11557 17559 11560
rect 25313 11557 25379 11560
rect 0 11424 11714 11484
rect 0 11394 480 11424
rect 2405 11348 2471 11351
rect 6637 11348 6703 11351
rect 2405 11346 6703 11348
rect 2405 11290 2410 11346
rect 2466 11290 6642 11346
rect 6698 11290 6703 11346
rect 2405 11288 6703 11290
rect 11654 11348 11714 11424
rect 13721 11482 17418 11484
rect 13721 11426 13726 11482
rect 13782 11426 17418 11482
rect 13721 11424 17418 11426
rect 24117 11484 24183 11487
rect 29520 11484 30000 11514
rect 24117 11482 30000 11484
rect 24117 11426 24122 11482
rect 24178 11426 30000 11482
rect 24117 11424 30000 11426
rect 13721 11421 13787 11424
rect 24117 11421 24183 11424
rect 29520 11394 30000 11424
rect 17217 11348 17283 11351
rect 11654 11346 17283 11348
rect 11654 11290 17222 11346
rect 17278 11290 17283 11346
rect 11654 11288 17283 11290
rect 2405 11285 2471 11288
rect 6637 11285 6703 11288
rect 17217 11285 17283 11288
rect 10944 11282 11264 11283
rect 10944 11218 10952 11282
rect 11016 11218 11032 11282
rect 11096 11218 11112 11282
rect 11176 11218 11192 11282
rect 11256 11218 11264 11282
rect 10944 11217 11264 11218
rect 20944 11282 21264 11283
rect 20944 11218 20952 11282
rect 21016 11218 21032 11282
rect 21096 11218 21112 11282
rect 21176 11218 21192 11282
rect 21256 11218 21264 11282
rect 20944 11217 21264 11218
rect 2497 11212 2563 11215
rect 7097 11212 7163 11215
rect 2497 11210 7163 11212
rect 2497 11154 2502 11210
rect 2558 11154 7102 11210
rect 7158 11154 7163 11210
rect 2497 11152 7163 11154
rect 2497 11149 2563 11152
rect 7097 11149 7163 11152
rect 12433 11212 12499 11215
rect 12433 11210 17786 11212
rect 12433 11154 12438 11210
rect 12494 11154 17786 11210
rect 12433 11152 17786 11154
rect 12433 11149 12499 11152
rect 2037 11076 2103 11079
rect 17493 11076 17559 11079
rect 2037 11074 17559 11076
rect 2037 11018 2042 11074
rect 2098 11018 17498 11074
rect 17554 11018 17559 11074
rect 2037 11016 17559 11018
rect 17726 11076 17786 11152
rect 25129 11076 25195 11079
rect 17726 11074 25195 11076
rect 17726 11018 25134 11074
rect 25190 11018 25195 11074
rect 17726 11016 25195 11018
rect 2037 11013 2103 11016
rect 17493 11013 17559 11016
rect 25129 11013 25195 11016
rect 0 10940 480 10970
rect 3417 10940 3483 10943
rect 0 10938 3483 10940
rect 0 10882 3422 10938
rect 3478 10882 3483 10938
rect 0 10880 3483 10882
rect 0 10850 480 10880
rect 3417 10877 3483 10880
rect 8109 10940 8175 10943
rect 12433 10940 12499 10943
rect 8109 10938 12499 10940
rect 8109 10882 8114 10938
rect 8170 10882 12438 10938
rect 12494 10882 12499 10938
rect 8109 10880 12499 10882
rect 8109 10877 8175 10880
rect 12433 10877 12499 10880
rect 24761 10940 24827 10943
rect 29520 10940 30000 10970
rect 24761 10938 30000 10940
rect 24761 10882 24766 10938
rect 24822 10882 30000 10938
rect 24761 10880 30000 10882
rect 24761 10877 24827 10880
rect 29520 10850 30000 10880
rect 5944 10738 6264 10739
rect 5944 10674 5952 10738
rect 6016 10674 6032 10738
rect 6096 10674 6112 10738
rect 6176 10674 6192 10738
rect 6256 10674 6264 10738
rect 5944 10673 6264 10674
rect 15944 10738 16264 10739
rect 15944 10674 15952 10738
rect 16016 10674 16032 10738
rect 16096 10674 16112 10738
rect 16176 10674 16192 10738
rect 16256 10674 16264 10738
rect 15944 10673 16264 10674
rect 25944 10738 26264 10739
rect 25944 10674 25952 10738
rect 26016 10674 26032 10738
rect 26096 10674 26112 10738
rect 26176 10674 26192 10738
rect 26256 10674 26264 10738
rect 25944 10673 26264 10674
rect 24117 10532 24183 10535
rect 3374 10530 24183 10532
rect 3374 10474 24122 10530
rect 24178 10474 24183 10530
rect 3374 10472 24183 10474
rect 0 10260 480 10290
rect 3374 10260 3434 10472
rect 24117 10469 24183 10472
rect 8293 10396 8359 10399
rect 24945 10396 25011 10399
rect 8293 10394 25011 10396
rect 8293 10338 8298 10394
rect 8354 10338 24950 10394
rect 25006 10338 25011 10394
rect 8293 10336 25011 10338
rect 8293 10333 8359 10336
rect 24945 10333 25011 10336
rect 0 10200 3434 10260
rect 25037 10260 25103 10263
rect 29520 10260 30000 10290
rect 25037 10258 30000 10260
rect 25037 10202 25042 10258
rect 25098 10202 30000 10258
rect 25037 10200 30000 10202
rect 0 10170 480 10200
rect 25037 10197 25103 10200
rect 10944 10194 11264 10195
rect 10944 10130 10952 10194
rect 11016 10130 11032 10194
rect 11096 10130 11112 10194
rect 11176 10130 11192 10194
rect 11256 10130 11264 10194
rect 10944 10129 11264 10130
rect 20944 10194 21264 10195
rect 20944 10130 20952 10194
rect 21016 10130 21032 10194
rect 21096 10130 21112 10194
rect 21176 10130 21192 10194
rect 21256 10130 21264 10194
rect 29520 10170 30000 10200
rect 20944 10129 21264 10130
rect 3601 10124 3667 10127
rect 7833 10124 7899 10127
rect 3601 10122 7899 10124
rect 3601 10066 3606 10122
rect 3662 10066 7838 10122
rect 7894 10066 7899 10122
rect 3601 10064 7899 10066
rect 3601 10061 3667 10064
rect 7833 10061 7899 10064
rect 1393 9988 1459 9991
rect 8293 9988 8359 9991
rect 1393 9986 8359 9988
rect 1393 9930 1398 9986
rect 1454 9930 8298 9986
rect 8354 9930 8359 9986
rect 1393 9928 8359 9930
rect 1393 9925 1459 9928
rect 8293 9925 8359 9928
rect 2037 9852 2103 9855
rect 19701 9852 19767 9855
rect 2037 9850 19767 9852
rect 2037 9794 2042 9850
rect 2098 9794 19706 9850
rect 19762 9794 19767 9850
rect 2037 9792 19767 9794
rect 2037 9789 2103 9792
rect 19701 9789 19767 9792
rect 24853 9852 24919 9855
rect 24853 9850 27906 9852
rect 24853 9794 24858 9850
rect 24914 9794 27906 9850
rect 24853 9792 27906 9794
rect 24853 9789 24919 9792
rect 0 9716 480 9746
rect 1577 9716 1643 9719
rect 0 9714 1643 9716
rect 0 9658 1582 9714
rect 1638 9658 1643 9714
rect 0 9656 1643 9658
rect 27846 9716 27906 9792
rect 29520 9716 30000 9746
rect 27846 9656 30000 9716
rect 0 9626 480 9656
rect 1577 9653 1643 9656
rect 5944 9650 6264 9651
rect 5944 9586 5952 9650
rect 6016 9586 6032 9650
rect 6096 9586 6112 9650
rect 6176 9586 6192 9650
rect 6256 9586 6264 9650
rect 5944 9585 6264 9586
rect 15944 9650 16264 9651
rect 15944 9586 15952 9650
rect 16016 9586 16032 9650
rect 16096 9586 16112 9650
rect 16176 9586 16192 9650
rect 16256 9586 16264 9650
rect 15944 9585 16264 9586
rect 25944 9650 26264 9651
rect 25944 9586 25952 9650
rect 26016 9586 26032 9650
rect 26096 9586 26112 9650
rect 26176 9586 26192 9650
rect 26256 9586 26264 9650
rect 29520 9626 30000 9656
rect 25944 9585 26264 9586
rect 23657 9444 23723 9447
rect 3374 9442 23723 9444
rect 3374 9386 23662 9442
rect 23718 9386 23723 9442
rect 3374 9384 23723 9386
rect 0 9172 480 9202
rect 3374 9172 3434 9384
rect 23657 9381 23723 9384
rect 3693 9308 3759 9311
rect 23933 9308 23999 9311
rect 3693 9306 23999 9308
rect 3693 9250 3698 9306
rect 3754 9250 23938 9306
rect 23994 9250 23999 9306
rect 3693 9248 23999 9250
rect 3693 9245 3759 9248
rect 23933 9245 23999 9248
rect 0 9112 3434 9172
rect 24117 9172 24183 9175
rect 29520 9172 30000 9202
rect 24117 9170 30000 9172
rect 24117 9114 24122 9170
rect 24178 9114 30000 9170
rect 24117 9112 30000 9114
rect 0 9082 480 9112
rect 24117 9109 24183 9112
rect 10944 9106 11264 9107
rect 10944 9042 10952 9106
rect 11016 9042 11032 9106
rect 11096 9042 11112 9106
rect 11176 9042 11192 9106
rect 11256 9042 11264 9106
rect 10944 9041 11264 9042
rect 20944 9106 21264 9107
rect 20944 9042 20952 9106
rect 21016 9042 21032 9106
rect 21096 9042 21112 9106
rect 21176 9042 21192 9106
rect 21256 9042 21264 9106
rect 29520 9082 30000 9112
rect 20944 9041 21264 9042
rect 3325 9036 3391 9039
rect 4797 9036 4863 9039
rect 3325 9034 4863 9036
rect 3325 8978 3330 9034
rect 3386 8978 4802 9034
rect 4858 8978 4863 9034
rect 3325 8976 4863 8978
rect 3325 8973 3391 8976
rect 4797 8973 4863 8976
rect 23749 8900 23815 8903
rect 3558 8898 23815 8900
rect 3558 8842 23754 8898
rect 23810 8842 23815 8898
rect 3558 8840 23815 8842
rect 0 8492 480 8522
rect 3558 8492 3618 8840
rect 23749 8837 23815 8840
rect 5944 8562 6264 8563
rect 5944 8498 5952 8562
rect 6016 8498 6032 8562
rect 6096 8498 6112 8562
rect 6176 8498 6192 8562
rect 6256 8498 6264 8562
rect 5944 8497 6264 8498
rect 15944 8562 16264 8563
rect 15944 8498 15952 8562
rect 16016 8498 16032 8562
rect 16096 8498 16112 8562
rect 16176 8498 16192 8562
rect 16256 8498 16264 8562
rect 15944 8497 16264 8498
rect 25944 8562 26264 8563
rect 25944 8498 25952 8562
rect 26016 8498 26032 8562
rect 26096 8498 26112 8562
rect 26176 8498 26192 8562
rect 26256 8498 26264 8562
rect 25944 8497 26264 8498
rect 29520 8492 30000 8522
rect 0 8432 3618 8492
rect 27846 8432 30000 8492
rect 0 8402 480 8432
rect 24117 8356 24183 8359
rect 27846 8356 27906 8432
rect 29520 8402 30000 8432
rect 24117 8354 27906 8356
rect 24117 8298 24122 8354
rect 24178 8298 27906 8354
rect 24117 8296 27906 8298
rect 24117 8293 24183 8296
rect 3969 8220 4035 8223
rect 24485 8220 24551 8223
rect 3969 8218 24551 8220
rect 3969 8162 3974 8218
rect 4030 8162 24490 8218
rect 24546 8162 24551 8218
rect 3969 8160 24551 8162
rect 3969 8157 4035 8160
rect 24485 8157 24551 8160
rect 3049 8084 3115 8087
rect 3601 8084 3667 8087
rect 10777 8084 10843 8087
rect 3049 8082 3667 8084
rect 3049 8026 3054 8082
rect 3110 8026 3606 8082
rect 3662 8026 3667 8082
rect 3049 8024 3667 8026
rect 3049 8021 3115 8024
rect 3601 8021 3667 8024
rect 3742 8082 10843 8084
rect 3742 8026 10782 8082
rect 10838 8026 10843 8082
rect 3742 8024 10843 8026
rect 0 7948 480 7978
rect 3742 7948 3802 8024
rect 10777 8021 10843 8024
rect 11329 8084 11395 8087
rect 11329 8082 17234 8084
rect 11329 8026 11334 8082
rect 11390 8026 17234 8082
rect 11329 8024 17234 8026
rect 11329 8021 11395 8024
rect 10944 8018 11264 8019
rect 10944 7954 10952 8018
rect 11016 7954 11032 8018
rect 11096 7954 11112 8018
rect 11176 7954 11192 8018
rect 11256 7954 11264 8018
rect 10944 7953 11264 7954
rect 0 7888 3802 7948
rect 0 7858 480 7888
rect 3693 7812 3759 7815
rect 17174 7812 17234 8024
rect 20944 8018 21264 8019
rect 20944 7954 20952 8018
rect 21016 7954 21032 8018
rect 21096 7954 21112 8018
rect 21176 7954 21192 8018
rect 21256 7954 21264 8018
rect 20944 7953 21264 7954
rect 24117 7948 24183 7951
rect 29520 7948 30000 7978
rect 24117 7946 30000 7948
rect 24117 7890 24122 7946
rect 24178 7890 30000 7946
rect 24117 7888 30000 7890
rect 24117 7885 24183 7888
rect 29520 7858 30000 7888
rect 23473 7812 23539 7815
rect 3693 7810 17050 7812
rect 3693 7754 3698 7810
rect 3754 7754 17050 7810
rect 3693 7752 17050 7754
rect 17174 7810 23539 7812
rect 17174 7754 23478 7810
rect 23534 7754 23539 7810
rect 17174 7752 23539 7754
rect 3693 7749 3759 7752
rect 3601 7676 3667 7679
rect 10869 7676 10935 7679
rect 3601 7674 10935 7676
rect 3601 7618 3606 7674
rect 3662 7618 10874 7674
rect 10930 7618 10935 7674
rect 3601 7616 10935 7618
rect 3601 7613 3667 7616
rect 10869 7613 10935 7616
rect 16990 7540 17050 7752
rect 23473 7749 23539 7752
rect 22645 7540 22711 7543
rect 16990 7538 22711 7540
rect 16990 7482 22650 7538
rect 22706 7482 22711 7538
rect 16990 7480 22711 7482
rect 22645 7477 22711 7480
rect 5944 7474 6264 7475
rect 5944 7410 5952 7474
rect 6016 7410 6032 7474
rect 6096 7410 6112 7474
rect 6176 7410 6192 7474
rect 6256 7410 6264 7474
rect 5944 7409 6264 7410
rect 15944 7474 16264 7475
rect 15944 7410 15952 7474
rect 16016 7410 16032 7474
rect 16096 7410 16112 7474
rect 16176 7410 16192 7474
rect 16256 7410 16264 7474
rect 15944 7409 16264 7410
rect 25944 7474 26264 7475
rect 25944 7410 25952 7474
rect 26016 7410 26032 7474
rect 26096 7410 26112 7474
rect 26176 7410 26192 7474
rect 26256 7410 26264 7474
rect 25944 7409 26264 7410
rect 0 7268 480 7298
rect 3693 7268 3759 7271
rect 0 7266 3759 7268
rect 0 7210 3698 7266
rect 3754 7210 3759 7266
rect 0 7208 3759 7210
rect 0 7178 480 7208
rect 3693 7205 3759 7208
rect 3877 7268 3943 7271
rect 18689 7268 18755 7271
rect 3877 7266 18755 7268
rect 3877 7210 3882 7266
rect 3938 7210 18694 7266
rect 18750 7210 18755 7266
rect 3877 7208 18755 7210
rect 3877 7205 3943 7208
rect 18689 7205 18755 7208
rect 18873 7268 18939 7271
rect 29520 7268 30000 7298
rect 18873 7266 30000 7268
rect 18873 7210 18878 7266
rect 18934 7210 30000 7266
rect 18873 7208 30000 7210
rect 18873 7205 18939 7208
rect 29520 7178 30000 7208
rect 3785 7132 3851 7135
rect 23933 7132 23999 7135
rect 3785 7130 23999 7132
rect 3785 7074 3790 7130
rect 3846 7074 23938 7130
rect 23994 7074 23999 7130
rect 3785 7072 23999 7074
rect 3785 7069 3851 7072
rect 23933 7069 23999 7072
rect 10944 6930 11264 6931
rect 10944 6866 10952 6930
rect 11016 6866 11032 6930
rect 11096 6866 11112 6930
rect 11176 6866 11192 6930
rect 11256 6866 11264 6930
rect 10944 6865 11264 6866
rect 20944 6930 21264 6931
rect 20944 6866 20952 6930
rect 21016 6866 21032 6930
rect 21096 6866 21112 6930
rect 21176 6866 21192 6930
rect 21256 6866 21264 6930
rect 20944 6865 21264 6866
rect 0 6724 480 6754
rect 29520 6724 30000 6754
rect 0 6664 674 6724
rect 0 6634 480 6664
rect 614 6588 674 6664
rect 24534 6664 30000 6724
rect 24117 6588 24183 6591
rect 614 6586 24183 6588
rect 614 6530 24122 6586
rect 24178 6530 24183 6586
rect 614 6528 24183 6530
rect 24117 6525 24183 6528
rect 17217 6452 17283 6455
rect 24534 6452 24594 6664
rect 29520 6634 30000 6664
rect 17217 6450 24594 6452
rect 17217 6394 17222 6450
rect 17278 6394 24594 6450
rect 17217 6392 24594 6394
rect 17217 6389 17283 6392
rect 5944 6386 6264 6387
rect 5944 6322 5952 6386
rect 6016 6322 6032 6386
rect 6096 6322 6112 6386
rect 6176 6322 6192 6386
rect 6256 6322 6264 6386
rect 5944 6321 6264 6322
rect 15944 6386 16264 6387
rect 15944 6322 15952 6386
rect 16016 6322 16032 6386
rect 16096 6322 16112 6386
rect 16176 6322 16192 6386
rect 16256 6322 16264 6386
rect 15944 6321 16264 6322
rect 25944 6386 26264 6387
rect 25944 6322 25952 6386
rect 26016 6322 26032 6386
rect 26096 6322 26112 6386
rect 26176 6322 26192 6386
rect 26256 6322 26264 6386
rect 25944 6321 26264 6322
rect 0 6180 480 6210
rect 2129 6180 2195 6183
rect 0 6178 2195 6180
rect 0 6122 2134 6178
rect 2190 6122 2195 6178
rect 0 6120 2195 6122
rect 0 6090 480 6120
rect 2129 6117 2195 6120
rect 11053 6180 11119 6183
rect 14825 6180 14891 6183
rect 29520 6180 30000 6210
rect 11053 6178 14704 6180
rect 11053 6122 11058 6178
rect 11114 6122 14704 6178
rect 11053 6120 14704 6122
rect 11053 6117 11119 6120
rect 12801 6044 12867 6047
rect 3190 6042 12867 6044
rect 3190 5986 12806 6042
rect 12862 5986 12867 6042
rect 3190 5984 12867 5986
rect 14644 6044 14704 6120
rect 14825 6178 30000 6180
rect 14825 6122 14830 6178
rect 14886 6122 30000 6178
rect 14825 6120 30000 6122
rect 14825 6117 14891 6120
rect 29520 6090 30000 6120
rect 17217 6044 17283 6047
rect 14644 6042 17283 6044
rect 14644 5986 17222 6042
rect 17278 5986 17283 6042
rect 14644 5984 17283 5986
rect 0 5500 480 5530
rect 3190 5500 3250 5984
rect 12801 5981 12867 5984
rect 17217 5981 17283 5984
rect 10944 5842 11264 5843
rect 10944 5778 10952 5842
rect 11016 5778 11032 5842
rect 11096 5778 11112 5842
rect 11176 5778 11192 5842
rect 11256 5778 11264 5842
rect 10944 5777 11264 5778
rect 20944 5842 21264 5843
rect 20944 5778 20952 5842
rect 21016 5778 21032 5842
rect 21096 5778 21112 5842
rect 21176 5778 21192 5842
rect 21256 5778 21264 5842
rect 20944 5777 21264 5778
rect 12617 5636 12683 5639
rect 25773 5636 25839 5639
rect 12617 5634 25839 5636
rect 12617 5578 12622 5634
rect 12678 5578 25778 5634
rect 25834 5578 25839 5634
rect 12617 5576 25839 5578
rect 12617 5573 12683 5576
rect 25773 5573 25839 5576
rect 0 5440 3250 5500
rect 4981 5500 5047 5503
rect 29520 5500 30000 5530
rect 4981 5498 30000 5500
rect 4981 5442 4986 5498
rect 5042 5442 30000 5498
rect 4981 5440 30000 5442
rect 0 5410 480 5440
rect 4981 5437 5047 5440
rect 29520 5410 30000 5440
rect 5944 5298 6264 5299
rect 5944 5234 5952 5298
rect 6016 5234 6032 5298
rect 6096 5234 6112 5298
rect 6176 5234 6192 5298
rect 6256 5234 6264 5298
rect 5944 5233 6264 5234
rect 15944 5298 16264 5299
rect 15944 5234 15952 5298
rect 16016 5234 16032 5298
rect 16096 5234 16112 5298
rect 16176 5234 16192 5298
rect 16256 5234 16264 5298
rect 15944 5233 16264 5234
rect 25944 5298 26264 5299
rect 25944 5234 25952 5298
rect 26016 5234 26032 5298
rect 26096 5234 26112 5298
rect 26176 5234 26192 5298
rect 26256 5234 26264 5298
rect 25944 5233 26264 5234
rect 16389 5228 16455 5231
rect 16389 5226 24410 5228
rect 16389 5170 16394 5226
rect 16450 5170 24410 5226
rect 16389 5168 24410 5170
rect 16389 5165 16455 5168
rect 3509 5092 3575 5095
rect 13721 5092 13787 5095
rect 3509 5090 13787 5092
rect 3509 5034 3514 5090
rect 3570 5034 13726 5090
rect 13782 5034 13787 5090
rect 3509 5032 13787 5034
rect 3509 5029 3575 5032
rect 13721 5029 13787 5032
rect 0 4956 480 4986
rect 24117 4956 24183 4959
rect 0 4954 24183 4956
rect 0 4898 24122 4954
rect 24178 4898 24183 4954
rect 0 4896 24183 4898
rect 24350 4956 24410 5168
rect 29520 4956 30000 4986
rect 24350 4896 30000 4956
rect 0 4866 480 4896
rect 24117 4893 24183 4896
rect 29520 4866 30000 4896
rect 10944 4754 11264 4755
rect 10944 4690 10952 4754
rect 11016 4690 11032 4754
rect 11096 4690 11112 4754
rect 11176 4690 11192 4754
rect 11256 4690 11264 4754
rect 10944 4689 11264 4690
rect 20944 4754 21264 4755
rect 20944 4690 20952 4754
rect 21016 4690 21032 4754
rect 21096 4690 21112 4754
rect 21176 4690 21192 4754
rect 21256 4690 21264 4754
rect 20944 4689 21264 4690
rect 3877 4548 3943 4551
rect 20713 4548 20779 4551
rect 3877 4546 20779 4548
rect 3877 4490 3882 4546
rect 3938 4490 20718 4546
rect 20774 4490 20779 4546
rect 3877 4488 20779 4490
rect 3877 4485 3943 4488
rect 20713 4485 20779 4488
rect 16481 4412 16547 4415
rect 2638 4410 16547 4412
rect 2638 4354 16486 4410
rect 16542 4354 16547 4410
rect 2638 4352 16547 4354
rect 0 4276 480 4306
rect 2638 4276 2698 4352
rect 16481 4349 16547 4352
rect 20897 4412 20963 4415
rect 20897 4410 27906 4412
rect 20897 4354 20902 4410
rect 20958 4354 27906 4410
rect 20897 4352 27906 4354
rect 20897 4349 20963 4352
rect 0 4216 2698 4276
rect 27846 4276 27906 4352
rect 29520 4276 30000 4306
rect 27846 4216 30000 4276
rect 0 4186 480 4216
rect 5944 4210 6264 4211
rect 5944 4146 5952 4210
rect 6016 4146 6032 4210
rect 6096 4146 6112 4210
rect 6176 4146 6192 4210
rect 6256 4146 6264 4210
rect 5944 4145 6264 4146
rect 15944 4210 16264 4211
rect 15944 4146 15952 4210
rect 16016 4146 16032 4210
rect 16096 4146 16112 4210
rect 16176 4146 16192 4210
rect 16256 4146 16264 4210
rect 15944 4145 16264 4146
rect 25944 4210 26264 4211
rect 25944 4146 25952 4210
rect 26016 4146 26032 4210
rect 26096 4146 26112 4210
rect 26176 4146 26192 4210
rect 26256 4146 26264 4210
rect 29520 4186 30000 4216
rect 25944 4145 26264 4146
rect 16389 4004 16455 4007
rect 25681 4004 25747 4007
rect 16389 4002 25747 4004
rect 16389 3946 16394 4002
rect 16450 3946 25686 4002
rect 25742 3946 25747 4002
rect 16389 3944 25747 3946
rect 16389 3941 16455 3944
rect 25681 3941 25747 3944
rect 3417 3868 3483 3871
rect 23933 3868 23999 3871
rect 3417 3866 23999 3868
rect 3417 3810 3422 3866
rect 3478 3810 23938 3866
rect 23994 3810 23999 3866
rect 3417 3808 23999 3810
rect 3417 3805 3483 3808
rect 23933 3805 23999 3808
rect 0 3732 480 3762
rect 24117 3732 24183 3735
rect 29520 3732 30000 3762
rect 0 3672 674 3732
rect 0 3642 480 3672
rect 614 3460 674 3672
rect 24117 3730 30000 3732
rect 24117 3674 24122 3730
rect 24178 3674 30000 3730
rect 24117 3672 30000 3674
rect 24117 3669 24183 3672
rect 10944 3666 11264 3667
rect 10944 3602 10952 3666
rect 11016 3602 11032 3666
rect 11096 3602 11112 3666
rect 11176 3602 11192 3666
rect 11256 3602 11264 3666
rect 10944 3601 11264 3602
rect 20944 3666 21264 3667
rect 20944 3602 20952 3666
rect 21016 3602 21032 3666
rect 21096 3602 21112 3666
rect 21176 3602 21192 3666
rect 21256 3602 21264 3666
rect 29520 3642 30000 3672
rect 20944 3601 21264 3602
rect 22093 3596 22159 3599
rect 25497 3596 25563 3599
rect 22093 3594 25563 3596
rect 22093 3538 22098 3594
rect 22154 3538 25502 3594
rect 25558 3538 25563 3594
rect 22093 3536 25563 3538
rect 22093 3533 22159 3536
rect 25497 3533 25563 3536
rect 21633 3460 21699 3463
rect 614 3458 21699 3460
rect 614 3402 21638 3458
rect 21694 3402 21699 3458
rect 614 3400 21699 3402
rect 21633 3397 21699 3400
rect 24117 3324 24183 3327
rect 2638 3322 24183 3324
rect 2638 3266 24122 3322
rect 24178 3266 24183 3322
rect 2638 3264 24183 3266
rect 0 3188 480 3218
rect 2638 3188 2698 3264
rect 24117 3261 24183 3264
rect 29520 3188 30000 3218
rect 0 3128 2698 3188
rect 27846 3128 30000 3188
rect 0 3098 480 3128
rect 5944 3122 6264 3123
rect 5944 3058 5952 3122
rect 6016 3058 6032 3122
rect 6096 3058 6112 3122
rect 6176 3058 6192 3122
rect 6256 3058 6264 3122
rect 5944 3057 6264 3058
rect 15944 3122 16264 3123
rect 15944 3058 15952 3122
rect 16016 3058 16032 3122
rect 16096 3058 16112 3122
rect 16176 3058 16192 3122
rect 16256 3058 16264 3122
rect 15944 3057 16264 3058
rect 25944 3122 26264 3123
rect 25944 3058 25952 3122
rect 26016 3058 26032 3122
rect 26096 3058 26112 3122
rect 26176 3058 26192 3122
rect 26256 3058 26264 3122
rect 25944 3057 26264 3058
rect 7373 2916 7439 2919
rect 23933 2916 23999 2919
rect 7373 2914 23999 2916
rect 7373 2858 7378 2914
rect 7434 2858 23938 2914
rect 23994 2858 23999 2914
rect 7373 2856 23999 2858
rect 7373 2853 7439 2856
rect 23933 2853 23999 2856
rect 1853 2780 1919 2783
rect 27846 2780 27906 3128
rect 29520 3098 30000 3128
rect 1853 2778 27906 2780
rect 1853 2722 1858 2778
rect 1914 2722 27906 2778
rect 1853 2720 27906 2722
rect 1853 2717 1919 2720
rect 10944 2578 11264 2579
rect 0 2508 480 2538
rect 10944 2514 10952 2578
rect 11016 2514 11032 2578
rect 11096 2514 11112 2578
rect 11176 2514 11192 2578
rect 11256 2514 11264 2578
rect 10944 2513 11264 2514
rect 20944 2578 21264 2579
rect 20944 2514 20952 2578
rect 21016 2514 21032 2578
rect 21096 2514 21112 2578
rect 21176 2514 21192 2578
rect 21256 2514 21264 2578
rect 20944 2513 21264 2514
rect 1761 2508 1827 2511
rect 0 2506 1827 2508
rect 0 2450 1766 2506
rect 1822 2450 1827 2506
rect 0 2448 1827 2450
rect 0 2418 480 2448
rect 1761 2445 1827 2448
rect 24209 2508 24275 2511
rect 29520 2508 30000 2538
rect 24209 2506 30000 2508
rect 24209 2450 24214 2506
rect 24270 2450 30000 2506
rect 24209 2448 30000 2450
rect 24209 2445 24275 2448
rect 29520 2418 30000 2448
rect 2037 2372 2103 2375
rect 25589 2372 25655 2375
rect 2037 2370 25655 2372
rect 2037 2314 2042 2370
rect 2098 2314 25594 2370
rect 25650 2314 25655 2370
rect 2037 2312 25655 2314
rect 2037 2309 2103 2312
rect 25589 2309 25655 2312
rect 12525 2236 12591 2239
rect 24025 2236 24091 2239
rect 12525 2234 24091 2236
rect 12525 2178 12530 2234
rect 12586 2178 24030 2234
rect 24086 2178 24091 2234
rect 12525 2176 24091 2178
rect 12525 2173 12591 2176
rect 24025 2173 24091 2176
rect 5944 2034 6264 2035
rect 0 1964 480 1994
rect 5944 1970 5952 2034
rect 6016 1970 6032 2034
rect 6096 1970 6112 2034
rect 6176 1970 6192 2034
rect 6256 1970 6264 2034
rect 5944 1969 6264 1970
rect 15944 2034 16264 2035
rect 15944 1970 15952 2034
rect 16016 1970 16032 2034
rect 16096 1970 16112 2034
rect 16176 1970 16192 2034
rect 16256 1970 16264 2034
rect 15944 1969 16264 1970
rect 25944 2034 26264 2035
rect 25944 1970 25952 2034
rect 26016 1970 26032 2034
rect 26096 1970 26112 2034
rect 26176 1970 26192 2034
rect 26256 1970 26264 2034
rect 25944 1969 26264 1970
rect 1945 1964 2011 1967
rect 29520 1964 30000 1994
rect 0 1962 2011 1964
rect 0 1906 1950 1962
rect 2006 1906 2011 1962
rect 0 1904 2011 1906
rect 0 1874 480 1904
rect 1945 1901 2011 1904
rect 26926 1904 30000 1964
rect 8385 1828 8451 1831
rect 25129 1828 25195 1831
rect 8385 1826 25195 1828
rect 8385 1770 8390 1826
rect 8446 1770 25134 1826
rect 25190 1770 25195 1826
rect 8385 1768 25195 1770
rect 8385 1765 8451 1768
rect 25129 1765 25195 1768
rect 26926 1692 26986 1904
rect 29520 1874 30000 1904
rect 21958 1632 26986 1692
rect 2221 1556 2287 1559
rect 21958 1556 22018 1632
rect 2221 1554 7666 1556
rect 2221 1498 2226 1554
rect 2282 1498 7666 1554
rect 2221 1496 7666 1498
rect 2221 1493 2287 1496
rect 7606 1420 7666 1496
rect 12390 1496 22018 1556
rect 12390 1420 12450 1496
rect 7606 1360 12450 1420
rect 24853 1420 24919 1423
rect 24853 1418 29378 1420
rect 24853 1362 24858 1418
rect 24914 1362 29378 1418
rect 24853 1360 29378 1362
rect 24853 1357 24919 1360
rect 0 1284 480 1314
rect 1669 1284 1735 1287
rect 0 1282 1735 1284
rect 0 1226 1674 1282
rect 1730 1226 1735 1282
rect 0 1224 1735 1226
rect 29318 1284 29378 1360
rect 29520 1284 30000 1314
rect 29318 1224 30000 1284
rect 0 1194 480 1224
rect 1669 1221 1735 1224
rect 29520 1194 30000 1224
rect 0 740 480 770
rect 1577 740 1643 743
rect 29520 740 30000 770
rect 0 738 1643 740
rect 0 682 1582 738
rect 1638 682 1643 738
rect 0 680 1643 682
rect 0 650 480 680
rect 1577 677 1643 680
rect 29318 680 30000 740
rect 29318 332 29378 680
rect 29520 650 30000 680
rect 21958 272 29378 332
rect 0 196 480 226
rect 1485 196 1551 199
rect 0 194 1551 196
rect 0 138 1490 194
rect 1546 138 1551 194
rect 0 136 1551 138
rect 0 106 480 136
rect 1485 133 1551 136
rect 2681 196 2747 199
rect 21958 196 22018 272
rect 2681 194 7666 196
rect 2681 138 2686 194
rect 2742 138 7666 194
rect 2681 136 7666 138
rect 2681 133 2747 136
rect 7606 60 7666 136
rect 12390 136 22018 196
rect 25313 196 25379 199
rect 29520 196 30000 226
rect 25313 194 30000 196
rect 25313 138 25318 194
rect 25374 138 30000 194
rect 25313 136 30000 138
rect 12390 60 12450 136
rect 25313 133 25379 136
rect 29520 106 30000 136
rect 7606 0 12450 60
<< via3 >>
rect 5952 21614 6016 21618
rect 5952 21558 5956 21614
rect 5956 21558 6012 21614
rect 6012 21558 6016 21614
rect 5952 21554 6016 21558
rect 6032 21614 6096 21618
rect 6032 21558 6036 21614
rect 6036 21558 6092 21614
rect 6092 21558 6096 21614
rect 6032 21554 6096 21558
rect 6112 21614 6176 21618
rect 6112 21558 6116 21614
rect 6116 21558 6172 21614
rect 6172 21558 6176 21614
rect 6112 21554 6176 21558
rect 6192 21614 6256 21618
rect 6192 21558 6196 21614
rect 6196 21558 6252 21614
rect 6252 21558 6256 21614
rect 6192 21554 6256 21558
rect 15952 21614 16016 21618
rect 15952 21558 15956 21614
rect 15956 21558 16012 21614
rect 16012 21558 16016 21614
rect 15952 21554 16016 21558
rect 16032 21614 16096 21618
rect 16032 21558 16036 21614
rect 16036 21558 16092 21614
rect 16092 21558 16096 21614
rect 16032 21554 16096 21558
rect 16112 21614 16176 21618
rect 16112 21558 16116 21614
rect 16116 21558 16172 21614
rect 16172 21558 16176 21614
rect 16112 21554 16176 21558
rect 16192 21614 16256 21618
rect 16192 21558 16196 21614
rect 16196 21558 16252 21614
rect 16252 21558 16256 21614
rect 16192 21554 16256 21558
rect 25952 21614 26016 21618
rect 25952 21558 25956 21614
rect 25956 21558 26012 21614
rect 26012 21558 26016 21614
rect 25952 21554 26016 21558
rect 26032 21614 26096 21618
rect 26032 21558 26036 21614
rect 26036 21558 26092 21614
rect 26092 21558 26096 21614
rect 26032 21554 26096 21558
rect 26112 21614 26176 21618
rect 26112 21558 26116 21614
rect 26116 21558 26172 21614
rect 26172 21558 26176 21614
rect 26112 21554 26176 21558
rect 26192 21614 26256 21618
rect 26192 21558 26196 21614
rect 26196 21558 26252 21614
rect 26252 21558 26256 21614
rect 26192 21554 26256 21558
rect 10952 21070 11016 21074
rect 10952 21014 10956 21070
rect 10956 21014 11012 21070
rect 11012 21014 11016 21070
rect 10952 21010 11016 21014
rect 11032 21070 11096 21074
rect 11032 21014 11036 21070
rect 11036 21014 11092 21070
rect 11092 21014 11096 21070
rect 11032 21010 11096 21014
rect 11112 21070 11176 21074
rect 11112 21014 11116 21070
rect 11116 21014 11172 21070
rect 11172 21014 11176 21070
rect 11112 21010 11176 21014
rect 11192 21070 11256 21074
rect 11192 21014 11196 21070
rect 11196 21014 11252 21070
rect 11252 21014 11256 21070
rect 11192 21010 11256 21014
rect 20952 21070 21016 21074
rect 20952 21014 20956 21070
rect 20956 21014 21012 21070
rect 21012 21014 21016 21070
rect 20952 21010 21016 21014
rect 21032 21070 21096 21074
rect 21032 21014 21036 21070
rect 21036 21014 21092 21070
rect 21092 21014 21096 21070
rect 21032 21010 21096 21014
rect 21112 21070 21176 21074
rect 21112 21014 21116 21070
rect 21116 21014 21172 21070
rect 21172 21014 21176 21070
rect 21112 21010 21176 21014
rect 21192 21070 21256 21074
rect 21192 21014 21196 21070
rect 21196 21014 21252 21070
rect 21252 21014 21256 21070
rect 21192 21010 21256 21014
rect 5952 20526 6016 20530
rect 5952 20470 5956 20526
rect 5956 20470 6012 20526
rect 6012 20470 6016 20526
rect 5952 20466 6016 20470
rect 6032 20526 6096 20530
rect 6032 20470 6036 20526
rect 6036 20470 6092 20526
rect 6092 20470 6096 20526
rect 6032 20466 6096 20470
rect 6112 20526 6176 20530
rect 6112 20470 6116 20526
rect 6116 20470 6172 20526
rect 6172 20470 6176 20526
rect 6112 20466 6176 20470
rect 6192 20526 6256 20530
rect 6192 20470 6196 20526
rect 6196 20470 6252 20526
rect 6252 20470 6256 20526
rect 6192 20466 6256 20470
rect 15952 20526 16016 20530
rect 15952 20470 15956 20526
rect 15956 20470 16012 20526
rect 16012 20470 16016 20526
rect 15952 20466 16016 20470
rect 16032 20526 16096 20530
rect 16032 20470 16036 20526
rect 16036 20470 16092 20526
rect 16092 20470 16096 20526
rect 16032 20466 16096 20470
rect 16112 20526 16176 20530
rect 16112 20470 16116 20526
rect 16116 20470 16172 20526
rect 16172 20470 16176 20526
rect 16112 20466 16176 20470
rect 16192 20526 16256 20530
rect 16192 20470 16196 20526
rect 16196 20470 16252 20526
rect 16252 20470 16256 20526
rect 16192 20466 16256 20470
rect 25952 20526 26016 20530
rect 25952 20470 25956 20526
rect 25956 20470 26012 20526
rect 26012 20470 26016 20526
rect 25952 20466 26016 20470
rect 26032 20526 26096 20530
rect 26032 20470 26036 20526
rect 26036 20470 26092 20526
rect 26092 20470 26096 20526
rect 26032 20466 26096 20470
rect 26112 20526 26176 20530
rect 26112 20470 26116 20526
rect 26116 20470 26172 20526
rect 26172 20470 26176 20526
rect 26112 20466 26176 20470
rect 26192 20526 26256 20530
rect 26192 20470 26196 20526
rect 26196 20470 26252 20526
rect 26252 20470 26256 20526
rect 26192 20466 26256 20470
rect 10952 19982 11016 19986
rect 10952 19926 10956 19982
rect 10956 19926 11012 19982
rect 11012 19926 11016 19982
rect 10952 19922 11016 19926
rect 11032 19982 11096 19986
rect 11032 19926 11036 19982
rect 11036 19926 11092 19982
rect 11092 19926 11096 19982
rect 11032 19922 11096 19926
rect 11112 19982 11176 19986
rect 11112 19926 11116 19982
rect 11116 19926 11172 19982
rect 11172 19926 11176 19982
rect 11112 19922 11176 19926
rect 11192 19982 11256 19986
rect 11192 19926 11196 19982
rect 11196 19926 11252 19982
rect 11252 19926 11256 19982
rect 11192 19922 11256 19926
rect 20952 19982 21016 19986
rect 20952 19926 20956 19982
rect 20956 19926 21012 19982
rect 21012 19926 21016 19982
rect 20952 19922 21016 19926
rect 21032 19982 21096 19986
rect 21032 19926 21036 19982
rect 21036 19926 21092 19982
rect 21092 19926 21096 19982
rect 21032 19922 21096 19926
rect 21112 19982 21176 19986
rect 21112 19926 21116 19982
rect 21116 19926 21172 19982
rect 21172 19926 21176 19982
rect 21112 19922 21176 19926
rect 21192 19982 21256 19986
rect 21192 19926 21196 19982
rect 21196 19926 21252 19982
rect 21252 19926 21256 19982
rect 21192 19922 21256 19926
rect 5952 19438 6016 19442
rect 5952 19382 5956 19438
rect 5956 19382 6012 19438
rect 6012 19382 6016 19438
rect 5952 19378 6016 19382
rect 6032 19438 6096 19442
rect 6032 19382 6036 19438
rect 6036 19382 6092 19438
rect 6092 19382 6096 19438
rect 6032 19378 6096 19382
rect 6112 19438 6176 19442
rect 6112 19382 6116 19438
rect 6116 19382 6172 19438
rect 6172 19382 6176 19438
rect 6112 19378 6176 19382
rect 6192 19438 6256 19442
rect 6192 19382 6196 19438
rect 6196 19382 6252 19438
rect 6252 19382 6256 19438
rect 6192 19378 6256 19382
rect 15952 19438 16016 19442
rect 15952 19382 15956 19438
rect 15956 19382 16012 19438
rect 16012 19382 16016 19438
rect 15952 19378 16016 19382
rect 16032 19438 16096 19442
rect 16032 19382 16036 19438
rect 16036 19382 16092 19438
rect 16092 19382 16096 19438
rect 16032 19378 16096 19382
rect 16112 19438 16176 19442
rect 16112 19382 16116 19438
rect 16116 19382 16172 19438
rect 16172 19382 16176 19438
rect 16112 19378 16176 19382
rect 16192 19438 16256 19442
rect 16192 19382 16196 19438
rect 16196 19382 16252 19438
rect 16252 19382 16256 19438
rect 16192 19378 16256 19382
rect 25952 19438 26016 19442
rect 25952 19382 25956 19438
rect 25956 19382 26012 19438
rect 26012 19382 26016 19438
rect 25952 19378 26016 19382
rect 26032 19438 26096 19442
rect 26032 19382 26036 19438
rect 26036 19382 26092 19438
rect 26092 19382 26096 19438
rect 26032 19378 26096 19382
rect 26112 19438 26176 19442
rect 26112 19382 26116 19438
rect 26116 19382 26172 19438
rect 26172 19382 26176 19438
rect 26112 19378 26176 19382
rect 26192 19438 26256 19442
rect 26192 19382 26196 19438
rect 26196 19382 26252 19438
rect 26252 19382 26256 19438
rect 26192 19378 26256 19382
rect 10952 18894 11016 18898
rect 10952 18838 10956 18894
rect 10956 18838 11012 18894
rect 11012 18838 11016 18894
rect 10952 18834 11016 18838
rect 11032 18894 11096 18898
rect 11032 18838 11036 18894
rect 11036 18838 11092 18894
rect 11092 18838 11096 18894
rect 11032 18834 11096 18838
rect 11112 18894 11176 18898
rect 11112 18838 11116 18894
rect 11116 18838 11172 18894
rect 11172 18838 11176 18894
rect 11112 18834 11176 18838
rect 11192 18894 11256 18898
rect 11192 18838 11196 18894
rect 11196 18838 11252 18894
rect 11252 18838 11256 18894
rect 11192 18834 11256 18838
rect 20952 18894 21016 18898
rect 20952 18838 20956 18894
rect 20956 18838 21012 18894
rect 21012 18838 21016 18894
rect 20952 18834 21016 18838
rect 21032 18894 21096 18898
rect 21032 18838 21036 18894
rect 21036 18838 21092 18894
rect 21092 18838 21096 18894
rect 21032 18834 21096 18838
rect 21112 18894 21176 18898
rect 21112 18838 21116 18894
rect 21116 18838 21172 18894
rect 21172 18838 21176 18894
rect 21112 18834 21176 18838
rect 21192 18894 21256 18898
rect 21192 18838 21196 18894
rect 21196 18838 21252 18894
rect 21252 18838 21256 18894
rect 21192 18834 21256 18838
rect 5952 18350 6016 18354
rect 5952 18294 5956 18350
rect 5956 18294 6012 18350
rect 6012 18294 6016 18350
rect 5952 18290 6016 18294
rect 6032 18350 6096 18354
rect 6032 18294 6036 18350
rect 6036 18294 6092 18350
rect 6092 18294 6096 18350
rect 6032 18290 6096 18294
rect 6112 18350 6176 18354
rect 6112 18294 6116 18350
rect 6116 18294 6172 18350
rect 6172 18294 6176 18350
rect 6112 18290 6176 18294
rect 6192 18350 6256 18354
rect 6192 18294 6196 18350
rect 6196 18294 6252 18350
rect 6252 18294 6256 18350
rect 6192 18290 6256 18294
rect 15952 18350 16016 18354
rect 15952 18294 15956 18350
rect 15956 18294 16012 18350
rect 16012 18294 16016 18350
rect 15952 18290 16016 18294
rect 16032 18350 16096 18354
rect 16032 18294 16036 18350
rect 16036 18294 16092 18350
rect 16092 18294 16096 18350
rect 16032 18290 16096 18294
rect 16112 18350 16176 18354
rect 16112 18294 16116 18350
rect 16116 18294 16172 18350
rect 16172 18294 16176 18350
rect 16112 18290 16176 18294
rect 16192 18350 16256 18354
rect 16192 18294 16196 18350
rect 16196 18294 16252 18350
rect 16252 18294 16256 18350
rect 16192 18290 16256 18294
rect 25952 18350 26016 18354
rect 25952 18294 25956 18350
rect 25956 18294 26012 18350
rect 26012 18294 26016 18350
rect 25952 18290 26016 18294
rect 26032 18350 26096 18354
rect 26032 18294 26036 18350
rect 26036 18294 26092 18350
rect 26092 18294 26096 18350
rect 26032 18290 26096 18294
rect 26112 18350 26176 18354
rect 26112 18294 26116 18350
rect 26116 18294 26172 18350
rect 26172 18294 26176 18350
rect 26112 18290 26176 18294
rect 26192 18350 26256 18354
rect 26192 18294 26196 18350
rect 26196 18294 26252 18350
rect 26252 18294 26256 18350
rect 26192 18290 26256 18294
rect 10952 17806 11016 17810
rect 10952 17750 10956 17806
rect 10956 17750 11012 17806
rect 11012 17750 11016 17806
rect 10952 17746 11016 17750
rect 11032 17806 11096 17810
rect 11032 17750 11036 17806
rect 11036 17750 11092 17806
rect 11092 17750 11096 17806
rect 11032 17746 11096 17750
rect 11112 17806 11176 17810
rect 11112 17750 11116 17806
rect 11116 17750 11172 17806
rect 11172 17750 11176 17806
rect 11112 17746 11176 17750
rect 11192 17806 11256 17810
rect 11192 17750 11196 17806
rect 11196 17750 11252 17806
rect 11252 17750 11256 17806
rect 11192 17746 11256 17750
rect 20952 17806 21016 17810
rect 20952 17750 20956 17806
rect 20956 17750 21012 17806
rect 21012 17750 21016 17806
rect 20952 17746 21016 17750
rect 21032 17806 21096 17810
rect 21032 17750 21036 17806
rect 21036 17750 21092 17806
rect 21092 17750 21096 17806
rect 21032 17746 21096 17750
rect 21112 17806 21176 17810
rect 21112 17750 21116 17806
rect 21116 17750 21172 17806
rect 21172 17750 21176 17806
rect 21112 17746 21176 17750
rect 21192 17806 21256 17810
rect 21192 17750 21196 17806
rect 21196 17750 21252 17806
rect 21252 17750 21256 17806
rect 21192 17746 21256 17750
rect 5952 17262 6016 17266
rect 5952 17206 5956 17262
rect 5956 17206 6012 17262
rect 6012 17206 6016 17262
rect 5952 17202 6016 17206
rect 6032 17262 6096 17266
rect 6032 17206 6036 17262
rect 6036 17206 6092 17262
rect 6092 17206 6096 17262
rect 6032 17202 6096 17206
rect 6112 17262 6176 17266
rect 6112 17206 6116 17262
rect 6116 17206 6172 17262
rect 6172 17206 6176 17262
rect 6112 17202 6176 17206
rect 6192 17262 6256 17266
rect 6192 17206 6196 17262
rect 6196 17206 6252 17262
rect 6252 17206 6256 17262
rect 6192 17202 6256 17206
rect 15952 17262 16016 17266
rect 15952 17206 15956 17262
rect 15956 17206 16012 17262
rect 16012 17206 16016 17262
rect 15952 17202 16016 17206
rect 16032 17262 16096 17266
rect 16032 17206 16036 17262
rect 16036 17206 16092 17262
rect 16092 17206 16096 17262
rect 16032 17202 16096 17206
rect 16112 17262 16176 17266
rect 16112 17206 16116 17262
rect 16116 17206 16172 17262
rect 16172 17206 16176 17262
rect 16112 17202 16176 17206
rect 16192 17262 16256 17266
rect 16192 17206 16196 17262
rect 16196 17206 16252 17262
rect 16252 17206 16256 17262
rect 16192 17202 16256 17206
rect 25952 17262 26016 17266
rect 25952 17206 25956 17262
rect 25956 17206 26012 17262
rect 26012 17206 26016 17262
rect 25952 17202 26016 17206
rect 26032 17262 26096 17266
rect 26032 17206 26036 17262
rect 26036 17206 26092 17262
rect 26092 17206 26096 17262
rect 26032 17202 26096 17206
rect 26112 17262 26176 17266
rect 26112 17206 26116 17262
rect 26116 17206 26172 17262
rect 26172 17206 26176 17262
rect 26112 17202 26176 17206
rect 26192 17262 26256 17266
rect 26192 17206 26196 17262
rect 26196 17206 26252 17262
rect 26252 17206 26256 17262
rect 26192 17202 26256 17206
rect 10952 16718 11016 16722
rect 10952 16662 10956 16718
rect 10956 16662 11012 16718
rect 11012 16662 11016 16718
rect 10952 16658 11016 16662
rect 11032 16718 11096 16722
rect 11032 16662 11036 16718
rect 11036 16662 11092 16718
rect 11092 16662 11096 16718
rect 11032 16658 11096 16662
rect 11112 16718 11176 16722
rect 11112 16662 11116 16718
rect 11116 16662 11172 16718
rect 11172 16662 11176 16718
rect 11112 16658 11176 16662
rect 11192 16718 11256 16722
rect 11192 16662 11196 16718
rect 11196 16662 11252 16718
rect 11252 16662 11256 16718
rect 11192 16658 11256 16662
rect 20952 16718 21016 16722
rect 20952 16662 20956 16718
rect 20956 16662 21012 16718
rect 21012 16662 21016 16718
rect 20952 16658 21016 16662
rect 21032 16718 21096 16722
rect 21032 16662 21036 16718
rect 21036 16662 21092 16718
rect 21092 16662 21096 16718
rect 21032 16658 21096 16662
rect 21112 16718 21176 16722
rect 21112 16662 21116 16718
rect 21116 16662 21172 16718
rect 21172 16662 21176 16718
rect 21112 16658 21176 16662
rect 21192 16718 21256 16722
rect 21192 16662 21196 16718
rect 21196 16662 21252 16718
rect 21252 16662 21256 16718
rect 21192 16658 21256 16662
rect 5952 16174 6016 16178
rect 5952 16118 5956 16174
rect 5956 16118 6012 16174
rect 6012 16118 6016 16174
rect 5952 16114 6016 16118
rect 6032 16174 6096 16178
rect 6032 16118 6036 16174
rect 6036 16118 6092 16174
rect 6092 16118 6096 16174
rect 6032 16114 6096 16118
rect 6112 16174 6176 16178
rect 6112 16118 6116 16174
rect 6116 16118 6172 16174
rect 6172 16118 6176 16174
rect 6112 16114 6176 16118
rect 6192 16174 6256 16178
rect 6192 16118 6196 16174
rect 6196 16118 6252 16174
rect 6252 16118 6256 16174
rect 6192 16114 6256 16118
rect 15952 16174 16016 16178
rect 15952 16118 15956 16174
rect 15956 16118 16012 16174
rect 16012 16118 16016 16174
rect 15952 16114 16016 16118
rect 16032 16174 16096 16178
rect 16032 16118 16036 16174
rect 16036 16118 16092 16174
rect 16092 16118 16096 16174
rect 16032 16114 16096 16118
rect 16112 16174 16176 16178
rect 16112 16118 16116 16174
rect 16116 16118 16172 16174
rect 16172 16118 16176 16174
rect 16112 16114 16176 16118
rect 16192 16174 16256 16178
rect 16192 16118 16196 16174
rect 16196 16118 16252 16174
rect 16252 16118 16256 16174
rect 16192 16114 16256 16118
rect 25952 16174 26016 16178
rect 25952 16118 25956 16174
rect 25956 16118 26012 16174
rect 26012 16118 26016 16174
rect 25952 16114 26016 16118
rect 26032 16174 26096 16178
rect 26032 16118 26036 16174
rect 26036 16118 26092 16174
rect 26092 16118 26096 16174
rect 26032 16114 26096 16118
rect 26112 16174 26176 16178
rect 26112 16118 26116 16174
rect 26116 16118 26172 16174
rect 26172 16118 26176 16174
rect 26112 16114 26176 16118
rect 26192 16174 26256 16178
rect 26192 16118 26196 16174
rect 26196 16118 26252 16174
rect 26252 16118 26256 16174
rect 26192 16114 26256 16118
rect 10952 15630 11016 15634
rect 10952 15574 10956 15630
rect 10956 15574 11012 15630
rect 11012 15574 11016 15630
rect 10952 15570 11016 15574
rect 11032 15630 11096 15634
rect 11032 15574 11036 15630
rect 11036 15574 11092 15630
rect 11092 15574 11096 15630
rect 11032 15570 11096 15574
rect 11112 15630 11176 15634
rect 11112 15574 11116 15630
rect 11116 15574 11172 15630
rect 11172 15574 11176 15630
rect 11112 15570 11176 15574
rect 11192 15630 11256 15634
rect 11192 15574 11196 15630
rect 11196 15574 11252 15630
rect 11252 15574 11256 15630
rect 11192 15570 11256 15574
rect 20952 15630 21016 15634
rect 20952 15574 20956 15630
rect 20956 15574 21012 15630
rect 21012 15574 21016 15630
rect 20952 15570 21016 15574
rect 21032 15630 21096 15634
rect 21032 15574 21036 15630
rect 21036 15574 21092 15630
rect 21092 15574 21096 15630
rect 21032 15570 21096 15574
rect 21112 15630 21176 15634
rect 21112 15574 21116 15630
rect 21116 15574 21172 15630
rect 21172 15574 21176 15630
rect 21112 15570 21176 15574
rect 21192 15630 21256 15634
rect 21192 15574 21196 15630
rect 21196 15574 21252 15630
rect 21252 15574 21256 15630
rect 21192 15570 21256 15574
rect 5952 15086 6016 15090
rect 5952 15030 5956 15086
rect 5956 15030 6012 15086
rect 6012 15030 6016 15086
rect 5952 15026 6016 15030
rect 6032 15086 6096 15090
rect 6032 15030 6036 15086
rect 6036 15030 6092 15086
rect 6092 15030 6096 15086
rect 6032 15026 6096 15030
rect 6112 15086 6176 15090
rect 6112 15030 6116 15086
rect 6116 15030 6172 15086
rect 6172 15030 6176 15086
rect 6112 15026 6176 15030
rect 6192 15086 6256 15090
rect 6192 15030 6196 15086
rect 6196 15030 6252 15086
rect 6252 15030 6256 15086
rect 6192 15026 6256 15030
rect 15952 15086 16016 15090
rect 15952 15030 15956 15086
rect 15956 15030 16012 15086
rect 16012 15030 16016 15086
rect 15952 15026 16016 15030
rect 16032 15086 16096 15090
rect 16032 15030 16036 15086
rect 16036 15030 16092 15086
rect 16092 15030 16096 15086
rect 16032 15026 16096 15030
rect 16112 15086 16176 15090
rect 16112 15030 16116 15086
rect 16116 15030 16172 15086
rect 16172 15030 16176 15086
rect 16112 15026 16176 15030
rect 16192 15086 16256 15090
rect 16192 15030 16196 15086
rect 16196 15030 16252 15086
rect 16252 15030 16256 15086
rect 16192 15026 16256 15030
rect 25952 15086 26016 15090
rect 25952 15030 25956 15086
rect 25956 15030 26012 15086
rect 26012 15030 26016 15086
rect 25952 15026 26016 15030
rect 26032 15086 26096 15090
rect 26032 15030 26036 15086
rect 26036 15030 26092 15086
rect 26092 15030 26096 15086
rect 26032 15026 26096 15030
rect 26112 15086 26176 15090
rect 26112 15030 26116 15086
rect 26116 15030 26172 15086
rect 26172 15030 26176 15086
rect 26112 15026 26176 15030
rect 26192 15086 26256 15090
rect 26192 15030 26196 15086
rect 26196 15030 26252 15086
rect 26252 15030 26256 15086
rect 26192 15026 26256 15030
rect 10952 14542 11016 14546
rect 10952 14486 10956 14542
rect 10956 14486 11012 14542
rect 11012 14486 11016 14542
rect 10952 14482 11016 14486
rect 11032 14542 11096 14546
rect 11032 14486 11036 14542
rect 11036 14486 11092 14542
rect 11092 14486 11096 14542
rect 11032 14482 11096 14486
rect 11112 14542 11176 14546
rect 11112 14486 11116 14542
rect 11116 14486 11172 14542
rect 11172 14486 11176 14542
rect 11112 14482 11176 14486
rect 11192 14542 11256 14546
rect 11192 14486 11196 14542
rect 11196 14486 11252 14542
rect 11252 14486 11256 14542
rect 11192 14482 11256 14486
rect 20952 14542 21016 14546
rect 20952 14486 20956 14542
rect 20956 14486 21012 14542
rect 21012 14486 21016 14542
rect 20952 14482 21016 14486
rect 21032 14542 21096 14546
rect 21032 14486 21036 14542
rect 21036 14486 21092 14542
rect 21092 14486 21096 14542
rect 21032 14482 21096 14486
rect 21112 14542 21176 14546
rect 21112 14486 21116 14542
rect 21116 14486 21172 14542
rect 21172 14486 21176 14542
rect 21112 14482 21176 14486
rect 21192 14542 21256 14546
rect 21192 14486 21196 14542
rect 21196 14486 21252 14542
rect 21252 14486 21256 14542
rect 21192 14482 21256 14486
rect 5952 13998 6016 14002
rect 5952 13942 5956 13998
rect 5956 13942 6012 13998
rect 6012 13942 6016 13998
rect 5952 13938 6016 13942
rect 6032 13998 6096 14002
rect 6032 13942 6036 13998
rect 6036 13942 6092 13998
rect 6092 13942 6096 13998
rect 6032 13938 6096 13942
rect 6112 13998 6176 14002
rect 6112 13942 6116 13998
rect 6116 13942 6172 13998
rect 6172 13942 6176 13998
rect 6112 13938 6176 13942
rect 6192 13998 6256 14002
rect 6192 13942 6196 13998
rect 6196 13942 6252 13998
rect 6252 13942 6256 13998
rect 6192 13938 6256 13942
rect 15952 13998 16016 14002
rect 15952 13942 15956 13998
rect 15956 13942 16012 13998
rect 16012 13942 16016 13998
rect 15952 13938 16016 13942
rect 16032 13998 16096 14002
rect 16032 13942 16036 13998
rect 16036 13942 16092 13998
rect 16092 13942 16096 13998
rect 16032 13938 16096 13942
rect 16112 13998 16176 14002
rect 16112 13942 16116 13998
rect 16116 13942 16172 13998
rect 16172 13942 16176 13998
rect 16112 13938 16176 13942
rect 16192 13998 16256 14002
rect 16192 13942 16196 13998
rect 16196 13942 16252 13998
rect 16252 13942 16256 13998
rect 16192 13938 16256 13942
rect 25952 13998 26016 14002
rect 25952 13942 25956 13998
rect 25956 13942 26012 13998
rect 26012 13942 26016 13998
rect 25952 13938 26016 13942
rect 26032 13998 26096 14002
rect 26032 13942 26036 13998
rect 26036 13942 26092 13998
rect 26092 13942 26096 13998
rect 26032 13938 26096 13942
rect 26112 13998 26176 14002
rect 26112 13942 26116 13998
rect 26116 13942 26172 13998
rect 26172 13942 26176 13998
rect 26112 13938 26176 13942
rect 26192 13998 26256 14002
rect 26192 13942 26196 13998
rect 26196 13942 26252 13998
rect 26252 13942 26256 13998
rect 26192 13938 26256 13942
rect 10952 13454 11016 13458
rect 10952 13398 10956 13454
rect 10956 13398 11012 13454
rect 11012 13398 11016 13454
rect 10952 13394 11016 13398
rect 11032 13454 11096 13458
rect 11032 13398 11036 13454
rect 11036 13398 11092 13454
rect 11092 13398 11096 13454
rect 11032 13394 11096 13398
rect 11112 13454 11176 13458
rect 11112 13398 11116 13454
rect 11116 13398 11172 13454
rect 11172 13398 11176 13454
rect 11112 13394 11176 13398
rect 11192 13454 11256 13458
rect 11192 13398 11196 13454
rect 11196 13398 11252 13454
rect 11252 13398 11256 13454
rect 11192 13394 11256 13398
rect 20952 13454 21016 13458
rect 20952 13398 20956 13454
rect 20956 13398 21012 13454
rect 21012 13398 21016 13454
rect 20952 13394 21016 13398
rect 21032 13454 21096 13458
rect 21032 13398 21036 13454
rect 21036 13398 21092 13454
rect 21092 13398 21096 13454
rect 21032 13394 21096 13398
rect 21112 13454 21176 13458
rect 21112 13398 21116 13454
rect 21116 13398 21172 13454
rect 21172 13398 21176 13454
rect 21112 13394 21176 13398
rect 21192 13454 21256 13458
rect 21192 13398 21196 13454
rect 21196 13398 21252 13454
rect 21252 13398 21256 13454
rect 21192 13394 21256 13398
rect 5952 12910 6016 12914
rect 5952 12854 5956 12910
rect 5956 12854 6012 12910
rect 6012 12854 6016 12910
rect 5952 12850 6016 12854
rect 6032 12910 6096 12914
rect 6032 12854 6036 12910
rect 6036 12854 6092 12910
rect 6092 12854 6096 12910
rect 6032 12850 6096 12854
rect 6112 12910 6176 12914
rect 6112 12854 6116 12910
rect 6116 12854 6172 12910
rect 6172 12854 6176 12910
rect 6112 12850 6176 12854
rect 6192 12910 6256 12914
rect 6192 12854 6196 12910
rect 6196 12854 6252 12910
rect 6252 12854 6256 12910
rect 6192 12850 6256 12854
rect 15952 12910 16016 12914
rect 15952 12854 15956 12910
rect 15956 12854 16012 12910
rect 16012 12854 16016 12910
rect 15952 12850 16016 12854
rect 16032 12910 16096 12914
rect 16032 12854 16036 12910
rect 16036 12854 16092 12910
rect 16092 12854 16096 12910
rect 16032 12850 16096 12854
rect 16112 12910 16176 12914
rect 16112 12854 16116 12910
rect 16116 12854 16172 12910
rect 16172 12854 16176 12910
rect 16112 12850 16176 12854
rect 16192 12910 16256 12914
rect 16192 12854 16196 12910
rect 16196 12854 16252 12910
rect 16252 12854 16256 12910
rect 16192 12850 16256 12854
rect 25952 12910 26016 12914
rect 25952 12854 25956 12910
rect 25956 12854 26012 12910
rect 26012 12854 26016 12910
rect 25952 12850 26016 12854
rect 26032 12910 26096 12914
rect 26032 12854 26036 12910
rect 26036 12854 26092 12910
rect 26092 12854 26096 12910
rect 26032 12850 26096 12854
rect 26112 12910 26176 12914
rect 26112 12854 26116 12910
rect 26116 12854 26172 12910
rect 26172 12854 26176 12910
rect 26112 12850 26176 12854
rect 26192 12910 26256 12914
rect 26192 12854 26196 12910
rect 26196 12854 26252 12910
rect 26252 12854 26256 12910
rect 26192 12850 26256 12854
rect 10952 12366 11016 12370
rect 10952 12310 10956 12366
rect 10956 12310 11012 12366
rect 11012 12310 11016 12366
rect 10952 12306 11016 12310
rect 11032 12366 11096 12370
rect 11032 12310 11036 12366
rect 11036 12310 11092 12366
rect 11092 12310 11096 12366
rect 11032 12306 11096 12310
rect 11112 12366 11176 12370
rect 11112 12310 11116 12366
rect 11116 12310 11172 12366
rect 11172 12310 11176 12366
rect 11112 12306 11176 12310
rect 11192 12366 11256 12370
rect 11192 12310 11196 12366
rect 11196 12310 11252 12366
rect 11252 12310 11256 12366
rect 11192 12306 11256 12310
rect 20952 12366 21016 12370
rect 20952 12310 20956 12366
rect 20956 12310 21012 12366
rect 21012 12310 21016 12366
rect 20952 12306 21016 12310
rect 21032 12366 21096 12370
rect 21032 12310 21036 12366
rect 21036 12310 21092 12366
rect 21092 12310 21096 12366
rect 21032 12306 21096 12310
rect 21112 12366 21176 12370
rect 21112 12310 21116 12366
rect 21116 12310 21172 12366
rect 21172 12310 21176 12366
rect 21112 12306 21176 12310
rect 21192 12366 21256 12370
rect 21192 12310 21196 12366
rect 21196 12310 21252 12366
rect 21252 12310 21256 12366
rect 21192 12306 21256 12310
rect 5952 11822 6016 11826
rect 5952 11766 5956 11822
rect 5956 11766 6012 11822
rect 6012 11766 6016 11822
rect 5952 11762 6016 11766
rect 6032 11822 6096 11826
rect 6032 11766 6036 11822
rect 6036 11766 6092 11822
rect 6092 11766 6096 11822
rect 6032 11762 6096 11766
rect 6112 11822 6176 11826
rect 6112 11766 6116 11822
rect 6116 11766 6172 11822
rect 6172 11766 6176 11822
rect 6112 11762 6176 11766
rect 6192 11822 6256 11826
rect 6192 11766 6196 11822
rect 6196 11766 6252 11822
rect 6252 11766 6256 11822
rect 6192 11762 6256 11766
rect 15952 11822 16016 11826
rect 15952 11766 15956 11822
rect 15956 11766 16012 11822
rect 16012 11766 16016 11822
rect 15952 11762 16016 11766
rect 16032 11822 16096 11826
rect 16032 11766 16036 11822
rect 16036 11766 16092 11822
rect 16092 11766 16096 11822
rect 16032 11762 16096 11766
rect 16112 11822 16176 11826
rect 16112 11766 16116 11822
rect 16116 11766 16172 11822
rect 16172 11766 16176 11822
rect 16112 11762 16176 11766
rect 16192 11822 16256 11826
rect 16192 11766 16196 11822
rect 16196 11766 16252 11822
rect 16252 11766 16256 11822
rect 16192 11762 16256 11766
rect 25952 11822 26016 11826
rect 25952 11766 25956 11822
rect 25956 11766 26012 11822
rect 26012 11766 26016 11822
rect 25952 11762 26016 11766
rect 26032 11822 26096 11826
rect 26032 11766 26036 11822
rect 26036 11766 26092 11822
rect 26092 11766 26096 11822
rect 26032 11762 26096 11766
rect 26112 11822 26176 11826
rect 26112 11766 26116 11822
rect 26116 11766 26172 11822
rect 26172 11766 26176 11822
rect 26112 11762 26176 11766
rect 26192 11822 26256 11826
rect 26192 11766 26196 11822
rect 26196 11766 26252 11822
rect 26252 11766 26256 11822
rect 26192 11762 26256 11766
rect 10952 11278 11016 11282
rect 10952 11222 10956 11278
rect 10956 11222 11012 11278
rect 11012 11222 11016 11278
rect 10952 11218 11016 11222
rect 11032 11278 11096 11282
rect 11032 11222 11036 11278
rect 11036 11222 11092 11278
rect 11092 11222 11096 11278
rect 11032 11218 11096 11222
rect 11112 11278 11176 11282
rect 11112 11222 11116 11278
rect 11116 11222 11172 11278
rect 11172 11222 11176 11278
rect 11112 11218 11176 11222
rect 11192 11278 11256 11282
rect 11192 11222 11196 11278
rect 11196 11222 11252 11278
rect 11252 11222 11256 11278
rect 11192 11218 11256 11222
rect 20952 11278 21016 11282
rect 20952 11222 20956 11278
rect 20956 11222 21012 11278
rect 21012 11222 21016 11278
rect 20952 11218 21016 11222
rect 21032 11278 21096 11282
rect 21032 11222 21036 11278
rect 21036 11222 21092 11278
rect 21092 11222 21096 11278
rect 21032 11218 21096 11222
rect 21112 11278 21176 11282
rect 21112 11222 21116 11278
rect 21116 11222 21172 11278
rect 21172 11222 21176 11278
rect 21112 11218 21176 11222
rect 21192 11278 21256 11282
rect 21192 11222 21196 11278
rect 21196 11222 21252 11278
rect 21252 11222 21256 11278
rect 21192 11218 21256 11222
rect 5952 10734 6016 10738
rect 5952 10678 5956 10734
rect 5956 10678 6012 10734
rect 6012 10678 6016 10734
rect 5952 10674 6016 10678
rect 6032 10734 6096 10738
rect 6032 10678 6036 10734
rect 6036 10678 6092 10734
rect 6092 10678 6096 10734
rect 6032 10674 6096 10678
rect 6112 10734 6176 10738
rect 6112 10678 6116 10734
rect 6116 10678 6172 10734
rect 6172 10678 6176 10734
rect 6112 10674 6176 10678
rect 6192 10734 6256 10738
rect 6192 10678 6196 10734
rect 6196 10678 6252 10734
rect 6252 10678 6256 10734
rect 6192 10674 6256 10678
rect 15952 10734 16016 10738
rect 15952 10678 15956 10734
rect 15956 10678 16012 10734
rect 16012 10678 16016 10734
rect 15952 10674 16016 10678
rect 16032 10734 16096 10738
rect 16032 10678 16036 10734
rect 16036 10678 16092 10734
rect 16092 10678 16096 10734
rect 16032 10674 16096 10678
rect 16112 10734 16176 10738
rect 16112 10678 16116 10734
rect 16116 10678 16172 10734
rect 16172 10678 16176 10734
rect 16112 10674 16176 10678
rect 16192 10734 16256 10738
rect 16192 10678 16196 10734
rect 16196 10678 16252 10734
rect 16252 10678 16256 10734
rect 16192 10674 16256 10678
rect 25952 10734 26016 10738
rect 25952 10678 25956 10734
rect 25956 10678 26012 10734
rect 26012 10678 26016 10734
rect 25952 10674 26016 10678
rect 26032 10734 26096 10738
rect 26032 10678 26036 10734
rect 26036 10678 26092 10734
rect 26092 10678 26096 10734
rect 26032 10674 26096 10678
rect 26112 10734 26176 10738
rect 26112 10678 26116 10734
rect 26116 10678 26172 10734
rect 26172 10678 26176 10734
rect 26112 10674 26176 10678
rect 26192 10734 26256 10738
rect 26192 10678 26196 10734
rect 26196 10678 26252 10734
rect 26252 10678 26256 10734
rect 26192 10674 26256 10678
rect 10952 10190 11016 10194
rect 10952 10134 10956 10190
rect 10956 10134 11012 10190
rect 11012 10134 11016 10190
rect 10952 10130 11016 10134
rect 11032 10190 11096 10194
rect 11032 10134 11036 10190
rect 11036 10134 11092 10190
rect 11092 10134 11096 10190
rect 11032 10130 11096 10134
rect 11112 10190 11176 10194
rect 11112 10134 11116 10190
rect 11116 10134 11172 10190
rect 11172 10134 11176 10190
rect 11112 10130 11176 10134
rect 11192 10190 11256 10194
rect 11192 10134 11196 10190
rect 11196 10134 11252 10190
rect 11252 10134 11256 10190
rect 11192 10130 11256 10134
rect 20952 10190 21016 10194
rect 20952 10134 20956 10190
rect 20956 10134 21012 10190
rect 21012 10134 21016 10190
rect 20952 10130 21016 10134
rect 21032 10190 21096 10194
rect 21032 10134 21036 10190
rect 21036 10134 21092 10190
rect 21092 10134 21096 10190
rect 21032 10130 21096 10134
rect 21112 10190 21176 10194
rect 21112 10134 21116 10190
rect 21116 10134 21172 10190
rect 21172 10134 21176 10190
rect 21112 10130 21176 10134
rect 21192 10190 21256 10194
rect 21192 10134 21196 10190
rect 21196 10134 21252 10190
rect 21252 10134 21256 10190
rect 21192 10130 21256 10134
rect 5952 9646 6016 9650
rect 5952 9590 5956 9646
rect 5956 9590 6012 9646
rect 6012 9590 6016 9646
rect 5952 9586 6016 9590
rect 6032 9646 6096 9650
rect 6032 9590 6036 9646
rect 6036 9590 6092 9646
rect 6092 9590 6096 9646
rect 6032 9586 6096 9590
rect 6112 9646 6176 9650
rect 6112 9590 6116 9646
rect 6116 9590 6172 9646
rect 6172 9590 6176 9646
rect 6112 9586 6176 9590
rect 6192 9646 6256 9650
rect 6192 9590 6196 9646
rect 6196 9590 6252 9646
rect 6252 9590 6256 9646
rect 6192 9586 6256 9590
rect 15952 9646 16016 9650
rect 15952 9590 15956 9646
rect 15956 9590 16012 9646
rect 16012 9590 16016 9646
rect 15952 9586 16016 9590
rect 16032 9646 16096 9650
rect 16032 9590 16036 9646
rect 16036 9590 16092 9646
rect 16092 9590 16096 9646
rect 16032 9586 16096 9590
rect 16112 9646 16176 9650
rect 16112 9590 16116 9646
rect 16116 9590 16172 9646
rect 16172 9590 16176 9646
rect 16112 9586 16176 9590
rect 16192 9646 16256 9650
rect 16192 9590 16196 9646
rect 16196 9590 16252 9646
rect 16252 9590 16256 9646
rect 16192 9586 16256 9590
rect 25952 9646 26016 9650
rect 25952 9590 25956 9646
rect 25956 9590 26012 9646
rect 26012 9590 26016 9646
rect 25952 9586 26016 9590
rect 26032 9646 26096 9650
rect 26032 9590 26036 9646
rect 26036 9590 26092 9646
rect 26092 9590 26096 9646
rect 26032 9586 26096 9590
rect 26112 9646 26176 9650
rect 26112 9590 26116 9646
rect 26116 9590 26172 9646
rect 26172 9590 26176 9646
rect 26112 9586 26176 9590
rect 26192 9646 26256 9650
rect 26192 9590 26196 9646
rect 26196 9590 26252 9646
rect 26252 9590 26256 9646
rect 26192 9586 26256 9590
rect 10952 9102 11016 9106
rect 10952 9046 10956 9102
rect 10956 9046 11012 9102
rect 11012 9046 11016 9102
rect 10952 9042 11016 9046
rect 11032 9102 11096 9106
rect 11032 9046 11036 9102
rect 11036 9046 11092 9102
rect 11092 9046 11096 9102
rect 11032 9042 11096 9046
rect 11112 9102 11176 9106
rect 11112 9046 11116 9102
rect 11116 9046 11172 9102
rect 11172 9046 11176 9102
rect 11112 9042 11176 9046
rect 11192 9102 11256 9106
rect 11192 9046 11196 9102
rect 11196 9046 11252 9102
rect 11252 9046 11256 9102
rect 11192 9042 11256 9046
rect 20952 9102 21016 9106
rect 20952 9046 20956 9102
rect 20956 9046 21012 9102
rect 21012 9046 21016 9102
rect 20952 9042 21016 9046
rect 21032 9102 21096 9106
rect 21032 9046 21036 9102
rect 21036 9046 21092 9102
rect 21092 9046 21096 9102
rect 21032 9042 21096 9046
rect 21112 9102 21176 9106
rect 21112 9046 21116 9102
rect 21116 9046 21172 9102
rect 21172 9046 21176 9102
rect 21112 9042 21176 9046
rect 21192 9102 21256 9106
rect 21192 9046 21196 9102
rect 21196 9046 21252 9102
rect 21252 9046 21256 9102
rect 21192 9042 21256 9046
rect 5952 8558 6016 8562
rect 5952 8502 5956 8558
rect 5956 8502 6012 8558
rect 6012 8502 6016 8558
rect 5952 8498 6016 8502
rect 6032 8558 6096 8562
rect 6032 8502 6036 8558
rect 6036 8502 6092 8558
rect 6092 8502 6096 8558
rect 6032 8498 6096 8502
rect 6112 8558 6176 8562
rect 6112 8502 6116 8558
rect 6116 8502 6172 8558
rect 6172 8502 6176 8558
rect 6112 8498 6176 8502
rect 6192 8558 6256 8562
rect 6192 8502 6196 8558
rect 6196 8502 6252 8558
rect 6252 8502 6256 8558
rect 6192 8498 6256 8502
rect 15952 8558 16016 8562
rect 15952 8502 15956 8558
rect 15956 8502 16012 8558
rect 16012 8502 16016 8558
rect 15952 8498 16016 8502
rect 16032 8558 16096 8562
rect 16032 8502 16036 8558
rect 16036 8502 16092 8558
rect 16092 8502 16096 8558
rect 16032 8498 16096 8502
rect 16112 8558 16176 8562
rect 16112 8502 16116 8558
rect 16116 8502 16172 8558
rect 16172 8502 16176 8558
rect 16112 8498 16176 8502
rect 16192 8558 16256 8562
rect 16192 8502 16196 8558
rect 16196 8502 16252 8558
rect 16252 8502 16256 8558
rect 16192 8498 16256 8502
rect 25952 8558 26016 8562
rect 25952 8502 25956 8558
rect 25956 8502 26012 8558
rect 26012 8502 26016 8558
rect 25952 8498 26016 8502
rect 26032 8558 26096 8562
rect 26032 8502 26036 8558
rect 26036 8502 26092 8558
rect 26092 8502 26096 8558
rect 26032 8498 26096 8502
rect 26112 8558 26176 8562
rect 26112 8502 26116 8558
rect 26116 8502 26172 8558
rect 26172 8502 26176 8558
rect 26112 8498 26176 8502
rect 26192 8558 26256 8562
rect 26192 8502 26196 8558
rect 26196 8502 26252 8558
rect 26252 8502 26256 8558
rect 26192 8498 26256 8502
rect 10952 8014 11016 8018
rect 10952 7958 10956 8014
rect 10956 7958 11012 8014
rect 11012 7958 11016 8014
rect 10952 7954 11016 7958
rect 11032 8014 11096 8018
rect 11032 7958 11036 8014
rect 11036 7958 11092 8014
rect 11092 7958 11096 8014
rect 11032 7954 11096 7958
rect 11112 8014 11176 8018
rect 11112 7958 11116 8014
rect 11116 7958 11172 8014
rect 11172 7958 11176 8014
rect 11112 7954 11176 7958
rect 11192 8014 11256 8018
rect 11192 7958 11196 8014
rect 11196 7958 11252 8014
rect 11252 7958 11256 8014
rect 11192 7954 11256 7958
rect 20952 8014 21016 8018
rect 20952 7958 20956 8014
rect 20956 7958 21012 8014
rect 21012 7958 21016 8014
rect 20952 7954 21016 7958
rect 21032 8014 21096 8018
rect 21032 7958 21036 8014
rect 21036 7958 21092 8014
rect 21092 7958 21096 8014
rect 21032 7954 21096 7958
rect 21112 8014 21176 8018
rect 21112 7958 21116 8014
rect 21116 7958 21172 8014
rect 21172 7958 21176 8014
rect 21112 7954 21176 7958
rect 21192 8014 21256 8018
rect 21192 7958 21196 8014
rect 21196 7958 21252 8014
rect 21252 7958 21256 8014
rect 21192 7954 21256 7958
rect 5952 7470 6016 7474
rect 5952 7414 5956 7470
rect 5956 7414 6012 7470
rect 6012 7414 6016 7470
rect 5952 7410 6016 7414
rect 6032 7470 6096 7474
rect 6032 7414 6036 7470
rect 6036 7414 6092 7470
rect 6092 7414 6096 7470
rect 6032 7410 6096 7414
rect 6112 7470 6176 7474
rect 6112 7414 6116 7470
rect 6116 7414 6172 7470
rect 6172 7414 6176 7470
rect 6112 7410 6176 7414
rect 6192 7470 6256 7474
rect 6192 7414 6196 7470
rect 6196 7414 6252 7470
rect 6252 7414 6256 7470
rect 6192 7410 6256 7414
rect 15952 7470 16016 7474
rect 15952 7414 15956 7470
rect 15956 7414 16012 7470
rect 16012 7414 16016 7470
rect 15952 7410 16016 7414
rect 16032 7470 16096 7474
rect 16032 7414 16036 7470
rect 16036 7414 16092 7470
rect 16092 7414 16096 7470
rect 16032 7410 16096 7414
rect 16112 7470 16176 7474
rect 16112 7414 16116 7470
rect 16116 7414 16172 7470
rect 16172 7414 16176 7470
rect 16112 7410 16176 7414
rect 16192 7470 16256 7474
rect 16192 7414 16196 7470
rect 16196 7414 16252 7470
rect 16252 7414 16256 7470
rect 16192 7410 16256 7414
rect 25952 7470 26016 7474
rect 25952 7414 25956 7470
rect 25956 7414 26012 7470
rect 26012 7414 26016 7470
rect 25952 7410 26016 7414
rect 26032 7470 26096 7474
rect 26032 7414 26036 7470
rect 26036 7414 26092 7470
rect 26092 7414 26096 7470
rect 26032 7410 26096 7414
rect 26112 7470 26176 7474
rect 26112 7414 26116 7470
rect 26116 7414 26172 7470
rect 26172 7414 26176 7470
rect 26112 7410 26176 7414
rect 26192 7470 26256 7474
rect 26192 7414 26196 7470
rect 26196 7414 26252 7470
rect 26252 7414 26256 7470
rect 26192 7410 26256 7414
rect 10952 6926 11016 6930
rect 10952 6870 10956 6926
rect 10956 6870 11012 6926
rect 11012 6870 11016 6926
rect 10952 6866 11016 6870
rect 11032 6926 11096 6930
rect 11032 6870 11036 6926
rect 11036 6870 11092 6926
rect 11092 6870 11096 6926
rect 11032 6866 11096 6870
rect 11112 6926 11176 6930
rect 11112 6870 11116 6926
rect 11116 6870 11172 6926
rect 11172 6870 11176 6926
rect 11112 6866 11176 6870
rect 11192 6926 11256 6930
rect 11192 6870 11196 6926
rect 11196 6870 11252 6926
rect 11252 6870 11256 6926
rect 11192 6866 11256 6870
rect 20952 6926 21016 6930
rect 20952 6870 20956 6926
rect 20956 6870 21012 6926
rect 21012 6870 21016 6926
rect 20952 6866 21016 6870
rect 21032 6926 21096 6930
rect 21032 6870 21036 6926
rect 21036 6870 21092 6926
rect 21092 6870 21096 6926
rect 21032 6866 21096 6870
rect 21112 6926 21176 6930
rect 21112 6870 21116 6926
rect 21116 6870 21172 6926
rect 21172 6870 21176 6926
rect 21112 6866 21176 6870
rect 21192 6926 21256 6930
rect 21192 6870 21196 6926
rect 21196 6870 21252 6926
rect 21252 6870 21256 6926
rect 21192 6866 21256 6870
rect 5952 6382 6016 6386
rect 5952 6326 5956 6382
rect 5956 6326 6012 6382
rect 6012 6326 6016 6382
rect 5952 6322 6016 6326
rect 6032 6382 6096 6386
rect 6032 6326 6036 6382
rect 6036 6326 6092 6382
rect 6092 6326 6096 6382
rect 6032 6322 6096 6326
rect 6112 6382 6176 6386
rect 6112 6326 6116 6382
rect 6116 6326 6172 6382
rect 6172 6326 6176 6382
rect 6112 6322 6176 6326
rect 6192 6382 6256 6386
rect 6192 6326 6196 6382
rect 6196 6326 6252 6382
rect 6252 6326 6256 6382
rect 6192 6322 6256 6326
rect 15952 6382 16016 6386
rect 15952 6326 15956 6382
rect 15956 6326 16012 6382
rect 16012 6326 16016 6382
rect 15952 6322 16016 6326
rect 16032 6382 16096 6386
rect 16032 6326 16036 6382
rect 16036 6326 16092 6382
rect 16092 6326 16096 6382
rect 16032 6322 16096 6326
rect 16112 6382 16176 6386
rect 16112 6326 16116 6382
rect 16116 6326 16172 6382
rect 16172 6326 16176 6382
rect 16112 6322 16176 6326
rect 16192 6382 16256 6386
rect 16192 6326 16196 6382
rect 16196 6326 16252 6382
rect 16252 6326 16256 6382
rect 16192 6322 16256 6326
rect 25952 6382 26016 6386
rect 25952 6326 25956 6382
rect 25956 6326 26012 6382
rect 26012 6326 26016 6382
rect 25952 6322 26016 6326
rect 26032 6382 26096 6386
rect 26032 6326 26036 6382
rect 26036 6326 26092 6382
rect 26092 6326 26096 6382
rect 26032 6322 26096 6326
rect 26112 6382 26176 6386
rect 26112 6326 26116 6382
rect 26116 6326 26172 6382
rect 26172 6326 26176 6382
rect 26112 6322 26176 6326
rect 26192 6382 26256 6386
rect 26192 6326 26196 6382
rect 26196 6326 26252 6382
rect 26252 6326 26256 6382
rect 26192 6322 26256 6326
rect 10952 5838 11016 5842
rect 10952 5782 10956 5838
rect 10956 5782 11012 5838
rect 11012 5782 11016 5838
rect 10952 5778 11016 5782
rect 11032 5838 11096 5842
rect 11032 5782 11036 5838
rect 11036 5782 11092 5838
rect 11092 5782 11096 5838
rect 11032 5778 11096 5782
rect 11112 5838 11176 5842
rect 11112 5782 11116 5838
rect 11116 5782 11172 5838
rect 11172 5782 11176 5838
rect 11112 5778 11176 5782
rect 11192 5838 11256 5842
rect 11192 5782 11196 5838
rect 11196 5782 11252 5838
rect 11252 5782 11256 5838
rect 11192 5778 11256 5782
rect 20952 5838 21016 5842
rect 20952 5782 20956 5838
rect 20956 5782 21012 5838
rect 21012 5782 21016 5838
rect 20952 5778 21016 5782
rect 21032 5838 21096 5842
rect 21032 5782 21036 5838
rect 21036 5782 21092 5838
rect 21092 5782 21096 5838
rect 21032 5778 21096 5782
rect 21112 5838 21176 5842
rect 21112 5782 21116 5838
rect 21116 5782 21172 5838
rect 21172 5782 21176 5838
rect 21112 5778 21176 5782
rect 21192 5838 21256 5842
rect 21192 5782 21196 5838
rect 21196 5782 21252 5838
rect 21252 5782 21256 5838
rect 21192 5778 21256 5782
rect 5952 5294 6016 5298
rect 5952 5238 5956 5294
rect 5956 5238 6012 5294
rect 6012 5238 6016 5294
rect 5952 5234 6016 5238
rect 6032 5294 6096 5298
rect 6032 5238 6036 5294
rect 6036 5238 6092 5294
rect 6092 5238 6096 5294
rect 6032 5234 6096 5238
rect 6112 5294 6176 5298
rect 6112 5238 6116 5294
rect 6116 5238 6172 5294
rect 6172 5238 6176 5294
rect 6112 5234 6176 5238
rect 6192 5294 6256 5298
rect 6192 5238 6196 5294
rect 6196 5238 6252 5294
rect 6252 5238 6256 5294
rect 6192 5234 6256 5238
rect 15952 5294 16016 5298
rect 15952 5238 15956 5294
rect 15956 5238 16012 5294
rect 16012 5238 16016 5294
rect 15952 5234 16016 5238
rect 16032 5294 16096 5298
rect 16032 5238 16036 5294
rect 16036 5238 16092 5294
rect 16092 5238 16096 5294
rect 16032 5234 16096 5238
rect 16112 5294 16176 5298
rect 16112 5238 16116 5294
rect 16116 5238 16172 5294
rect 16172 5238 16176 5294
rect 16112 5234 16176 5238
rect 16192 5294 16256 5298
rect 16192 5238 16196 5294
rect 16196 5238 16252 5294
rect 16252 5238 16256 5294
rect 16192 5234 16256 5238
rect 25952 5294 26016 5298
rect 25952 5238 25956 5294
rect 25956 5238 26012 5294
rect 26012 5238 26016 5294
rect 25952 5234 26016 5238
rect 26032 5294 26096 5298
rect 26032 5238 26036 5294
rect 26036 5238 26092 5294
rect 26092 5238 26096 5294
rect 26032 5234 26096 5238
rect 26112 5294 26176 5298
rect 26112 5238 26116 5294
rect 26116 5238 26172 5294
rect 26172 5238 26176 5294
rect 26112 5234 26176 5238
rect 26192 5294 26256 5298
rect 26192 5238 26196 5294
rect 26196 5238 26252 5294
rect 26252 5238 26256 5294
rect 26192 5234 26256 5238
rect 10952 4750 11016 4754
rect 10952 4694 10956 4750
rect 10956 4694 11012 4750
rect 11012 4694 11016 4750
rect 10952 4690 11016 4694
rect 11032 4750 11096 4754
rect 11032 4694 11036 4750
rect 11036 4694 11092 4750
rect 11092 4694 11096 4750
rect 11032 4690 11096 4694
rect 11112 4750 11176 4754
rect 11112 4694 11116 4750
rect 11116 4694 11172 4750
rect 11172 4694 11176 4750
rect 11112 4690 11176 4694
rect 11192 4750 11256 4754
rect 11192 4694 11196 4750
rect 11196 4694 11252 4750
rect 11252 4694 11256 4750
rect 11192 4690 11256 4694
rect 20952 4750 21016 4754
rect 20952 4694 20956 4750
rect 20956 4694 21012 4750
rect 21012 4694 21016 4750
rect 20952 4690 21016 4694
rect 21032 4750 21096 4754
rect 21032 4694 21036 4750
rect 21036 4694 21092 4750
rect 21092 4694 21096 4750
rect 21032 4690 21096 4694
rect 21112 4750 21176 4754
rect 21112 4694 21116 4750
rect 21116 4694 21172 4750
rect 21172 4694 21176 4750
rect 21112 4690 21176 4694
rect 21192 4750 21256 4754
rect 21192 4694 21196 4750
rect 21196 4694 21252 4750
rect 21252 4694 21256 4750
rect 21192 4690 21256 4694
rect 5952 4206 6016 4210
rect 5952 4150 5956 4206
rect 5956 4150 6012 4206
rect 6012 4150 6016 4206
rect 5952 4146 6016 4150
rect 6032 4206 6096 4210
rect 6032 4150 6036 4206
rect 6036 4150 6092 4206
rect 6092 4150 6096 4206
rect 6032 4146 6096 4150
rect 6112 4206 6176 4210
rect 6112 4150 6116 4206
rect 6116 4150 6172 4206
rect 6172 4150 6176 4206
rect 6112 4146 6176 4150
rect 6192 4206 6256 4210
rect 6192 4150 6196 4206
rect 6196 4150 6252 4206
rect 6252 4150 6256 4206
rect 6192 4146 6256 4150
rect 15952 4206 16016 4210
rect 15952 4150 15956 4206
rect 15956 4150 16012 4206
rect 16012 4150 16016 4206
rect 15952 4146 16016 4150
rect 16032 4206 16096 4210
rect 16032 4150 16036 4206
rect 16036 4150 16092 4206
rect 16092 4150 16096 4206
rect 16032 4146 16096 4150
rect 16112 4206 16176 4210
rect 16112 4150 16116 4206
rect 16116 4150 16172 4206
rect 16172 4150 16176 4206
rect 16112 4146 16176 4150
rect 16192 4206 16256 4210
rect 16192 4150 16196 4206
rect 16196 4150 16252 4206
rect 16252 4150 16256 4206
rect 16192 4146 16256 4150
rect 25952 4206 26016 4210
rect 25952 4150 25956 4206
rect 25956 4150 26012 4206
rect 26012 4150 26016 4206
rect 25952 4146 26016 4150
rect 26032 4206 26096 4210
rect 26032 4150 26036 4206
rect 26036 4150 26092 4206
rect 26092 4150 26096 4206
rect 26032 4146 26096 4150
rect 26112 4206 26176 4210
rect 26112 4150 26116 4206
rect 26116 4150 26172 4206
rect 26172 4150 26176 4206
rect 26112 4146 26176 4150
rect 26192 4206 26256 4210
rect 26192 4150 26196 4206
rect 26196 4150 26252 4206
rect 26252 4150 26256 4206
rect 26192 4146 26256 4150
rect 10952 3662 11016 3666
rect 10952 3606 10956 3662
rect 10956 3606 11012 3662
rect 11012 3606 11016 3662
rect 10952 3602 11016 3606
rect 11032 3662 11096 3666
rect 11032 3606 11036 3662
rect 11036 3606 11092 3662
rect 11092 3606 11096 3662
rect 11032 3602 11096 3606
rect 11112 3662 11176 3666
rect 11112 3606 11116 3662
rect 11116 3606 11172 3662
rect 11172 3606 11176 3662
rect 11112 3602 11176 3606
rect 11192 3662 11256 3666
rect 11192 3606 11196 3662
rect 11196 3606 11252 3662
rect 11252 3606 11256 3662
rect 11192 3602 11256 3606
rect 20952 3662 21016 3666
rect 20952 3606 20956 3662
rect 20956 3606 21012 3662
rect 21012 3606 21016 3662
rect 20952 3602 21016 3606
rect 21032 3662 21096 3666
rect 21032 3606 21036 3662
rect 21036 3606 21092 3662
rect 21092 3606 21096 3662
rect 21032 3602 21096 3606
rect 21112 3662 21176 3666
rect 21112 3606 21116 3662
rect 21116 3606 21172 3662
rect 21172 3606 21176 3662
rect 21112 3602 21176 3606
rect 21192 3662 21256 3666
rect 21192 3606 21196 3662
rect 21196 3606 21252 3662
rect 21252 3606 21256 3662
rect 21192 3602 21256 3606
rect 5952 3118 6016 3122
rect 5952 3062 5956 3118
rect 5956 3062 6012 3118
rect 6012 3062 6016 3118
rect 5952 3058 6016 3062
rect 6032 3118 6096 3122
rect 6032 3062 6036 3118
rect 6036 3062 6092 3118
rect 6092 3062 6096 3118
rect 6032 3058 6096 3062
rect 6112 3118 6176 3122
rect 6112 3062 6116 3118
rect 6116 3062 6172 3118
rect 6172 3062 6176 3118
rect 6112 3058 6176 3062
rect 6192 3118 6256 3122
rect 6192 3062 6196 3118
rect 6196 3062 6252 3118
rect 6252 3062 6256 3118
rect 6192 3058 6256 3062
rect 15952 3118 16016 3122
rect 15952 3062 15956 3118
rect 15956 3062 16012 3118
rect 16012 3062 16016 3118
rect 15952 3058 16016 3062
rect 16032 3118 16096 3122
rect 16032 3062 16036 3118
rect 16036 3062 16092 3118
rect 16092 3062 16096 3118
rect 16032 3058 16096 3062
rect 16112 3118 16176 3122
rect 16112 3062 16116 3118
rect 16116 3062 16172 3118
rect 16172 3062 16176 3118
rect 16112 3058 16176 3062
rect 16192 3118 16256 3122
rect 16192 3062 16196 3118
rect 16196 3062 16252 3118
rect 16252 3062 16256 3118
rect 16192 3058 16256 3062
rect 25952 3118 26016 3122
rect 25952 3062 25956 3118
rect 25956 3062 26012 3118
rect 26012 3062 26016 3118
rect 25952 3058 26016 3062
rect 26032 3118 26096 3122
rect 26032 3062 26036 3118
rect 26036 3062 26092 3118
rect 26092 3062 26096 3118
rect 26032 3058 26096 3062
rect 26112 3118 26176 3122
rect 26112 3062 26116 3118
rect 26116 3062 26172 3118
rect 26172 3062 26176 3118
rect 26112 3058 26176 3062
rect 26192 3118 26256 3122
rect 26192 3062 26196 3118
rect 26196 3062 26252 3118
rect 26252 3062 26256 3118
rect 26192 3058 26256 3062
rect 10952 2574 11016 2578
rect 10952 2518 10956 2574
rect 10956 2518 11012 2574
rect 11012 2518 11016 2574
rect 10952 2514 11016 2518
rect 11032 2574 11096 2578
rect 11032 2518 11036 2574
rect 11036 2518 11092 2574
rect 11092 2518 11096 2574
rect 11032 2514 11096 2518
rect 11112 2574 11176 2578
rect 11112 2518 11116 2574
rect 11116 2518 11172 2574
rect 11172 2518 11176 2574
rect 11112 2514 11176 2518
rect 11192 2574 11256 2578
rect 11192 2518 11196 2574
rect 11196 2518 11252 2574
rect 11252 2518 11256 2574
rect 11192 2514 11256 2518
rect 20952 2574 21016 2578
rect 20952 2518 20956 2574
rect 20956 2518 21012 2574
rect 21012 2518 21016 2574
rect 20952 2514 21016 2518
rect 21032 2574 21096 2578
rect 21032 2518 21036 2574
rect 21036 2518 21092 2574
rect 21092 2518 21096 2574
rect 21032 2514 21096 2518
rect 21112 2574 21176 2578
rect 21112 2518 21116 2574
rect 21116 2518 21172 2574
rect 21172 2518 21176 2574
rect 21112 2514 21176 2518
rect 21192 2574 21256 2578
rect 21192 2518 21196 2574
rect 21196 2518 21252 2574
rect 21252 2518 21256 2574
rect 21192 2514 21256 2518
rect 5952 2030 6016 2034
rect 5952 1974 5956 2030
rect 5956 1974 6012 2030
rect 6012 1974 6016 2030
rect 5952 1970 6016 1974
rect 6032 2030 6096 2034
rect 6032 1974 6036 2030
rect 6036 1974 6092 2030
rect 6092 1974 6096 2030
rect 6032 1970 6096 1974
rect 6112 2030 6176 2034
rect 6112 1974 6116 2030
rect 6116 1974 6172 2030
rect 6172 1974 6176 2030
rect 6112 1970 6176 1974
rect 6192 2030 6256 2034
rect 6192 1974 6196 2030
rect 6196 1974 6252 2030
rect 6252 1974 6256 2030
rect 6192 1970 6256 1974
rect 15952 2030 16016 2034
rect 15952 1974 15956 2030
rect 15956 1974 16012 2030
rect 16012 1974 16016 2030
rect 15952 1970 16016 1974
rect 16032 2030 16096 2034
rect 16032 1974 16036 2030
rect 16036 1974 16092 2030
rect 16092 1974 16096 2030
rect 16032 1970 16096 1974
rect 16112 2030 16176 2034
rect 16112 1974 16116 2030
rect 16116 1974 16172 2030
rect 16172 1974 16176 2030
rect 16112 1970 16176 1974
rect 16192 2030 16256 2034
rect 16192 1974 16196 2030
rect 16196 1974 16252 2030
rect 16252 1974 16256 2030
rect 16192 1970 16256 1974
rect 25952 2030 26016 2034
rect 25952 1974 25956 2030
rect 25956 1974 26012 2030
rect 26012 1974 26016 2030
rect 25952 1970 26016 1974
rect 26032 2030 26096 2034
rect 26032 1974 26036 2030
rect 26036 1974 26092 2030
rect 26092 1974 26096 2030
rect 26032 1970 26096 1974
rect 26112 2030 26176 2034
rect 26112 1974 26116 2030
rect 26116 1974 26172 2030
rect 26172 1974 26176 2030
rect 26112 1970 26176 1974
rect 26192 2030 26256 2034
rect 26192 1974 26196 2030
rect 26196 1974 26252 2030
rect 26252 1974 26256 2030
rect 26192 1970 26256 1974
<< metal4 >>
rect 5944 21618 6264 21634
rect 5944 21554 5952 21618
rect 6016 21554 6032 21618
rect 6096 21554 6112 21618
rect 6176 21554 6192 21618
rect 6256 21554 6264 21618
rect 5944 20530 6264 21554
rect 5944 20466 5952 20530
rect 6016 20466 6032 20530
rect 6096 20466 6112 20530
rect 6176 20466 6192 20530
rect 6256 20466 6264 20530
rect 5944 19442 6264 20466
rect 5944 19378 5952 19442
rect 6016 19378 6032 19442
rect 6096 19378 6112 19442
rect 6176 19378 6192 19442
rect 6256 19378 6264 19442
rect 5944 18354 6264 19378
rect 5944 18290 5952 18354
rect 6016 18290 6032 18354
rect 6096 18290 6112 18354
rect 6176 18290 6192 18354
rect 6256 18290 6264 18354
rect 5944 17266 6264 18290
rect 5944 17202 5952 17266
rect 6016 17202 6032 17266
rect 6096 17202 6112 17266
rect 6176 17202 6192 17266
rect 6256 17202 6264 17266
rect 5944 16178 6264 17202
rect 5944 16114 5952 16178
rect 6016 16114 6032 16178
rect 6096 16114 6112 16178
rect 6176 16114 6192 16178
rect 6256 16114 6264 16178
rect 5944 15090 6264 16114
rect 5944 15026 5952 15090
rect 6016 15026 6032 15090
rect 6096 15026 6112 15090
rect 6176 15026 6192 15090
rect 6256 15026 6264 15090
rect 5944 14002 6264 15026
rect 5944 13938 5952 14002
rect 6016 13938 6032 14002
rect 6096 13938 6112 14002
rect 6176 13938 6192 14002
rect 6256 13938 6264 14002
rect 5944 12914 6264 13938
rect 5944 12850 5952 12914
rect 6016 12850 6032 12914
rect 6096 12850 6112 12914
rect 6176 12850 6192 12914
rect 6256 12850 6264 12914
rect 5944 11826 6264 12850
rect 5944 11762 5952 11826
rect 6016 11762 6032 11826
rect 6096 11762 6112 11826
rect 6176 11762 6192 11826
rect 6256 11762 6264 11826
rect 5944 10738 6264 11762
rect 5944 10674 5952 10738
rect 6016 10674 6032 10738
rect 6096 10674 6112 10738
rect 6176 10674 6192 10738
rect 6256 10674 6264 10738
rect 5944 9650 6264 10674
rect 5944 9586 5952 9650
rect 6016 9586 6032 9650
rect 6096 9586 6112 9650
rect 6176 9586 6192 9650
rect 6256 9586 6264 9650
rect 5944 8562 6264 9586
rect 5944 8498 5952 8562
rect 6016 8498 6032 8562
rect 6096 8498 6112 8562
rect 6176 8498 6192 8562
rect 6256 8498 6264 8562
rect 5944 7474 6264 8498
rect 5944 7410 5952 7474
rect 6016 7410 6032 7474
rect 6096 7410 6112 7474
rect 6176 7410 6192 7474
rect 6256 7410 6264 7474
rect 5944 6386 6264 7410
rect 5944 6322 5952 6386
rect 6016 6322 6032 6386
rect 6096 6322 6112 6386
rect 6176 6322 6192 6386
rect 6256 6322 6264 6386
rect 5944 5298 6264 6322
rect 5944 5234 5952 5298
rect 6016 5234 6032 5298
rect 6096 5234 6112 5298
rect 6176 5234 6192 5298
rect 6256 5234 6264 5298
rect 5944 4210 6264 5234
rect 5944 4146 5952 4210
rect 6016 4146 6032 4210
rect 6096 4146 6112 4210
rect 6176 4146 6192 4210
rect 6256 4146 6264 4210
rect 5944 3122 6264 4146
rect 5944 3058 5952 3122
rect 6016 3058 6032 3122
rect 6096 3058 6112 3122
rect 6176 3058 6192 3122
rect 6256 3058 6264 3122
rect 5944 2034 6264 3058
rect 5944 1970 5952 2034
rect 6016 1970 6032 2034
rect 6096 1970 6112 2034
rect 6176 1970 6192 2034
rect 6256 1970 6264 2034
rect 5944 1954 6264 1970
rect 10944 21074 11264 21634
rect 10944 21010 10952 21074
rect 11016 21010 11032 21074
rect 11096 21010 11112 21074
rect 11176 21010 11192 21074
rect 11256 21010 11264 21074
rect 10944 19986 11264 21010
rect 10944 19922 10952 19986
rect 11016 19922 11032 19986
rect 11096 19922 11112 19986
rect 11176 19922 11192 19986
rect 11256 19922 11264 19986
rect 10944 18898 11264 19922
rect 10944 18834 10952 18898
rect 11016 18834 11032 18898
rect 11096 18834 11112 18898
rect 11176 18834 11192 18898
rect 11256 18834 11264 18898
rect 10944 17810 11264 18834
rect 10944 17746 10952 17810
rect 11016 17746 11032 17810
rect 11096 17746 11112 17810
rect 11176 17746 11192 17810
rect 11256 17746 11264 17810
rect 10944 16722 11264 17746
rect 10944 16658 10952 16722
rect 11016 16658 11032 16722
rect 11096 16658 11112 16722
rect 11176 16658 11192 16722
rect 11256 16658 11264 16722
rect 10944 15634 11264 16658
rect 10944 15570 10952 15634
rect 11016 15570 11032 15634
rect 11096 15570 11112 15634
rect 11176 15570 11192 15634
rect 11256 15570 11264 15634
rect 10944 14546 11264 15570
rect 10944 14482 10952 14546
rect 11016 14482 11032 14546
rect 11096 14482 11112 14546
rect 11176 14482 11192 14546
rect 11256 14482 11264 14546
rect 10944 13458 11264 14482
rect 10944 13394 10952 13458
rect 11016 13394 11032 13458
rect 11096 13394 11112 13458
rect 11176 13394 11192 13458
rect 11256 13394 11264 13458
rect 10944 12370 11264 13394
rect 10944 12306 10952 12370
rect 11016 12306 11032 12370
rect 11096 12306 11112 12370
rect 11176 12306 11192 12370
rect 11256 12306 11264 12370
rect 10944 11282 11264 12306
rect 10944 11218 10952 11282
rect 11016 11218 11032 11282
rect 11096 11218 11112 11282
rect 11176 11218 11192 11282
rect 11256 11218 11264 11282
rect 10944 10194 11264 11218
rect 10944 10130 10952 10194
rect 11016 10130 11032 10194
rect 11096 10130 11112 10194
rect 11176 10130 11192 10194
rect 11256 10130 11264 10194
rect 10944 9106 11264 10130
rect 10944 9042 10952 9106
rect 11016 9042 11032 9106
rect 11096 9042 11112 9106
rect 11176 9042 11192 9106
rect 11256 9042 11264 9106
rect 10944 8018 11264 9042
rect 10944 7954 10952 8018
rect 11016 7954 11032 8018
rect 11096 7954 11112 8018
rect 11176 7954 11192 8018
rect 11256 7954 11264 8018
rect 10944 6930 11264 7954
rect 10944 6866 10952 6930
rect 11016 6866 11032 6930
rect 11096 6866 11112 6930
rect 11176 6866 11192 6930
rect 11256 6866 11264 6930
rect 10944 5842 11264 6866
rect 10944 5778 10952 5842
rect 11016 5778 11032 5842
rect 11096 5778 11112 5842
rect 11176 5778 11192 5842
rect 11256 5778 11264 5842
rect 10944 4754 11264 5778
rect 10944 4690 10952 4754
rect 11016 4690 11032 4754
rect 11096 4690 11112 4754
rect 11176 4690 11192 4754
rect 11256 4690 11264 4754
rect 10944 3666 11264 4690
rect 10944 3602 10952 3666
rect 11016 3602 11032 3666
rect 11096 3602 11112 3666
rect 11176 3602 11192 3666
rect 11256 3602 11264 3666
rect 10944 2578 11264 3602
rect 10944 2514 10952 2578
rect 11016 2514 11032 2578
rect 11096 2514 11112 2578
rect 11176 2514 11192 2578
rect 11256 2514 11264 2578
rect 10944 1954 11264 2514
rect 15944 21618 16264 21634
rect 15944 21554 15952 21618
rect 16016 21554 16032 21618
rect 16096 21554 16112 21618
rect 16176 21554 16192 21618
rect 16256 21554 16264 21618
rect 15944 20530 16264 21554
rect 15944 20466 15952 20530
rect 16016 20466 16032 20530
rect 16096 20466 16112 20530
rect 16176 20466 16192 20530
rect 16256 20466 16264 20530
rect 15944 19442 16264 20466
rect 15944 19378 15952 19442
rect 16016 19378 16032 19442
rect 16096 19378 16112 19442
rect 16176 19378 16192 19442
rect 16256 19378 16264 19442
rect 15944 18354 16264 19378
rect 15944 18290 15952 18354
rect 16016 18290 16032 18354
rect 16096 18290 16112 18354
rect 16176 18290 16192 18354
rect 16256 18290 16264 18354
rect 15944 17266 16264 18290
rect 15944 17202 15952 17266
rect 16016 17202 16032 17266
rect 16096 17202 16112 17266
rect 16176 17202 16192 17266
rect 16256 17202 16264 17266
rect 15944 16178 16264 17202
rect 15944 16114 15952 16178
rect 16016 16114 16032 16178
rect 16096 16114 16112 16178
rect 16176 16114 16192 16178
rect 16256 16114 16264 16178
rect 15944 15090 16264 16114
rect 15944 15026 15952 15090
rect 16016 15026 16032 15090
rect 16096 15026 16112 15090
rect 16176 15026 16192 15090
rect 16256 15026 16264 15090
rect 15944 14002 16264 15026
rect 15944 13938 15952 14002
rect 16016 13938 16032 14002
rect 16096 13938 16112 14002
rect 16176 13938 16192 14002
rect 16256 13938 16264 14002
rect 15944 12914 16264 13938
rect 15944 12850 15952 12914
rect 16016 12850 16032 12914
rect 16096 12850 16112 12914
rect 16176 12850 16192 12914
rect 16256 12850 16264 12914
rect 15944 11826 16264 12850
rect 15944 11762 15952 11826
rect 16016 11762 16032 11826
rect 16096 11762 16112 11826
rect 16176 11762 16192 11826
rect 16256 11762 16264 11826
rect 15944 10738 16264 11762
rect 15944 10674 15952 10738
rect 16016 10674 16032 10738
rect 16096 10674 16112 10738
rect 16176 10674 16192 10738
rect 16256 10674 16264 10738
rect 15944 9650 16264 10674
rect 15944 9586 15952 9650
rect 16016 9586 16032 9650
rect 16096 9586 16112 9650
rect 16176 9586 16192 9650
rect 16256 9586 16264 9650
rect 15944 8562 16264 9586
rect 15944 8498 15952 8562
rect 16016 8498 16032 8562
rect 16096 8498 16112 8562
rect 16176 8498 16192 8562
rect 16256 8498 16264 8562
rect 15944 7474 16264 8498
rect 15944 7410 15952 7474
rect 16016 7410 16032 7474
rect 16096 7410 16112 7474
rect 16176 7410 16192 7474
rect 16256 7410 16264 7474
rect 15944 6386 16264 7410
rect 15944 6322 15952 6386
rect 16016 6322 16032 6386
rect 16096 6322 16112 6386
rect 16176 6322 16192 6386
rect 16256 6322 16264 6386
rect 15944 5298 16264 6322
rect 15944 5234 15952 5298
rect 16016 5234 16032 5298
rect 16096 5234 16112 5298
rect 16176 5234 16192 5298
rect 16256 5234 16264 5298
rect 15944 4210 16264 5234
rect 15944 4146 15952 4210
rect 16016 4146 16032 4210
rect 16096 4146 16112 4210
rect 16176 4146 16192 4210
rect 16256 4146 16264 4210
rect 15944 3122 16264 4146
rect 15944 3058 15952 3122
rect 16016 3058 16032 3122
rect 16096 3058 16112 3122
rect 16176 3058 16192 3122
rect 16256 3058 16264 3122
rect 15944 2034 16264 3058
rect 15944 1970 15952 2034
rect 16016 1970 16032 2034
rect 16096 1970 16112 2034
rect 16176 1970 16192 2034
rect 16256 1970 16264 2034
rect 15944 1954 16264 1970
rect 20944 21074 21264 21634
rect 20944 21010 20952 21074
rect 21016 21010 21032 21074
rect 21096 21010 21112 21074
rect 21176 21010 21192 21074
rect 21256 21010 21264 21074
rect 20944 19986 21264 21010
rect 20944 19922 20952 19986
rect 21016 19922 21032 19986
rect 21096 19922 21112 19986
rect 21176 19922 21192 19986
rect 21256 19922 21264 19986
rect 20944 18898 21264 19922
rect 20944 18834 20952 18898
rect 21016 18834 21032 18898
rect 21096 18834 21112 18898
rect 21176 18834 21192 18898
rect 21256 18834 21264 18898
rect 20944 17810 21264 18834
rect 20944 17746 20952 17810
rect 21016 17746 21032 17810
rect 21096 17746 21112 17810
rect 21176 17746 21192 17810
rect 21256 17746 21264 17810
rect 20944 16722 21264 17746
rect 20944 16658 20952 16722
rect 21016 16658 21032 16722
rect 21096 16658 21112 16722
rect 21176 16658 21192 16722
rect 21256 16658 21264 16722
rect 20944 15634 21264 16658
rect 20944 15570 20952 15634
rect 21016 15570 21032 15634
rect 21096 15570 21112 15634
rect 21176 15570 21192 15634
rect 21256 15570 21264 15634
rect 20944 14546 21264 15570
rect 20944 14482 20952 14546
rect 21016 14482 21032 14546
rect 21096 14482 21112 14546
rect 21176 14482 21192 14546
rect 21256 14482 21264 14546
rect 20944 13458 21264 14482
rect 20944 13394 20952 13458
rect 21016 13394 21032 13458
rect 21096 13394 21112 13458
rect 21176 13394 21192 13458
rect 21256 13394 21264 13458
rect 20944 12370 21264 13394
rect 20944 12306 20952 12370
rect 21016 12306 21032 12370
rect 21096 12306 21112 12370
rect 21176 12306 21192 12370
rect 21256 12306 21264 12370
rect 20944 11282 21264 12306
rect 20944 11218 20952 11282
rect 21016 11218 21032 11282
rect 21096 11218 21112 11282
rect 21176 11218 21192 11282
rect 21256 11218 21264 11282
rect 20944 10194 21264 11218
rect 20944 10130 20952 10194
rect 21016 10130 21032 10194
rect 21096 10130 21112 10194
rect 21176 10130 21192 10194
rect 21256 10130 21264 10194
rect 20944 9106 21264 10130
rect 20944 9042 20952 9106
rect 21016 9042 21032 9106
rect 21096 9042 21112 9106
rect 21176 9042 21192 9106
rect 21256 9042 21264 9106
rect 20944 8018 21264 9042
rect 20944 7954 20952 8018
rect 21016 7954 21032 8018
rect 21096 7954 21112 8018
rect 21176 7954 21192 8018
rect 21256 7954 21264 8018
rect 20944 6930 21264 7954
rect 20944 6866 20952 6930
rect 21016 6866 21032 6930
rect 21096 6866 21112 6930
rect 21176 6866 21192 6930
rect 21256 6866 21264 6930
rect 20944 5842 21264 6866
rect 20944 5778 20952 5842
rect 21016 5778 21032 5842
rect 21096 5778 21112 5842
rect 21176 5778 21192 5842
rect 21256 5778 21264 5842
rect 20944 4754 21264 5778
rect 20944 4690 20952 4754
rect 21016 4690 21032 4754
rect 21096 4690 21112 4754
rect 21176 4690 21192 4754
rect 21256 4690 21264 4754
rect 20944 3666 21264 4690
rect 20944 3602 20952 3666
rect 21016 3602 21032 3666
rect 21096 3602 21112 3666
rect 21176 3602 21192 3666
rect 21256 3602 21264 3666
rect 20944 2578 21264 3602
rect 20944 2514 20952 2578
rect 21016 2514 21032 2578
rect 21096 2514 21112 2578
rect 21176 2514 21192 2578
rect 21256 2514 21264 2578
rect 20944 1954 21264 2514
rect 25944 21618 26264 21634
rect 25944 21554 25952 21618
rect 26016 21554 26032 21618
rect 26096 21554 26112 21618
rect 26176 21554 26192 21618
rect 26256 21554 26264 21618
rect 25944 20530 26264 21554
rect 25944 20466 25952 20530
rect 26016 20466 26032 20530
rect 26096 20466 26112 20530
rect 26176 20466 26192 20530
rect 26256 20466 26264 20530
rect 25944 19442 26264 20466
rect 25944 19378 25952 19442
rect 26016 19378 26032 19442
rect 26096 19378 26112 19442
rect 26176 19378 26192 19442
rect 26256 19378 26264 19442
rect 25944 18354 26264 19378
rect 25944 18290 25952 18354
rect 26016 18290 26032 18354
rect 26096 18290 26112 18354
rect 26176 18290 26192 18354
rect 26256 18290 26264 18354
rect 25944 17266 26264 18290
rect 25944 17202 25952 17266
rect 26016 17202 26032 17266
rect 26096 17202 26112 17266
rect 26176 17202 26192 17266
rect 26256 17202 26264 17266
rect 25944 16178 26264 17202
rect 25944 16114 25952 16178
rect 26016 16114 26032 16178
rect 26096 16114 26112 16178
rect 26176 16114 26192 16178
rect 26256 16114 26264 16178
rect 25944 15090 26264 16114
rect 25944 15026 25952 15090
rect 26016 15026 26032 15090
rect 26096 15026 26112 15090
rect 26176 15026 26192 15090
rect 26256 15026 26264 15090
rect 25944 14002 26264 15026
rect 25944 13938 25952 14002
rect 26016 13938 26032 14002
rect 26096 13938 26112 14002
rect 26176 13938 26192 14002
rect 26256 13938 26264 14002
rect 25944 12914 26264 13938
rect 25944 12850 25952 12914
rect 26016 12850 26032 12914
rect 26096 12850 26112 12914
rect 26176 12850 26192 12914
rect 26256 12850 26264 12914
rect 25944 11826 26264 12850
rect 25944 11762 25952 11826
rect 26016 11762 26032 11826
rect 26096 11762 26112 11826
rect 26176 11762 26192 11826
rect 26256 11762 26264 11826
rect 25944 10738 26264 11762
rect 25944 10674 25952 10738
rect 26016 10674 26032 10738
rect 26096 10674 26112 10738
rect 26176 10674 26192 10738
rect 26256 10674 26264 10738
rect 25944 9650 26264 10674
rect 25944 9586 25952 9650
rect 26016 9586 26032 9650
rect 26096 9586 26112 9650
rect 26176 9586 26192 9650
rect 26256 9586 26264 9650
rect 25944 8562 26264 9586
rect 25944 8498 25952 8562
rect 26016 8498 26032 8562
rect 26096 8498 26112 8562
rect 26176 8498 26192 8562
rect 26256 8498 26264 8562
rect 25944 7474 26264 8498
rect 25944 7410 25952 7474
rect 26016 7410 26032 7474
rect 26096 7410 26112 7474
rect 26176 7410 26192 7474
rect 26256 7410 26264 7474
rect 25944 6386 26264 7410
rect 25944 6322 25952 6386
rect 26016 6322 26032 6386
rect 26096 6322 26112 6386
rect 26176 6322 26192 6386
rect 26256 6322 26264 6386
rect 25944 5298 26264 6322
rect 25944 5234 25952 5298
rect 26016 5234 26032 5298
rect 26096 5234 26112 5298
rect 26176 5234 26192 5298
rect 26256 5234 26264 5298
rect 25944 4210 26264 5234
rect 25944 4146 25952 4210
rect 26016 4146 26032 4210
rect 26096 4146 26112 4210
rect 26176 4146 26192 4210
rect 26256 4146 26264 4210
rect 25944 3122 26264 4146
rect 25944 3058 25952 3122
rect 26016 3058 26032 3122
rect 26096 3058 26112 3122
rect 26176 3058 26192 3122
rect 26256 3058 26264 3122
rect 25944 2034 26264 3058
rect 25944 1970 25952 2034
rect 26016 1970 26032 2034
rect 26096 1970 26112 2034
rect 26176 1970 26192 2034
rect 26256 1970 26264 2034
rect 25944 1954 26264 1970
use sky130_fd_sc_hd__fill_2  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1748 0 1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7
timestamp 1604666999
transform 1 0 1748 0 -1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1932 0 -1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__15__A
timestamp 1604666999
transform 1 0 1932 0 1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1104 0 1 2546
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604666999
transform 1 0 1104 0 -1 2546
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _35_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 2546
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1604666999
transform 1 0 1380 0 1 2546
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2116 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_11
timestamp 1604666999
transform 1 0 2116 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604666999
transform 1 0 3956 0 1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3220 0 -1 2546
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604666999
transform 1 0 4048 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_23
timestamp 1604666999
transform 1 0 3220 0 1 2546
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1604666999
transform 1 0 4048 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604666999
transform 1 0 5152 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6256 0 -1 2546
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1604666999
transform 1 0 5152 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1604666999
transform 1 0 6256 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604666999
transform 1 0 6808 0 -1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604666999
transform 1 0 6900 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604666999
transform 1 0 8004 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1604666999
transform 1 0 7360 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604666999
transform 1 0 9660 0 -1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604666999
transform 1 0 9568 0 1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604666999
transform 1 0 9108 0 -1 2546
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604666999
transform 1 0 9752 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1604666999
transform 1 0 8464 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1604666999
transform 1 0 9660 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604666999
transform 1 0 10856 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604666999
transform 1 0 11960 0 -1 2546
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_105
timestamp 1604666999
transform 1 0 10764 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1604666999
transform 1 0 11868 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604666999
transform 1 0 12512 0 -1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604666999
transform 1 0 12604 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604666999
transform 1 0 13708 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1604666999
transform 1 0 12972 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604666999
transform 1 0 15364 0 -1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604666999
transform 1 0 15180 0 1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604666999
transform 1 0 14812 0 -1 2546
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604666999
transform 1 0 15456 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_141
timestamp 1604666999
transform 1 0 14076 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1604666999
transform 1 0 15272 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604666999
transform 1 0 16560 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_166
timestamp 1604666999
transform 1 0 16376 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_178
timestamp 1604666999
transform 1 0 17480 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604666999
transform 1 0 18216 0 -1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604666999
transform 1 0 17664 0 -1 2546
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604666999
transform 1 0 18308 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1604666999
transform 1 0 18584 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604666999
transform 1 0 21068 0 -1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604666999
transform 1 0 20792 0 1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604666999
transform 1 0 19412 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604666999
transform 1 0 20516 0 -1 2546
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604666999
transform 1 0 21160 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_202
timestamp 1604666999
transform 1 0 19688 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_215
timestamp 1604666999
transform 1 0 20884 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604666999
transform 1 0 22264 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_227
timestamp 1604666999
transform 1 0 21988 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_245 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 23644 0 1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_239
timestamp 1604666999
transform 1 0 23092 0 1 2546
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604666999
transform 1 0 23368 0 -1 2546
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1604666999
transform 1 0 23736 0 1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_252
timestamp 1604666999
transform 1 0 24288 0 1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 24748 0 -1 2546
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1604666999
transform 1 0 24380 0 -1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__12__A
timestamp 1604666999
transform 1 0 24564 0 -1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__14__A
timestamp 1604666999
transform 1 0 24472 0 1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604666999
transform 1 0 23920 0 -1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1604666999
transform 1 0 23920 0 1 2546
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1604666999
transform 1 0 24012 0 -1 2546
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_256
timestamp 1604666999
transform 1 0 24656 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1604666999
transform 1 0 25116 0 -1 2546
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604666999
transform 1 0 26404 0 1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__16__A
timestamp 1604666999
transform 1 0 25668 0 -1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_265
timestamp 1604666999
transform 1 0 25484 0 -1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269
timestamp 1604666999
transform 1 0 25852 0 -1 2546
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_277
timestamp 1604666999
transform 1 0 26588 0 -1 2546
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_268
timestamp 1604666999
transform 1 0 25760 0 1 2546
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_274
timestamp 1604666999
transform 1 0 26312 0 1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_276
timestamp 1604666999
transform 1 0 26496 0 1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604666999
transform 1 0 26772 0 -1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1604666999
transform 1 0 26864 0 -1 2546
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_292
timestamp 1604666999
transform 1 0 27968 0 -1 2546
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_288
timestamp 1604666999
transform 1 0 27600 0 1 2546
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_296
timestamp 1604666999
transform 1 0 28336 0 1 2546
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 28888 0 -1 2546
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 28888 0 1 2546
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298
timestamp 1604666999
transform 1 0 28520 0 -1 2546
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604666999
transform 1 0 1380 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604666999
transform 1 0 2484 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1604666999
transform 1 0 4692 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_51
timestamp 1604666999
transform 1 0 5796 0 -1 3634
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59
timestamp 1604666999
transform 1 0 6532 0 -1 3634
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604666999
transform 1 0 6716 0 -1 3634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1604666999
transform 1 0 6808 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_74
timestamp 1604666999
transform 1 0 7912 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_86
timestamp 1604666999
transform 1 0 9016 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_98
timestamp 1604666999
transform 1 0 10120 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_110
timestamp 1604666999
transform 1 0 11224 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604666999
transform 1 0 12328 0 -1 3634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1604666999
transform 1 0 12420 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_135
timestamp 1604666999
transform 1 0 13524 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_147
timestamp 1604666999
transform 1 0 14628 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_159
timestamp 1604666999
transform 1 0 15732 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1604666999
transform 1 0 16836 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604666999
transform 1 0 17940 0 -1 3634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1604666999
transform 1 0 18032 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_196
timestamp 1604666999
transform 1 0 19136 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_208
timestamp 1604666999
transform 1 0 20240 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_220
timestamp 1604666999
transform 1 0 21344 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_232
timestamp 1604666999
transform 1 0 22448 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1604666999
transform 1 0 23920 0 -1 3634
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604666999
transform 1 0 23552 0 -1 3634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_245
timestamp 1604666999
transform 1 0 23644 0 -1 3634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_252
timestamp 1604666999
transform 1 0 24288 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_264
timestamp 1604666999
transform 1 0 25392 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1604666999
transform 1 0 26496 0 -1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_288
timestamp 1604666999
transform 1 0 27600 0 -1 3634
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_296
timestamp 1604666999
transform 1 0 28336 0 -1 3634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 28888 0 -1 3634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604666999
transform 1 0 2484 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604666999
transform 1 0 3956 0 1 3634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1604666999
transform 1 0 3588 0 1 3634
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1604666999
transform 1 0 4048 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1604666999
transform 1 0 5152 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_56
timestamp 1604666999
transform 1 0 6256 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1604666999
transform 1 0 7360 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604666999
transform 1 0 9568 0 1 3634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1604666999
transform 1 0 8464 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1604666999
transform 1 0 9660 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_105
timestamp 1604666999
transform 1 0 10764 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_117
timestamp 1604666999
transform 1 0 11868 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_129
timestamp 1604666999
transform 1 0 12972 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604666999
transform 1 0 15180 0 1 3634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_141
timestamp 1604666999
transform 1 0 14076 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_154
timestamp 1604666999
transform 1 0 15272 0 1 3634
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1604666999
transform 1 0 16284 0 1 3634
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_162
timestamp 1604666999
transform 1 0 16008 0 1 3634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_167
timestamp 1604666999
transform 1 0 16468 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_179
timestamp 1604666999
transform 1 0 17572 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_191
timestamp 1604666999
transform 1 0 18676 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604666999
transform 1 0 20792 0 1 3634
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__09__A
timestamp 1604666999
transform 1 0 21068 0 1 3634
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_203
timestamp 1604666999
transform 1 0 19780 0 1 3634
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_211
timestamp 1604666999
transform 1 0 20516 0 1 3634
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_215
timestamp 1604666999
transform 1 0 20884 0 1 3634
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1604666999
transform 1 0 21436 0 1 3634
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1604666999
transform 1 0 21988 0 1 3634
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_219
timestamp 1604666999
transform 1 0 21252 0 1 3634
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1604666999
transform 1 0 21804 0 1 3634
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_229
timestamp 1604666999
transform 1 0 22172 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1604666999
transform 1 0 23920 0 1 3634
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__10__A
timestamp 1604666999
transform 1 0 24472 0 1 3634
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_241
timestamp 1604666999
transform 1 0 23276 0 1 3634
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_247
timestamp 1604666999
transform 1 0 23828 0 1 3634
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_252
timestamp 1604666999
transform 1 0 24288 0 1 3634
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_256
timestamp 1604666999
transform 1 0 24656 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604666999
transform 1 0 26404 0 1 3634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_268
timestamp 1604666999
transform 1 0 25760 0 1 3634
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_274
timestamp 1604666999
transform 1 0 26312 0 1 3634
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_276
timestamp 1604666999
transform 1 0 26496 0 1 3634
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_288
timestamp 1604666999
transform 1 0 27600 0 1 3634
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_296
timestamp 1604666999
transform 1 0 28336 0 1 3634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 28888 0 1 3634
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604666999
transform 1 0 1380 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604666999
transform 1 0 2484 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_27
timestamp 1604666999
transform 1 0 3588 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_39
timestamp 1604666999
transform 1 0 4692 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_51
timestamp 1604666999
transform 1 0 5796 0 -1 4722
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1604666999
transform 1 0 6532 0 -1 4722
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604666999
transform 1 0 6716 0 -1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1604666999
transform 1 0 6808 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_74
timestamp 1604666999
transform 1 0 7912 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_86
timestamp 1604666999
transform 1 0 9016 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1604666999
transform 1 0 10120 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1604666999
transform 1 0 11224 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604666999
transform 1 0 12328 0 -1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1604666999
transform 1 0 12420 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_135
timestamp 1604666999
transform 1 0 13524 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_147
timestamp 1604666999
transform 1 0 14628 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1604666999
transform 1 0 16284 0 -1 4722
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_159
timestamp 1604666999
transform 1 0 15732 0 -1 4722
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_169
timestamp 1604666999
transform 1 0 16652 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604666999
transform 1 0 17940 0 -1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_181
timestamp 1604666999
transform 1 0 17756 0 -1 4722
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1604666999
transform 1 0 18032 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1604666999
transform 1 0 19136 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _09_
timestamp 1604666999
transform 1 0 20700 0 -1 4722
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_208
timestamp 1604666999
transform 1 0 20240 0 -1 4722
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_212
timestamp 1604666999
transform 1 0 20608 0 -1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_217
timestamp 1604666999
transform 1 0 21068 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_229
timestamp 1604666999
transform 1 0 22172 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604666999
transform 1 0 23552 0 -1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_241
timestamp 1604666999
transform 1 0 23276 0 -1 4722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_245
timestamp 1604666999
transform 1 0 23644 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_257
timestamp 1604666999
transform 1 0 24748 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_269
timestamp 1604666999
transform 1 0 25852 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_281
timestamp 1604666999
transform 1 0 26956 0 -1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_293
timestamp 1604666999
transform 1 0 28060 0 -1 4722
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 28888 0 -1 4722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604666999
transform 1 0 1380 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604666999
transform 1 0 2484 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604666999
transform 1 0 3956 0 1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1604666999
transform 1 0 3588 0 1 4722
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_32
timestamp 1604666999
transform 1 0 4048 0 1 4722
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__07__A
timestamp 1604666999
transform 1 0 4784 0 1 4722
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_42
timestamp 1604666999
transform 1 0 4968 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_54
timestamp 1604666999
transform 1 0 6072 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_66
timestamp 1604666999
transform 1 0 7176 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_78
timestamp 1604666999
transform 1 0 8280 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604666999
transform 1 0 9568 0 1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_90
timestamp 1604666999
transform 1 0 9384 0 1 4722
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1604666999
transform 1 0 9660 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_105
timestamp 1604666999
transform 1 0 10764 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_117
timestamp 1604666999
transform 1 0 11868 0 1 4722
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1604666999
transform 1 0 13708 0 1 4722
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1604666999
transform 1 0 12604 0 1 4722
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_127
timestamp 1604666999
transform 1 0 12788 0 1 4722
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_135
timestamp 1604666999
transform 1 0 13524 0 1 4722
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604666999
transform 1 0 15180 0 1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__08__A
timestamp 1604666999
transform 1 0 14260 0 1 4722
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_141
timestamp 1604666999
transform 1 0 14076 0 1 4722
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_145
timestamp 1604666999
transform 1 0 14444 0 1 4722
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_154
timestamp 1604666999
transform 1 0 15272 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_166
timestamp 1604666999
transform 1 0 16376 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_178
timestamp 1604666999
transform 1 0 17480 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_190
timestamp 1604666999
transform 1 0 18584 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604666999
transform 1 0 20792 0 1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_202
timestamp 1604666999
transform 1 0 19688 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_215
timestamp 1604666999
transform 1 0 20884 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_227
timestamp 1604666999
transform 1 0 21988 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1604666999
transform 1 0 23920 0 1 4722
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1604666999
transform 1 0 24472 0 1 4722
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_239
timestamp 1604666999
transform 1 0 23092 0 1 4722
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_247
timestamp 1604666999
transform 1 0 23828 0 1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_252
timestamp 1604666999
transform 1 0 24288 0 1 4722
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_256
timestamp 1604666999
transform 1 0 24656 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604666999
transform 1 0 26404 0 1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_268
timestamp 1604666999
transform 1 0 25760 0 1 4722
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_274
timestamp 1604666999
transform 1 0 26312 0 1 4722
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_276
timestamp 1604666999
transform 1 0 26496 0 1 4722
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_288
timestamp 1604666999
transform 1 0 27600 0 1 4722
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_296
timestamp 1604666999
transform 1 0 28336 0 1 4722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 28888 0 1 4722
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604666999
transform 1 0 1380 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604666999
transform 1 0 2484 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604666999
transform 1 0 1380 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604666999
transform 1 0 2484 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604666999
transform 1 0 3956 0 1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_27
timestamp 1604666999
transform 1 0 3588 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_39
timestamp 1604666999
transform 1 0 4692 0 -1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1604666999
transform 1 0 3588 0 1 5810
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1604666999
transform 1 0 4048 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _07_
timestamp 1604666999
transform 1 0 4784 0 -1 5810
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604666999
transform 1 0 5152 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_56
timestamp 1604666999
transform 1 0 6256 0 -1 5810
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1604666999
transform 1 0 5152 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_56
timestamp 1604666999
transform 1 0 6256 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604666999
transform 1 0 6716 0 -1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_60
timestamp 1604666999
transform 1 0 6624 0 -1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_62
timestamp 1604666999
transform 1 0 6808 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1604666999
transform 1 0 7912 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1604666999
transform 1 0 7360 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604666999
transform 1 0 9568 0 1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_86
timestamp 1604666999
transform 1 0 9016 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_98
timestamp 1604666999
transform 1 0 10120 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1604666999
transform 1 0 8464 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1604666999
transform 1 0 9660 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__05__A
timestamp 1604666999
transform 1 0 10856 0 1 5810
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_110
timestamp 1604666999
transform 1 0 11224 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_105
timestamp 1604666999
transform 1 0 10764 0 1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_108
timestamp 1604666999
transform 1 0 11040 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1604666999
transform 1 0 12604 0 -1 5810
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604666999
transform 1 0 12328 0 -1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_123
timestamp 1604666999
transform 1 0 12420 0 -1 5810
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604666999
transform 1 0 12972 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_120
timestamp 1604666999
transform 1 0 12144 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_132
timestamp 1604666999
transform 1 0 13248 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604666999
transform 1 0 15180 0 1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__06__A
timestamp 1604666999
transform 1 0 14628 0 1 5810
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604666999
transform 1 0 14076 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1604666999
transform 1 0 15180 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_144
timestamp 1604666999
transform 1 0 14352 0 1 5810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_149
timestamp 1604666999
transform 1 0 14812 0 1 5810
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_154
timestamp 1604666999
transform 1 0 15272 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1604666999
transform 1 0 16284 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_177
timestamp 1604666999
transform 1 0 17388 0 -1 5810
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_166
timestamp 1604666999
transform 1 0 16376 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_178
timestamp 1604666999
transform 1 0 17480 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604666999
transform 1 0 17940 0 -1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1604666999
transform 1 0 18032 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1604666999
transform 1 0 19136 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_190
timestamp 1604666999
transform 1 0 18584 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604666999
transform 1 0 20792 0 1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_208
timestamp 1604666999
transform 1 0 20240 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_202
timestamp 1604666999
transform 1 0 19688 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_215
timestamp 1604666999
transform 1 0 20884 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_220
timestamp 1604666999
transform 1 0 21344 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_232
timestamp 1604666999
transform 1 0 22448 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_227
timestamp 1604666999
transform 1 0 21988 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604666999
transform 1 0 23552 0 -1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1604666999
transform 1 0 23920 0 1 5810
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_245
timestamp 1604666999
transform 1 0 23644 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_257
timestamp 1604666999
transform 1 0 24748 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_239
timestamp 1604666999
transform 1 0 23092 0 1 5810
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_247
timestamp 1604666999
transform 1 0 23828 0 1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_250
timestamp 1604666999
transform 1 0 24104 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604666999
transform 1 0 26404 0 1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_269
timestamp 1604666999
transform 1 0 25852 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_262
timestamp 1604666999
transform 1 0 25208 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_274
timestamp 1604666999
transform 1 0 26312 0 1 5810
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_276
timestamp 1604666999
transform 1 0 26496 0 1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_281
timestamp 1604666999
transform 1 0 26956 0 -1 5810
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_293
timestamp 1604666999
transform 1 0 28060 0 -1 5810
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_288
timestamp 1604666999
transform 1 0 27600 0 1 5810
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_296
timestamp 1604666999
transform 1 0 28336 0 1 5810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 28888 0 -1 5810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 28888 0 1 5810
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 6898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604666999
transform 1 0 1380 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604666999
transform 1 0 2484 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_27
timestamp 1604666999
transform 1 0 3588 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_39
timestamp 1604666999
transform 1 0 4692 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1604666999
transform 1 0 5796 0 -1 6898
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1604666999
transform 1 0 6532 0 -1 6898
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604666999
transform 1 0 6716 0 -1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1604666999
transform 1 0 6808 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_74
timestamp 1604666999
transform 1 0 7912 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_86
timestamp 1604666999
transform 1 0 9016 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_98
timestamp 1604666999
transform 1 0 10120 0 -1 6898
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1604666999
transform 1 0 10856 0 -1 6898
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_110
timestamp 1604666999
transform 1 0 11224 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604666999
transform 1 0 12328 0 -1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1604666999
transform 1 0 12420 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_135
timestamp 1604666999
transform 1 0 13524 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _06_
timestamp 1604666999
transform 1 0 14628 0 -1 6898
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_151
timestamp 1604666999
transform 1 0 14996 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_163
timestamp 1604666999
transform 1 0 16100 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_175
timestamp 1604666999
transform 1 0 17204 0 -1 6898
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604666999
transform 1 0 17940 0 -1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1604666999
transform 1 0 18032 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_196
timestamp 1604666999
transform 1 0 19136 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_208
timestamp 1604666999
transform 1 0 20240 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_220
timestamp 1604666999
transform 1 0 21344 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_232
timestamp 1604666999
transform 1 0 22448 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1604666999
transform 1 0 23920 0 -1 6898
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604666999
transform 1 0 23552 0 -1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_245
timestamp 1604666999
transform 1 0 23644 0 -1 6898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_252
timestamp 1604666999
transform 1 0 24288 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_264
timestamp 1604666999
transform 1 0 25392 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_276
timestamp 1604666999
transform 1 0 26496 0 -1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_288
timestamp 1604666999
transform 1 0 27600 0 -1 6898
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_296
timestamp 1604666999
transform 1 0 28336 0 -1 6898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 28888 0 -1 6898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 6898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604666999
transform 1 0 1380 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604666999
transform 1 0 2484 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604666999
transform 1 0 3956 0 1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1604666999
transform 1 0 3588 0 1 6898
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1604666999
transform 1 0 4048 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1604666999
transform 1 0 5152 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_56
timestamp 1604666999
transform 1 0 6256 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_68
timestamp 1604666999
transform 1 0 7360 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604666999
transform 1 0 9568 0 1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_80
timestamp 1604666999
transform 1 0 8464 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1604666999
transform 1 0 9660 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_105
timestamp 1604666999
transform 1 0 10764 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_117
timestamp 1604666999
transform 1 0 11868 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_129
timestamp 1604666999
transform 1 0 12972 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604666999
transform 1 0 15180 0 1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_141
timestamp 1604666999
transform 1 0 14076 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_154
timestamp 1604666999
transform 1 0 15272 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_166
timestamp 1604666999
transform 1 0 16376 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_178
timestamp 1604666999
transform 1 0 17480 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _04_
timestamp 1604666999
transform 1 0 18676 0 1 6898
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__04__A
timestamp 1604666999
transform 1 0 19228 0 1 6898
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_190
timestamp 1604666999
transform 1 0 18584 0 1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_195
timestamp 1604666999
transform 1 0 19044 0 1 6898
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604666999
transform 1 0 20792 0 1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_199
timestamp 1604666999
transform 1 0 19412 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_211
timestamp 1604666999
transform 1 0 20516 0 1 6898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_215
timestamp 1604666999
transform 1 0 20884 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1604666999
transform 1 0 22448 0 1 6898
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1604666999
transform 1 0 23000 0 1 6898
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_227
timestamp 1604666999
transform 1 0 21988 0 1 6898
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_231
timestamp 1604666999
transform 1 0 22356 0 1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1604666999
transform 1 0 22816 0 1 6898
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__03__A
timestamp 1604666999
transform 1 0 23920 0 1 6898
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_240
timestamp 1604666999
transform 1 0 23184 0 1 6898
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_250
timestamp 1604666999
transform 1 0 24104 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604666999
transform 1 0 26404 0 1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_262
timestamp 1604666999
transform 1 0 25208 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_274
timestamp 1604666999
transform 1 0 26312 0 1 6898
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_276
timestamp 1604666999
transform 1 0 26496 0 1 6898
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_288
timestamp 1604666999
transform 1 0 27600 0 1 6898
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_296
timestamp 1604666999
transform 1 0 28336 0 1 6898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 28888 0 1 6898
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 7986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604666999
transform 1 0 1380 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604666999
transform 1 0 2484 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1604666999
transform 1 0 3588 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1604666999
transform 1 0 4692 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1604666999
transform 1 0 5796 0 -1 7986
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1604666999
transform 1 0 6532 0 -1 7986
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604666999
transform 1 0 6716 0 -1 7986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_62
timestamp 1604666999
transform 1 0 6808 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1604666999
transform 1 0 7912 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_86
timestamp 1604666999
transform 1 0 9016 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_98
timestamp 1604666999
transform 1 0 10120 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_110
timestamp 1604666999
transform 1 0 11224 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604666999
transform 1 0 12328 0 -1 7986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1604666999
transform 1 0 12420 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_135
timestamp 1604666999
transform 1 0 13524 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_147
timestamp 1604666999
transform 1 0 14628 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_159
timestamp 1604666999
transform 1 0 15732 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_171
timestamp 1604666999
transform 1 0 16836 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604666999
transform 1 0 17940 0 -1 7986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_184
timestamp 1604666999
transform 1 0 18032 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_196
timestamp 1604666999
transform 1 0 19136 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_208
timestamp 1604666999
transform 1 0 20240 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_220
timestamp 1604666999
transform 1 0 21344 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_232
timestamp 1604666999
transform 1 0 22448 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _03_
timestamp 1604666999
transform 1 0 23920 0 -1 7986
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604666999
transform 1 0 23552 0 -1 7986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_245
timestamp 1604666999
transform 1 0 23644 0 -1 7986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_252
timestamp 1604666999
transform 1 0 24288 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_264
timestamp 1604666999
transform 1 0 25392 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_276
timestamp 1604666999
transform 1 0 26496 0 -1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_288
timestamp 1604666999
transform 1 0 27600 0 -1 7986
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_296
timestamp 1604666999
transform 1 0 28336 0 -1 7986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 28888 0 -1 7986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 7986
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604666999
transform 1 0 1564 0 1 7986
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1604666999
transform 1 0 1380 0 1 7986
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_7
timestamp 1604666999
transform 1 0 1748 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_19
timestamp 1604666999
transform 1 0 2852 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604666999
transform 1 0 3956 0 1 7986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1604666999
transform 1 0 4048 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1604666999
transform 1 0 5152 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_56
timestamp 1604666999
transform 1 0 6256 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1604666999
transform 1 0 7360 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604666999
transform 1 0 9568 0 1 7986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1604666999
transform 1 0 8464 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1604666999
transform 1 0 9660 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_105
timestamp 1604666999
transform 1 0 10764 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_117
timestamp 1604666999
transform 1 0 11868 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_129
timestamp 1604666999
transform 1 0 12972 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604666999
transform 1 0 15180 0 1 7986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_141
timestamp 1604666999
transform 1 0 14076 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_154
timestamp 1604666999
transform 1 0 15272 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_166
timestamp 1604666999
transform 1 0 16376 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_178
timestamp 1604666999
transform 1 0 17480 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_190
timestamp 1604666999
transform 1 0 18584 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604666999
transform 1 0 20792 0 1 7986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_202
timestamp 1604666999
transform 1 0 19688 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_215
timestamp 1604666999
transform 1 0 20884 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_227
timestamp 1604666999
transform 1 0 21988 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1604666999
transform 1 0 23920 0 1 7986
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__02__A
timestamp 1604666999
transform 1 0 24472 0 1 7986
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1604666999
transform 1 0 23736 0 1 7986
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_239
timestamp 1604666999
transform 1 0 23092 0 1 7986
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_245
timestamp 1604666999
transform 1 0 23644 0 1 7986
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_252
timestamp 1604666999
transform 1 0 24288 0 1 7986
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_256
timestamp 1604666999
transform 1 0 24656 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604666999
transform 1 0 26404 0 1 7986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_268
timestamp 1604666999
transform 1 0 25760 0 1 7986
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_274
timestamp 1604666999
transform 1 0 26312 0 1 7986
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_276
timestamp 1604666999
transform 1 0 26496 0 1 7986
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_288
timestamp 1604666999
transform 1 0 27600 0 1 7986
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_296
timestamp 1604666999
transform 1 0 28336 0 1 7986
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 28888 0 1 7986
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604666999
transform 1 0 1380 0 -1 9074
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_7
timestamp 1604666999
transform 1 0 1748 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_19
timestamp 1604666999
transform 1 0 2852 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_31
timestamp 1604666999
transform 1 0 3956 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_43
timestamp 1604666999
transform 1 0 5060 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_55
timestamp 1604666999
transform 1 0 6164 0 -1 9074
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 6716 0 -1 9074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1604666999
transform 1 0 6808 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_74
timestamp 1604666999
transform 1 0 7912 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_86
timestamp 1604666999
transform 1 0 9016 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_98
timestamp 1604666999
transform 1 0 10120 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_110
timestamp 1604666999
transform 1 0 11224 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 12328 0 -1 9074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1604666999
transform 1 0 12420 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_135
timestamp 1604666999
transform 1 0 13524 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_147
timestamp 1604666999
transform 1 0 14628 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_159
timestamp 1604666999
transform 1 0 15732 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_171
timestamp 1604666999
transform 1 0 16836 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 17940 0 -1 9074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_184
timestamp 1604666999
transform 1 0 18032 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_196
timestamp 1604666999
transform 1 0 19136 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_208
timestamp 1604666999
transform 1 0 20240 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_220
timestamp 1604666999
transform 1 0 21344 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_232
timestamp 1604666999
transform 1 0 22448 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _02_
timestamp 1604666999
transform 1 0 23920 0 -1 9074
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 23552 0 -1 9074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_245
timestamp 1604666999
transform 1 0 23644 0 -1 9074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_252
timestamp 1604666999
transform 1 0 24288 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_264
timestamp 1604666999
transform 1 0 25392 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1604666999
transform 1 0 26496 0 -1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_288
timestamp 1604666999
transform 1 0 27600 0 -1 9074
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_296
timestamp 1604666999
transform 1 0 28336 0 -1 9074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 28888 0 -1 9074
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604666999
transform 1 0 1748 0 1 9074
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1604666999
transform 1 0 1932 0 1 9074
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10162
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9074
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604666999
transform 1 0 1380 0 1 9074
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1604666999
transform 1 0 1380 0 -1 10162
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1604666999
transform 1 0 2116 0 1 9074
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604666999
transform 1 0 2300 0 1 9074
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_19
timestamp 1604666999
transform 1 0 2852 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_7
timestamp 1604666999
transform 1 0 1748 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604666999
transform 1 0 2484 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 3956 0 1 9074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1604666999
transform 1 0 3588 0 1 9074
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1604666999
transform 1 0 4048 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_31
timestamp 1604666999
transform 1 0 3956 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1604666999
transform 1 0 5152 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_56
timestamp 1604666999
transform 1 0 6256 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_43
timestamp 1604666999
transform 1 0 5060 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_55
timestamp 1604666999
transform 1 0 6164 0 -1 10162
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 6716 0 -1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 7912 0 -1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8280 0 -1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_68
timestamp 1604666999
transform 1 0 7360 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_62
timestamp 1604666999
transform 1 0 6808 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_76
timestamp 1604666999
transform 1 0 8096 0 -1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 9568 0 1 9074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_80
timestamp 1604666999
transform 1 0 8464 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1604666999
transform 1 0 9660 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604666999
transform 1 0 8464 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_92
timestamp 1604666999
transform 1 0 9568 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_105
timestamp 1604666999
transform 1 0 10764 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_117
timestamp 1604666999
transform 1 0 11868 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_104
timestamp 1604666999
transform 1 0 10672 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_116
timestamp 1604666999
transform 1 0 11776 0 -1 10162
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 12328 0 -1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_129
timestamp 1604666999
transform 1 0 12972 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1604666999
transform 1 0 12420 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_135
timestamp 1604666999
transform 1 0 13524 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 15180 0 1 9074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_141
timestamp 1604666999
transform 1 0 14076 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_154
timestamp 1604666999
transform 1 0 15272 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_147
timestamp 1604666999
transform 1 0 14628 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_166
timestamp 1604666999
transform 1 0 16376 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_178
timestamp 1604666999
transform 1 0 17480 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_159
timestamp 1604666999
transform 1 0 15732 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_171
timestamp 1604666999
transform 1 0 16836 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 17940 0 -1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_190
timestamp 1604666999
transform 1 0 18584 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_184
timestamp 1604666999
transform 1 0 18032 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_196
timestamp 1604666999
transform 1 0 19136 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 20792 0 1 9074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_202
timestamp 1604666999
transform 1 0 19688 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_215
timestamp 1604666999
transform 1 0 20884 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_208
timestamp 1604666999
transform 1 0 20240 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_227
timestamp 1604666999
transform 1 0 21988 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_220
timestamp 1604666999
transform 1 0 21344 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_232
timestamp 1604666999
transform 1 0 22448 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604666999
transform 1 0 23920 0 1 9074
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 23552 0 -1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604666999
transform 1 0 24472 0 1 9074
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_239
timestamp 1604666999
transform 1 0 23092 0 1 9074
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_247
timestamp 1604666999
transform 1 0 23828 0 1 9074
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_252
timestamp 1604666999
transform 1 0 24288 0 1 9074
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_256
timestamp 1604666999
transform 1 0 24656 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_245
timestamp 1604666999
transform 1 0 23644 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_257
timestamp 1604666999
transform 1 0 24748 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 26404 0 1 9074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_268
timestamp 1604666999
transform 1 0 25760 0 1 9074
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_274
timestamp 1604666999
transform 1 0 26312 0 1 9074
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_276
timestamp 1604666999
transform 1 0 26496 0 1 9074
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_269
timestamp 1604666999
transform 1 0 25852 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_288
timestamp 1604666999
transform 1 0 27600 0 1 9074
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_296
timestamp 1604666999
transform 1 0 28336 0 1 9074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_281
timestamp 1604666999
transform 1 0 26956 0 -1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_293
timestamp 1604666999
transform 1 0 28060 0 -1 10162
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 28888 0 1 9074
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 28888 0 -1 10162
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604666999
transform 1 0 1380 0 1 10162
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10162
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1604666999
transform 1 0 1932 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1604666999
transform 1 0 2300 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1604666999
transform 1 0 1748 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_11
timestamp 1604666999
transform 1 0 2116 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1604666999
transform 1 0 2484 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 3956 0 1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1604666999
transform 1 0 3588 0 1 10162
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1604666999
transform 1 0 4048 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1604666999
transform 1 0 5152 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_56
timestamp 1604666999
transform 1 0 6256 0 1 10162
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 7912 0 1 10162
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 7728 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 7360 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6992 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1604666999
transform 1 0 7176 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp 1604666999
transform 1 0 7544 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 9568 0 1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 8924 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_83
timestamp 1604666999
transform 1 0 8740 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_87
timestamp 1604666999
transform 1 0 9108 0 1 10162
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_91
timestamp 1604666999
transform 1 0 9476 0 1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1604666999
transform 1 0 9660 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_105
timestamp 1604666999
transform 1 0 10764 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_117
timestamp 1604666999
transform 1 0 11868 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_129
timestamp 1604666999
transform 1 0 12972 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 15180 0 1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_141
timestamp 1604666999
transform 1 0 14076 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_154
timestamp 1604666999
transform 1 0 15272 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_166
timestamp 1604666999
transform 1 0 16376 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_178
timestamp 1604666999
transform 1 0 17480 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_190
timestamp 1604666999
transform 1 0 18584 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 20792 0 1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_202
timestamp 1604666999
transform 1 0 19688 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_215
timestamp 1604666999
transform 1 0 20884 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_227
timestamp 1604666999
transform 1 0 21988 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1604666999
transform 1 0 23920 0 1 10162
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_239
timestamp 1604666999
transform 1 0 23092 0 1 10162
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_247
timestamp 1604666999
transform 1 0 23828 0 1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_250
timestamp 1604666999
transform 1 0 24104 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 26404 0 1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_262
timestamp 1604666999
transform 1 0 25208 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_274
timestamp 1604666999
transform 1 0 26312 0 1 10162
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_276
timestamp 1604666999
transform 1 0 26496 0 1 10162
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_288
timestamp 1604666999
transform 1 0 27600 0 1 10162
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_296
timestamp 1604666999
transform 1 0 28336 0 1 10162
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 28888 0 1 10162
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604666999
transform 1 0 1380 0 -1 11250
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11250
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_7
timestamp 1604666999
transform 1 0 1748 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_19
timestamp 1604666999
transform 1 0 2852 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_31
timestamp 1604666999
transform 1 0 3956 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_43
timestamp 1604666999
transform 1 0 5060 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_55
timestamp 1604666999
transform 1 0 6164 0 -1 11250
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 7728 0 -1 11250
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 6716 0 -1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_62
timestamp 1604666999
transform 1 0 6808 0 -1 11250
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_70
timestamp 1604666999
transform 1 0 7544 0 -1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_81
timestamp 1604666999
transform 1 0 8556 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604666999
transform 1 0 9660 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 12052 0 -1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604666999
transform 1 0 10764 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_117
timestamp 1604666999
transform 1 0 11868 0 -1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 12328 0 -1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_121
timestamp 1604666999
transform 1 0 12236 0 -1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1604666999
transform 1 0 12420 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_135
timestamp 1604666999
transform 1 0 13524 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_147
timestamp 1604666999
transform 1 0 14628 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_159
timestamp 1604666999
transform 1 0 15732 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_171
timestamp 1604666999
transform 1 0 16836 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 17940 0 -1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_184
timestamp 1604666999
transform 1 0 18032 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_196
timestamp 1604666999
transform 1 0 19136 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_208
timestamp 1604666999
transform 1 0 20240 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_220
timestamp 1604666999
transform 1 0 21344 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_232
timestamp 1604666999
transform 1 0 22448 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1604666999
transform 1 0 23920 0 -1 11250
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 23552 0 -1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_245
timestamp 1604666999
transform 1 0 23644 0 -1 11250
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_252
timestamp 1604666999
transform 1 0 24288 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_264
timestamp 1604666999
transform 1 0 25392 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_276
timestamp 1604666999
transform 1 0 26496 0 -1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_288
timestamp 1604666999
transform 1 0 27600 0 -1 11250
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_296
timestamp 1604666999
transform 1 0 28336 0 -1 11250
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 28888 0 -1 11250
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1604666999
transform 1 0 1380 0 1 11250
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11250
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__13__A
timestamp 1604666999
transform 1 0 1932 0 1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604666999
transform 1 0 1748 0 1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_11
timestamp 1604666999
transform 1 0 2116 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 3956 0 1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_23
timestamp 1604666999
transform 1 0 3220 0 1 11250
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1604666999
transform 1 0 4048 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1604666999
transform 1 0 5152 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_56
timestamp 1604666999
transform 1 0 6256 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 7912 0 1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8280 0 1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_68
timestamp 1604666999
transform 1 0 7360 0 1 11250
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_76
timestamp 1604666999
transform 1 0 8096 0 1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 9568 0 1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8648 0 1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_80
timestamp 1604666999
transform 1 0 8464 0 1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_84
timestamp 1604666999
transform 1 0 8832 0 1 11250
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1604666999
transform 1 0 9660 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 12052 0 1 11250
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 11868 0 1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_105
timestamp 1604666999
transform 1 0 10764 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_128
timestamp 1604666999
transform 1 0 12880 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 15180 0 1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_140
timestamp 1604666999
transform 1 0 13984 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_152
timestamp 1604666999
transform 1 0 15088 0 1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_154
timestamp 1604666999
transform 1 0 15272 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_166
timestamp 1604666999
transform 1 0 16376 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_178
timestamp 1604666999
transform 1 0 17480 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_190
timestamp 1604666999
transform 1 0 18584 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 20792 0 1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_202
timestamp 1604666999
transform 1 0 19688 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_215
timestamp 1604666999
transform 1 0 20884 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_227
timestamp 1604666999
transform 1 0 21988 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604666999
transform 1 0 23920 0 1 11250
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604666999
transform 1 0 24472 0 1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_239
timestamp 1604666999
transform 1 0 23092 0 1 11250
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_247
timestamp 1604666999
transform 1 0 23828 0 1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_252
timestamp 1604666999
transform 1 0 24288 0 1 11250
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_256
timestamp 1604666999
transform 1 0 24656 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 26404 0 1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_268
timestamp 1604666999
transform 1 0 25760 0 1 11250
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_274
timestamp 1604666999
transform 1 0 26312 0 1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_276
timestamp 1604666999
transform 1 0 26496 0 1 11250
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_288
timestamp 1604666999
transform 1 0 27600 0 1 11250
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_296
timestamp 1604666999
transform 1 0 28336 0 1 11250
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 28888 0 1 11250
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12338
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1604666999
transform 1 0 1564 0 -1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604666999
transform 1 0 1380 0 -1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_7
timestamp 1604666999
transform 1 0 1748 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_19
timestamp 1604666999
transform 1 0 2852 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_31
timestamp 1604666999
transform 1 0 3956 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_43
timestamp 1604666999
transform 1 0 5060 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_55
timestamp 1604666999
transform 1 0 6164 0 -1 12338
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7912 0 -1 12338
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 6716 0 -1 12338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_62
timestamp 1604666999
transform 1 0 6808 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_83
timestamp 1604666999
transform 1 0 8740 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_95
timestamp 1604666999
transform 1 0 9844 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 12052 0 -1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_107
timestamp 1604666999
transform 1 0 10948 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 12328 0 -1 12338
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 13064 0 -1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 13524 0 -1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1604666999
transform 1 0 12236 0 -1 12338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_123
timestamp 1604666999
transform 1 0 12420 0 -1 12338
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_129
timestamp 1604666999
transform 1 0 12972 0 -1 12338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_132
timestamp 1604666999
transform 1 0 13248 0 -1 12338
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_137
timestamp 1604666999
transform 1 0 13708 0 -1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 13892 0 -1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1604666999
transform 1 0 14076 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1604666999
transform 1 0 15180 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1604666999
transform 1 0 16284 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_177
timestamp 1604666999
transform 1 0 17388 0 -1 12338
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 17940 0 -1 12338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_184
timestamp 1604666999
transform 1 0 18032 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_196
timestamp 1604666999
transform 1 0 19136 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_208
timestamp 1604666999
transform 1 0 20240 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_220
timestamp 1604666999
transform 1 0 21344 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_232
timestamp 1604666999
transform 1 0 22448 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 23552 0 -1 12338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_245
timestamp 1604666999
transform 1 0 23644 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_257
timestamp 1604666999
transform 1 0 24748 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_269
timestamp 1604666999
transform 1 0 25852 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_281
timestamp 1604666999
transform 1 0 26956 0 -1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_293
timestamp 1604666999
transform 1 0 28060 0 -1 12338
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 28888 0 -1 12338
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1604666999
transform 1 0 1380 0 1 12338
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1604666999
transform 1 0 1380 0 -1 13426
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13426
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__11__A
timestamp 1604666999
transform 1 0 1932 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1604666999
transform 1 0 1748 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_11
timestamp 1604666999
transform 1 0 2116 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_7
timestamp 1604666999
transform 1 0 1748 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_19
timestamp 1604666999
transform 1 0 2852 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 3956 0 1 12338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_23
timestamp 1604666999
transform 1 0 3220 0 1 12338
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1604666999
transform 1 0 4048 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_31
timestamp 1604666999
transform 1 0 3956 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1604666999
transform 1 0 5152 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_56
timestamp 1604666999
transform 1 0 6256 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_43
timestamp 1604666999
transform 1 0 5060 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_55
timestamp 1604666999
transform 1 0 6164 0 -1 13426
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 6716 0 -1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_68
timestamp 1604666999
transform 1 0 7360 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_62
timestamp 1604666999
transform 1 0 6808 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_74
timestamp 1604666999
transform 1 0 7912 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 9568 0 1 12338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_80
timestamp 1604666999
transform 1 0 8464 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1604666999
transform 1 0 9660 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_86
timestamp 1604666999
transform 1 0 9016 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_98
timestamp 1604666999
transform 1 0 10120 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_105
timestamp 1604666999
transform 1 0 10764 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_117
timestamp 1604666999
transform 1 0 11868 0 1 12338
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_110
timestamp 1604666999
transform 1 0 11224 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 13064 0 1 12338
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 13524 0 -1 13426
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 12328 0 -1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 12880 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 13064 0 -1 13426
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_125
timestamp 1604666999
transform 1 0 12604 0 1 12338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_123
timestamp 1604666999
transform 1 0 12420 0 -1 13426
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_129
timestamp 1604666999
transform 1 0 12972 0 -1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_132
timestamp 1604666999
transform 1 0 13248 0 -1 13426
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 15180 0 1 12338
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 14076 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_139
timestamp 1604666999
transform 1 0 13892 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_143
timestamp 1604666999
transform 1 0 14260 0 1 12338
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_151
timestamp 1604666999
transform 1 0 14996 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_154
timestamp 1604666999
transform 1 0 15272 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1604666999
transform 1 0 14352 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1604666999
transform 1 0 15456 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_166
timestamp 1604666999
transform 1 0 16376 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_178
timestamp 1604666999
transform 1 0 17480 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_168
timestamp 1604666999
transform 1 0 16560 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 17940 0 -1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_190
timestamp 1604666999
transform 1 0 18584 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_180
timestamp 1604666999
transform 1 0 17664 0 -1 13426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_184
timestamp 1604666999
transform 1 0 18032 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_196
timestamp 1604666999
transform 1 0 19136 0 -1 13426
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1604666999
transform 1 0 20240 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_204
timestamp 1604666999
transform 1 0 19872 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 20056 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 19688 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 19688 0 -1 13426
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_212
timestamp 1604666999
transform 1 0 20608 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 20424 0 1 12338
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 20792 0 1 12338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_211
timestamp 1604666999
transform 1 0 20516 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_215
timestamp 1604666999
transform 1 0 20884 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_227
timestamp 1604666999
transform 1 0 21988 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_223
timestamp 1604666999
transform 1 0 21620 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_235
timestamp 1604666999
transform 1 0 22724 0 -1 13426
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 23552 0 -1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_239
timestamp 1604666999
transform 1 0 23092 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_251
timestamp 1604666999
transform 1 0 24196 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_243
timestamp 1604666999
transform 1 0 23460 0 -1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_245
timestamp 1604666999
transform 1 0 23644 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_257
timestamp 1604666999
transform 1 0 24748 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 26404 0 1 12338
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_263
timestamp 1604666999
transform 1 0 25300 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_276
timestamp 1604666999
transform 1 0 26496 0 1 12338
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_269
timestamp 1604666999
transform 1 0 25852 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_288
timestamp 1604666999
transform 1 0 27600 0 1 12338
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_296
timestamp 1604666999
transform 1 0 28336 0 1 12338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_281
timestamp 1604666999
transform 1 0 26956 0 -1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_293
timestamp 1604666999
transform 1 0 28060 0 -1 13426
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 28888 0 1 12338
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 28888 0 -1 13426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604666999
transform 1 0 1380 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604666999
transform 1 0 2484 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 3956 0 1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1604666999
transform 1 0 3588 0 1 13426
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1604666999
transform 1 0 4048 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_44
timestamp 1604666999
transform 1 0 5152 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_56
timestamp 1604666999
transform 1 0 6256 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_68
timestamp 1604666999
transform 1 0 7360 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 9568 0 1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_80
timestamp 1604666999
transform 1 0 8464 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1604666999
transform 1 0 9660 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_105
timestamp 1604666999
transform 1 0 10764 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_117
timestamp 1604666999
transform 1 0 11868 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_129
timestamp 1604666999
transform 1 0 12972 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 15180 0 1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_141
timestamp 1604666999
transform 1 0 14076 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_154
timestamp 1604666999
transform 1 0 15272 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_166
timestamp 1604666999
transform 1 0 16376 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_178
timestamp 1604666999
transform 1 0 17480 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _01_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 19044 0 1 13426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_190
timestamp 1604666999
transform 1 0 18584 0 1 13426
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_194
timestamp 1604666999
transform 1 0 18952 0 1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_198
timestamp 1604666999
transform 1 0 19320 0 1 13426
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 20792 0 1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 19504 0 1 13426
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 19872 0 1 13426
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 20240 0 1 13426
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_202
timestamp 1604666999
transform 1 0 19688 0 1 13426
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1604666999
transform 1 0 20056 0 1 13426
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1604666999
transform 1 0 20424 0 1 13426
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_215
timestamp 1604666999
transform 1 0 20884 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_227
timestamp 1604666999
transform 1 0 21988 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_239
timestamp 1604666999
transform 1 0 23092 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_251
timestamp 1604666999
transform 1 0 24196 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 26404 0 1 13426
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_263
timestamp 1604666999
transform 1 0 25300 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_276
timestamp 1604666999
transform 1 0 26496 0 1 13426
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_288
timestamp 1604666999
transform 1 0 27600 0 1 13426
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_296
timestamp 1604666999
transform 1 0 28336 0 1 13426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 28888 0 1 13426
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604666999
transform 1 0 1380 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604666999
transform 1 0 2484 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_27
timestamp 1604666999
transform 1 0 3588 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_39
timestamp 1604666999
transform 1 0 4692 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_51
timestamp 1604666999
transform 1 0 5796 0 -1 14514
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1604666999
transform 1 0 6532 0 -1 14514
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 6716 0 -1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_62
timestamp 1604666999
transform 1 0 6808 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_74
timestamp 1604666999
transform 1 0 7912 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_86
timestamp 1604666999
transform 1 0 9016 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_98
timestamp 1604666999
transform 1 0 10120 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_110
timestamp 1604666999
transform 1 0 11224 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 12328 0 -1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1604666999
transform 1 0 12420 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_135
timestamp 1604666999
transform 1 0 13524 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_147
timestamp 1604666999
transform 1 0 14628 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_159
timestamp 1604666999
transform 1 0 15732 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_171
timestamp 1604666999
transform 1 0 16836 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 17940 0 -1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 18492 0 -1 14514
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_184
timestamp 1604666999
transform 1 0 18032 0 -1 14514
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_188
timestamp 1604666999
transform 1 0 18400 0 -1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_191
timestamp 1604666999
transform 1 0 18676 0 -1 14514
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 19412 0 -1 14514
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_208
timestamp 1604666999
transform 1 0 20240 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_220
timestamp 1604666999
transform 1 0 21344 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_232
timestamp 1604666999
transform 1 0 22448 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 23552 0 -1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_245
timestamp 1604666999
transform 1 0 23644 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_257
timestamp 1604666999
transform 1 0 24748 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_269
timestamp 1604666999
transform 1 0 25852 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_281
timestamp 1604666999
transform 1 0 26956 0 -1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_293
timestamp 1604666999
transform 1 0 28060 0 -1 14514
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 28888 0 -1 14514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1604666999
transform 1 0 1380 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1604666999
transform 1 0 2484 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 3956 0 1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1604666999
transform 1 0 3588 0 1 14514
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_32
timestamp 1604666999
transform 1 0 4048 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_44
timestamp 1604666999
transform 1 0 5152 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_56
timestamp 1604666999
transform 1 0 6256 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_68
timestamp 1604666999
transform 1 0 7360 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 9568 0 1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_80
timestamp 1604666999
transform 1 0 8464 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1604666999
transform 1 0 9660 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_105
timestamp 1604666999
transform 1 0 10764 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_117
timestamp 1604666999
transform 1 0 11868 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_129
timestamp 1604666999
transform 1 0 12972 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 15180 0 1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_141
timestamp 1604666999
transform 1 0 14076 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1604666999
transform 1 0 15272 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_166
timestamp 1604666999
transform 1 0 16376 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_178
timestamp 1604666999
transform 1 0 17480 0 1 14514
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 18492 0 1 14514
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 18308 0 1 14514
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_186
timestamp 1604666999
transform 1 0 18216 0 1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_198
timestamp 1604666999
transform 1 0 19320 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 20792 0 1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1604666999
transform 1 0 20424 0 1 14514
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_215
timestamp 1604666999
transform 1 0 20884 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_227
timestamp 1604666999
transform 1 0 21988 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1604666999
transform 1 0 23920 0 1 14514
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_239
timestamp 1604666999
transform 1 0 23092 0 1 14514
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_247
timestamp 1604666999
transform 1 0 23828 0 1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_250
timestamp 1604666999
transform 1 0 24104 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 26404 0 1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_262
timestamp 1604666999
transform 1 0 25208 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_274
timestamp 1604666999
transform 1 0 26312 0 1 14514
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_276
timestamp 1604666999
transform 1 0 26496 0 1 14514
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_288
timestamp 1604666999
transform 1 0 27600 0 1 14514
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_296
timestamp 1604666999
transform 1 0 28336 0 1 14514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 28888 0 1 14514
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604666999
transform 1 0 1380 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604666999
transform 1 0 2484 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_27
timestamp 1604666999
transform 1 0 3588 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_39
timestamp 1604666999
transform 1 0 4692 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_51
timestamp 1604666999
transform 1 0 5796 0 -1 15602
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_59
timestamp 1604666999
transform 1 0 6532 0 -1 15602
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 6716 0 -1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 7084 0 -1 15602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_62
timestamp 1604666999
transform 1 0 6808 0 -1 15602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_67
timestamp 1604666999
transform 1 0 7268 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_79
timestamp 1604666999
transform 1 0 8372 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_91
timestamp 1604666999
transform 1 0 9476 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_103
timestamp 1604666999
transform 1 0 10580 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_115
timestamp 1604666999
transform 1 0 11684 0 -1 15602
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 12328 0 -1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_121
timestamp 1604666999
transform 1 0 12236 0 -1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1604666999
transform 1 0 12420 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_135
timestamp 1604666999
transform 1 0 13524 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_147
timestamp 1604666999
transform 1 0 14628 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_159
timestamp 1604666999
transform 1 0 15732 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_171
timestamp 1604666999
transform 1 0 16836 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 17940 0 -1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 18492 0 -1 15602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_184
timestamp 1604666999
transform 1 0 18032 0 -1 15602
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_188
timestamp 1604666999
transform 1 0 18400 0 -1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_191
timestamp 1604666999
transform 1 0 18676 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_203
timestamp 1604666999
transform 1 0 19780 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604666999
transform 1 0 20884 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604666999
transform 1 0 21988 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1604666999
transform 1 0 23920 0 -1 15602
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 23552 0 -1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_239
timestamp 1604666999
transform 1 0 23092 0 -1 15602
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_243
timestamp 1604666999
transform 1 0 23460 0 -1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_245
timestamp 1604666999
transform 1 0 23644 0 -1 15602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_252
timestamp 1604666999
transform 1 0 24288 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_264
timestamp 1604666999
transform 1 0 25392 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_276
timestamp 1604666999
transform 1 0 26496 0 -1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_288
timestamp 1604666999
transform 1 0 27600 0 -1 15602
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_296
timestamp 1604666999
transform 1 0 28336 0 -1 15602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 28888 0 -1 15602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604666999
transform 1 0 1380 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604666999
transform 1 0 2484 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 3956 0 1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_27
timestamp 1604666999
transform 1 0 3588 0 1 15602
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_32
timestamp 1604666999
transform 1 0 4048 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_44
timestamp 1604666999
transform 1 0 5152 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_56
timestamp 1604666999
transform 1 0 6256 0 1 15602
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 7084 0 1 15602
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6900 0 1 15602
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1604666999
transform 1 0 6808 0 1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 9568 0 1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_84
timestamp 1604666999
transform 1 0 8832 0 1 15602
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1604666999
transform 1 0 9660 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_105
timestamp 1604666999
transform 1 0 10764 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_117
timestamp 1604666999
transform 1 0 11868 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 12972 0 1 15602
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13340 0 1 15602
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_131
timestamp 1604666999
transform 1 0 13156 0 1 15602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1604666999
transform 1 0 13524 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 15180 0 1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_147
timestamp 1604666999
transform 1 0 14628 0 1 15602
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_154
timestamp 1604666999
transform 1 0 15272 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_166
timestamp 1604666999
transform 1 0 16376 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_178
timestamp 1604666999
transform 1 0 17480 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_190
timestamp 1604666999
transform 1 0 18584 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 20792 0 1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_202
timestamp 1604666999
transform 1 0 19688 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_215
timestamp 1604666999
transform 1 0 20884 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_227
timestamp 1604666999
transform 1 0 21988 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1604666999
transform 1 0 23920 0 1 15602
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1604666999
transform 1 0 24472 0 1 15602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_239
timestamp 1604666999
transform 1 0 23092 0 1 15602
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_247
timestamp 1604666999
transform 1 0 23828 0 1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_252
timestamp 1604666999
transform 1 0 24288 0 1 15602
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_256
timestamp 1604666999
transform 1 0 24656 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 26404 0 1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_268
timestamp 1604666999
transform 1 0 25760 0 1 15602
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_274
timestamp 1604666999
transform 1 0 26312 0 1 15602
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_276
timestamp 1604666999
transform 1 0 26496 0 1 15602
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_288
timestamp 1604666999
transform 1 0 27600 0 1 15602
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_296
timestamp 1604666999
transform 1 0 28336 0 1 15602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 28888 0 1 15602
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604666999
transform 1 0 1380 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604666999
transform 1 0 2484 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604666999
transform 1 0 1380 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604666999
transform 1 0 2484 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 3956 0 1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_27
timestamp 1604666999
transform 1 0 3588 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_39
timestamp 1604666999
transform 1 0 4692 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1604666999
transform 1 0 3588 0 1 16690
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1604666999
transform 1 0 4048 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_51
timestamp 1604666999
transform 1 0 5796 0 -1 16690
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_59
timestamp 1604666999
transform 1 0 6532 0 -1 16690
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1604666999
transform 1 0 5152 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_56
timestamp 1604666999
transform 1 0 6256 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 6716 0 -1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_62
timestamp 1604666999
transform 1 0 6808 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_74
timestamp 1604666999
transform 1 0 7912 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_68
timestamp 1604666999
transform 1 0 7360 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 9568 0 1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_86
timestamp 1604666999
transform 1 0 9016 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_98
timestamp 1604666999
transform 1 0 10120 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_80
timestamp 1604666999
transform 1 0 8464 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1604666999
transform 1 0 9660 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_110
timestamp 1604666999
transform 1 0 11224 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_105
timestamp 1604666999
transform 1 0 10764 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_117
timestamp 1604666999
transform 1 0 11868 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 12972 0 -1 16690
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 12328 0 -1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_123
timestamp 1604666999
transform 1 0 12420 0 -1 16690
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_129
timestamp 1604666999
transform 1 0 12972 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 15180 0 1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_148
timestamp 1604666999
transform 1 0 14720 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_141
timestamp 1604666999
transform 1 0 14076 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_154
timestamp 1604666999
transform 1 0 15272 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 17480 0 1 16690
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_160
timestamp 1604666999
transform 1 0 15824 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_172
timestamp 1604666999
transform 1 0 16928 0 -1 16690
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_166
timestamp 1604666999
transform 1 0 16376 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 16690
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 17940 0 -1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 17848 0 1 16690
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 18216 0 -1 16690
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_180
timestamp 1604666999
transform 1 0 17664 0 -1 16690
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_184
timestamp 1604666999
transform 1 0 18032 0 -1 16690
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_188
timestamp 1604666999
transform 1 0 18400 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_180
timestamp 1604666999
transform 1 0 17664 0 1 16690
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1604666999
transform 1 0 18860 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 20792 0 1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_200
timestamp 1604666999
transform 1 0 19504 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_212
timestamp 1604666999
transform 1 0 20608 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_205
timestamp 1604666999
transform 1 0 19964 0 1 16690
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_213
timestamp 1604666999
transform 1 0 20700 0 1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_215
timestamp 1604666999
transform 1 0 20884 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_224
timestamp 1604666999
transform 1 0 21712 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_236
timestamp 1604666999
transform 1 0 22816 0 -1 16690
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_227
timestamp 1604666999
transform 1 0 21988 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 23552 0 -1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1604666999
transform 1 0 23920 0 1 16690
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_245
timestamp 1604666999
transform 1 0 23644 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_257
timestamp 1604666999
transform 1 0 24748 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_239
timestamp 1604666999
transform 1 0 23092 0 1 16690
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_247
timestamp 1604666999
transform 1 0 23828 0 1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_250
timestamp 1604666999
transform 1 0 24104 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 26404 0 1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_269
timestamp 1604666999
transform 1 0 25852 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_262
timestamp 1604666999
transform 1 0 25208 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_274
timestamp 1604666999
transform 1 0 26312 0 1 16690
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_276
timestamp 1604666999
transform 1 0 26496 0 1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_281
timestamp 1604666999
transform 1 0 26956 0 -1 16690
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_293
timestamp 1604666999
transform 1 0 28060 0 -1 16690
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_288
timestamp 1604666999
transform 1 0 27600 0 1 16690
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_296
timestamp 1604666999
transform 1 0 28336 0 1 16690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 28888 0 -1 16690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 28888 0 1 16690
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604666999
transform 1 0 1380 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604666999
transform 1 0 2484 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_27
timestamp 1604666999
transform 1 0 3588 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_39
timestamp 1604666999
transform 1 0 4692 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_51
timestamp 1604666999
transform 1 0 5796 0 -1 17778
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_59
timestamp 1604666999
transform 1 0 6532 0 -1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 6716 0 -1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_62
timestamp 1604666999
transform 1 0 6808 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_74
timestamp 1604666999
transform 1 0 7912 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_86
timestamp 1604666999
transform 1 0 9016 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_98
timestamp 1604666999
transform 1 0 10120 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_110
timestamp 1604666999
transform 1 0 11224 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 12328 0 -1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1604666999
transform 1 0 12420 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_135
timestamp 1604666999
transform 1 0 13524 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_147
timestamp 1604666999
transform 1 0 14628 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_159
timestamp 1604666999
transform 1 0 15732 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_171
timestamp 1604666999
transform 1 0 16836 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 17940 0 -1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_184
timestamp 1604666999
transform 1 0 18032 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_196
timestamp 1604666999
transform 1 0 19136 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_208
timestamp 1604666999
transform 1 0 20240 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_220
timestamp 1604666999
transform 1 0 21344 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_232
timestamp 1604666999
transform 1 0 22448 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1604666999
transform 1 0 23920 0 -1 17778
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 23552 0 -1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_245
timestamp 1604666999
transform 1 0 23644 0 -1 17778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_252
timestamp 1604666999
transform 1 0 24288 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_264
timestamp 1604666999
transform 1 0 25392 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1604666999
transform 1 0 26496 0 -1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_288
timestamp 1604666999
transform 1 0 27600 0 -1 17778
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1604666999
transform 1 0 28336 0 -1 17778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 28888 0 -1 17778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604666999
transform 1 0 1380 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604666999
transform 1 0 2484 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 3956 0 1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1604666999
transform 1 0 3588 0 1 17778
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1604666999
transform 1 0 4048 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1604666999
transform 1 0 5152 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_56
timestamp 1604666999
transform 1 0 6256 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_68
timestamp 1604666999
transform 1 0 7360 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 9568 0 1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 8556 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 8924 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_80
timestamp 1604666999
transform 1 0 8464 0 1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_83
timestamp 1604666999
transform 1 0 8740 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_87
timestamp 1604666999
transform 1 0 9108 0 1 17778
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_91
timestamp 1604666999
transform 1 0 9476 0 1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1604666999
transform 1 0 9660 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_105
timestamp 1604666999
transform 1 0 10764 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_117
timestamp 1604666999
transform 1 0 11868 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_129
timestamp 1604666999
transform 1 0 12972 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 15180 0 1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 15456 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_141
timestamp 1604666999
transform 1 0 14076 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_154
timestamp 1604666999
transform 1 0 15272 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_158
timestamp 1604666999
transform 1 0 15640 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 15824 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_162
timestamp 1604666999
transform 1 0 16008 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_174
timestamp 1604666999
transform 1 0 17112 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_186
timestamp 1604666999
transform 1 0 18216 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_198
timestamp 1604666999
transform 1 0 19320 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 20792 0 1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 20424 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_212
timestamp 1604666999
transform 1 0 20608 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_215
timestamp 1604666999
transform 1 0 20884 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_227
timestamp 1604666999
transform 1 0 21988 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604666999
transform 1 0 23920 0 1 17778
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604666999
transform 1 0 24472 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604666999
transform 1 0 23736 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_239
timestamp 1604666999
transform 1 0 23092 0 1 17778
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_245
timestamp 1604666999
transform 1 0 23644 0 1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_252
timestamp 1604666999
transform 1 0 24288 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_256
timestamp 1604666999
transform 1 0 24656 0 1 17778
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 26404 0 1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__17__A
timestamp 1604666999
transform 1 0 25024 0 1 17778
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_262
timestamp 1604666999
transform 1 0 25208 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_274
timestamp 1604666999
transform 1 0 26312 0 1 17778
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_276
timestamp 1604666999
transform 1 0 26496 0 1 17778
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_288
timestamp 1604666999
transform 1 0 27600 0 1 17778
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_296
timestamp 1604666999
transform 1 0 28336 0 1 17778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 28888 0 1 17778
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 18866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604666999
transform 1 0 1380 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604666999
transform 1 0 2484 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_27
timestamp 1604666999
transform 1 0 3588 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_39
timestamp 1604666999
transform 1 0 4692 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_51
timestamp 1604666999
transform 1 0 5796 0 -1 18866
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1604666999
transform 1 0 6532 0 -1 18866
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 6716 0 -1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_62
timestamp 1604666999
transform 1 0 6808 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_74
timestamp 1604666999
transform 1 0 7912 0 -1 18866
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8556 0 -1 18866
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_30_80
timestamp 1604666999
transform 1 0 8464 0 -1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_100
timestamp 1604666999
transform 1 0 10304 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_112
timestamp 1604666999
transform 1 0 11408 0 -1 18866
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 12328 0 -1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1604666999
transform 1 0 12144 0 -1 18866
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_123
timestamp 1604666999
transform 1 0 12420 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_135
timestamp 1604666999
transform 1 0 13524 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 15272 0 -1 18866
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_30_147
timestamp 1604666999
transform 1 0 14628 0 -1 18866
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_153
timestamp 1604666999
transform 1 0 15180 0 -1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_173
timestamp 1604666999
transform 1 0 17020 0 -1 18866
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 17940 0 -1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_181
timestamp 1604666999
transform 1 0 17756 0 -1 18866
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_184
timestamp 1604666999
transform 1 0 18032 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_196
timestamp 1604666999
transform 1 0 19136 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 20424 0 -1 18866
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_208
timestamp 1604666999
transform 1 0 20240 0 -1 18866
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_213
timestamp 1604666999
transform 1 0 20700 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_225
timestamp 1604666999
transform 1 0 21804 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_237
timestamp 1604666999
transform 1 0 22908 0 -1 18866
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604666999
transform 1 0 23920 0 -1 18866
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 23552 0 -1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_243
timestamp 1604666999
transform 1 0 23460 0 -1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_245
timestamp 1604666999
transform 1 0 23644 0 -1 18866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_252
timestamp 1604666999
transform 1 0 24288 0 -1 18866
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1604666999
transform 1 0 25024 0 -1 18866
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_264
timestamp 1604666999
transform 1 0 25392 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1604666999
transform 1 0 26496 0 -1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_288
timestamp 1604666999
transform 1 0 27600 0 -1 18866
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_296
timestamp 1604666999
transform 1 0 28336 0 -1 18866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 28888 0 -1 18866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 18866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604666999
transform 1 0 1380 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604666999
transform 1 0 2484 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 3956 0 1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_27
timestamp 1604666999
transform 1 0 3588 0 1 18866
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_32
timestamp 1604666999
transform 1 0 4048 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_44
timestamp 1604666999
transform 1 0 5152 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_56
timestamp 1604666999
transform 1 0 6256 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_68
timestamp 1604666999
transform 1 0 7360 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 9568 0 1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_80
timestamp 1604666999
transform 1 0 8464 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1604666999
transform 1 0 9660 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_105
timestamp 1604666999
transform 1 0 10764 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_117
timestamp 1604666999
transform 1 0 11868 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_129
timestamp 1604666999
transform 1 0 12972 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 15180 0 1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_141
timestamp 1604666999
transform 1 0 14076 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_154
timestamp 1604666999
transform 1 0 15272 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_166
timestamp 1604666999
transform 1 0 16376 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_178
timestamp 1604666999
transform 1 0 17480 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_190
timestamp 1604666999
transform 1 0 18584 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 20792 0 1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_202
timestamp 1604666999
transform 1 0 19688 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_215
timestamp 1604666999
transform 1 0 20884 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_227
timestamp 1604666999
transform 1 0 21988 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604666999
transform 1 0 23920 0 1 18866
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604666999
transform 1 0 24472 0 1 18866
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_239
timestamp 1604666999
transform 1 0 23092 0 1 18866
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_247
timestamp 1604666999
transform 1 0 23828 0 1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_252
timestamp 1604666999
transform 1 0 24288 0 1 18866
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_256
timestamp 1604666999
transform 1 0 24656 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 26404 0 1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_268
timestamp 1604666999
transform 1 0 25760 0 1 18866
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_274
timestamp 1604666999
transform 1 0 26312 0 1 18866
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_276
timestamp 1604666999
transform 1 0 26496 0 1 18866
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_288
timestamp 1604666999
transform 1 0 27600 0 1 18866
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_296
timestamp 1604666999
transform 1 0 28336 0 1 18866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 28888 0 1 18866
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 19954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604666999
transform 1 0 1380 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604666999
transform 1 0 2484 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_27
timestamp 1604666999
transform 1 0 3588 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_39
timestamp 1604666999
transform 1 0 4692 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_51
timestamp 1604666999
transform 1 0 5796 0 -1 19954
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_59
timestamp 1604666999
transform 1 0 6532 0 -1 19954
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 6716 0 -1 19954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_62
timestamp 1604666999
transform 1 0 6808 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_74
timestamp 1604666999
transform 1 0 7912 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_86
timestamp 1604666999
transform 1 0 9016 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_98
timestamp 1604666999
transform 1 0 10120 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_110
timestamp 1604666999
transform 1 0 11224 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 12328 0 -1 19954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1604666999
transform 1 0 12420 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_135
timestamp 1604666999
transform 1 0 13524 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_147
timestamp 1604666999
transform 1 0 14628 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_159
timestamp 1604666999
transform 1 0 15732 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_171
timestamp 1604666999
transform 1 0 16836 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 17940 0 -1 19954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_184
timestamp 1604666999
transform 1 0 18032 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_196
timestamp 1604666999
transform 1 0 19136 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_208
timestamp 1604666999
transform 1 0 20240 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_220
timestamp 1604666999
transform 1 0 21344 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_232
timestamp 1604666999
transform 1 0 22448 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 23552 0 -1 19954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_245
timestamp 1604666999
transform 1 0 23644 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_257
timestamp 1604666999
transform 1 0 24748 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_269
timestamp 1604666999
transform 1 0 25852 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_281
timestamp 1604666999
transform 1 0 26956 0 -1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_293
timestamp 1604666999
transform 1 0 28060 0 -1 19954
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 28888 0 -1 19954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 19954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604666999
transform 1 0 1380 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604666999
transform 1 0 2484 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604666999
transform 1 0 1380 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604666999
transform 1 0 2484 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 3956 0 1 19954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_27
timestamp 1604666999
transform 1 0 3588 0 1 19954
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1604666999
transform 1 0 4048 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_27
timestamp 1604666999
transform 1 0 3588 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_39
timestamp 1604666999
transform 1 0 4692 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1604666999
transform 1 0 5152 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_56
timestamp 1604666999
transform 1 0 6256 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_51
timestamp 1604666999
transform 1 0 5796 0 -1 21042
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_59
timestamp 1604666999
transform 1 0 6532 0 -1 21042
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 6716 0 -1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_68
timestamp 1604666999
transform 1 0 7360 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_62
timestamp 1604666999
transform 1 0 6808 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_74
timestamp 1604666999
transform 1 0 7912 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 9568 0 1 19954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_80
timestamp 1604666999
transform 1 0 8464 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1604666999
transform 1 0 9660 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_86
timestamp 1604666999
transform 1 0 9016 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_98
timestamp 1604666999
transform 1 0 10120 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_105
timestamp 1604666999
transform 1 0 10764 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_117
timestamp 1604666999
transform 1 0 11868 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_110
timestamp 1604666999
transform 1 0 11224 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 12328 0 -1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_129
timestamp 1604666999
transform 1 0 12972 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1604666999
transform 1 0 12420 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_135
timestamp 1604666999
transform 1 0 13524 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 15180 0 1 19954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_141
timestamp 1604666999
transform 1 0 14076 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_154
timestamp 1604666999
transform 1 0 15272 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_147
timestamp 1604666999
transform 1 0 14628 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_166
timestamp 1604666999
transform 1 0 16376 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_178
timestamp 1604666999
transform 1 0 17480 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_159
timestamp 1604666999
transform 1 0 15732 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_171
timestamp 1604666999
transform 1 0 16836 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 17940 0 -1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_190
timestamp 1604666999
transform 1 0 18584 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_184
timestamp 1604666999
transform 1 0 18032 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_196
timestamp 1604666999
transform 1 0 19136 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 20792 0 1 19954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_202
timestamp 1604666999
transform 1 0 19688 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_215
timestamp 1604666999
transform 1 0 20884 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_208
timestamp 1604666999
transform 1 0 20240 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_227
timestamp 1604666999
transform 1 0 21988 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_220
timestamp 1604666999
transform 1 0 21344 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_232
timestamp 1604666999
transform 1 0 22448 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 23552 0 -1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_239
timestamp 1604666999
transform 1 0 23092 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_251
timestamp 1604666999
transform 1 0 24196 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_245
timestamp 1604666999
transform 1 0 23644 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_257
timestamp 1604666999
transform 1 0 24748 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 26404 0 1 19954
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_263
timestamp 1604666999
transform 1 0 25300 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_276
timestamp 1604666999
transform 1 0 26496 0 1 19954
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_269
timestamp 1604666999
transform 1 0 25852 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_288
timestamp 1604666999
transform 1 0 27600 0 1 19954
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_296
timestamp 1604666999
transform 1 0 28336 0 1 19954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_281
timestamp 1604666999
transform 1 0 26956 0 -1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_293
timestamp 1604666999
transform 1 0 28060 0 -1 21042
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 28888 0 1 19954
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 28888 0 -1 21042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21042
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604666999
transform 1 0 1380 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604666999
transform 1 0 2484 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 3956 0 1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604666999
transform 1 0 3588 0 1 21042
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604666999
transform 1 0 4048 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604666999
transform 1 0 5152 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604666999
transform 1 0 6256 0 1 21042
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 6808 0 1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604666999
transform 1 0 6900 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604666999
transform 1 0 8004 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 9660 0 1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604666999
transform 1 0 9108 0 1 21042
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604666999
transform 1 0 9752 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604666999
transform 1 0 10856 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604666999
transform 1 0 11960 0 1 21042
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 12512 0 1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604666999
transform 1 0 12604 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604666999
transform 1 0 13708 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 15364 0 1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604666999
transform 1 0 14812 0 1 21042
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604666999
transform 1 0 15456 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604666999
transform 1 0 16560 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 18216 0 1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604666999
transform 1 0 17664 0 1 21042
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604666999
transform 1 0 18308 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 21068 0 1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604666999
transform 1 0 19412 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604666999
transform 1 0 20516 0 1 21042
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604666999
transform 1 0 21160 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604666999
transform 1 0 22264 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 23920 0 1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604666999
transform 1 0 23368 0 1 21042
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604666999
transform 1 0 24012 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604666999
transform 1 0 25116 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604666999
transform 1 0 26220 0 1 21042
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 26772 0 1 21042
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604666999
transform 1 0 26864 0 1 21042
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604666999
transform 1 0 27968 0 1 21042
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 28888 0 1 21042
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604666999
transform 1 0 28520 0 1 21042
box -38 -48 130 592
<< labels >>
rlabel metal2 s 11150 23346 11206 23826 6 ccff_head
port 0 nsew default input
rlabel metal2 s 18694 23346 18750 23826 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 12074 480 12194 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 18058 480 18178 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 18602 480 18722 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 19146 480 19266 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 19826 480 19946 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 20370 480 20490 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 21050 480 21170 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 21594 480 21714 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 22138 480 22258 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 22818 480 22938 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 23362 480 23482 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 12618 480 12738 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 13162 480 13282 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 13842 480 13962 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 14386 480 14506 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 15066 480 15186 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 15610 480 15730 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 16154 480 16274 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 16834 480 16954 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 17378 480 17498 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 106 480 226 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 6090 480 6210 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 6634 480 6754 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 7178 480 7298 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 7858 480 7978 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 8402 480 8522 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 9082 480 9202 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 9626 480 9746 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 10170 480 10290 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 10850 480 10970 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 11394 480 11514 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 650 480 770 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 1194 480 1314 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 1874 480 1994 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 2418 480 2538 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 3098 480 3218 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 3642 480 3762 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 4186 480 4306 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 4866 480 4986 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 5410 480 5530 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal3 s 29520 12074 30000 12194 6 chanx_right_in[0]
port 42 nsew default input
rlabel metal3 s 29520 18058 30000 18178 6 chanx_right_in[10]
port 43 nsew default input
rlabel metal3 s 29520 18602 30000 18722 6 chanx_right_in[11]
port 44 nsew default input
rlabel metal3 s 29520 19146 30000 19266 6 chanx_right_in[12]
port 45 nsew default input
rlabel metal3 s 29520 19826 30000 19946 6 chanx_right_in[13]
port 46 nsew default input
rlabel metal3 s 29520 20370 30000 20490 6 chanx_right_in[14]
port 47 nsew default input
rlabel metal3 s 29520 21050 30000 21170 6 chanx_right_in[15]
port 48 nsew default input
rlabel metal3 s 29520 21594 30000 21714 6 chanx_right_in[16]
port 49 nsew default input
rlabel metal3 s 29520 22138 30000 22258 6 chanx_right_in[17]
port 50 nsew default input
rlabel metal3 s 29520 22818 30000 22938 6 chanx_right_in[18]
port 51 nsew default input
rlabel metal3 s 29520 23362 30000 23482 6 chanx_right_in[19]
port 52 nsew default input
rlabel metal3 s 29520 12618 30000 12738 6 chanx_right_in[1]
port 53 nsew default input
rlabel metal3 s 29520 13162 30000 13282 6 chanx_right_in[2]
port 54 nsew default input
rlabel metal3 s 29520 13842 30000 13962 6 chanx_right_in[3]
port 55 nsew default input
rlabel metal3 s 29520 14386 30000 14506 6 chanx_right_in[4]
port 56 nsew default input
rlabel metal3 s 29520 15066 30000 15186 6 chanx_right_in[5]
port 57 nsew default input
rlabel metal3 s 29520 15610 30000 15730 6 chanx_right_in[6]
port 58 nsew default input
rlabel metal3 s 29520 16154 30000 16274 6 chanx_right_in[7]
port 59 nsew default input
rlabel metal3 s 29520 16834 30000 16954 6 chanx_right_in[8]
port 60 nsew default input
rlabel metal3 s 29520 17378 30000 17498 6 chanx_right_in[9]
port 61 nsew default input
rlabel metal3 s 29520 106 30000 226 6 chanx_right_out[0]
port 62 nsew default tristate
rlabel metal3 s 29520 6090 30000 6210 6 chanx_right_out[10]
port 63 nsew default tristate
rlabel metal3 s 29520 6634 30000 6754 6 chanx_right_out[11]
port 64 nsew default tristate
rlabel metal3 s 29520 7178 30000 7298 6 chanx_right_out[12]
port 65 nsew default tristate
rlabel metal3 s 29520 7858 30000 7978 6 chanx_right_out[13]
port 66 nsew default tristate
rlabel metal3 s 29520 8402 30000 8522 6 chanx_right_out[14]
port 67 nsew default tristate
rlabel metal3 s 29520 9082 30000 9202 6 chanx_right_out[15]
port 68 nsew default tristate
rlabel metal3 s 29520 9626 30000 9746 6 chanx_right_out[16]
port 69 nsew default tristate
rlabel metal3 s 29520 10170 30000 10290 6 chanx_right_out[17]
port 70 nsew default tristate
rlabel metal3 s 29520 10850 30000 10970 6 chanx_right_out[18]
port 71 nsew default tristate
rlabel metal3 s 29520 11394 30000 11514 6 chanx_right_out[19]
port 72 nsew default tristate
rlabel metal3 s 29520 650 30000 770 6 chanx_right_out[1]
port 73 nsew default tristate
rlabel metal3 s 29520 1194 30000 1314 6 chanx_right_out[2]
port 74 nsew default tristate
rlabel metal3 s 29520 1874 30000 1994 6 chanx_right_out[3]
port 75 nsew default tristate
rlabel metal3 s 29520 2418 30000 2538 6 chanx_right_out[4]
port 76 nsew default tristate
rlabel metal3 s 29520 3098 30000 3218 6 chanx_right_out[5]
port 77 nsew default tristate
rlabel metal3 s 29520 3642 30000 3762 6 chanx_right_out[6]
port 78 nsew default tristate
rlabel metal3 s 29520 4186 30000 4306 6 chanx_right_out[7]
port 79 nsew default tristate
rlabel metal3 s 29520 4866 30000 4986 6 chanx_right_out[8]
port 80 nsew default tristate
rlabel metal3 s 29520 5410 30000 5530 6 chanx_right_out[9]
port 81 nsew default tristate
rlabel metal2 s 3698 23346 3754 23826 6 prog_clk
port 82 nsew default input
rlabel metal2 s 26146 23346 26202 23826 6 top_grid_pin_0_
port 83 nsew default tristate
rlabel metal4 s 5944 1954 6264 21634 6 VPWR
port 84 nsew default input
rlabel metal4 s 10944 1954 11264 21634 6 VGND
port 85 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 23826
<< end >>
