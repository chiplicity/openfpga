magic
tech EFS8A
magscale 1 2
timestamp 1602529361
<< locali >>
rect 11471 25313 11506 25347
rect 10183 24225 10310 24259
rect 6135 22049 6170 22083
rect 11339 21097 11345 21131
rect 16491 21097 16497 21131
rect 11339 21029 11373 21097
rect 16491 21029 16525 21097
rect 9631 20961 9758 20995
rect 16399 20009 16405 20043
rect 16399 19941 16433 20009
rect 19751 19873 19786 19907
rect 13553 19159 13587 19329
rect 16583 18921 16589 18955
rect 3111 18853 3249 18887
rect 16583 18853 16617 18921
rect 2915 18785 3042 18819
rect 3795 18071 3829 18139
rect 7843 18071 7877 18139
rect 15111 18071 15145 18139
rect 3795 18037 3801 18071
rect 7843 18037 7849 18071
rect 15111 18037 15117 18071
rect 7751 17833 7757 17867
rect 7751 17765 7785 17833
rect 19199 17697 19234 17731
rect 6975 17289 7113 17323
rect 19947 17289 20085 17323
rect 4905 17051 4939 17221
rect 6779 17085 6906 17119
rect 10143 16745 10149 16779
rect 16767 16745 16773 16779
rect 10143 16677 10177 16745
rect 16767 16677 16801 16745
rect 15243 16609 15370 16643
rect 24535 16609 24662 16643
rect 6929 16031 6963 16065
rect 6929 15997 7090 16031
rect 16215 15657 16221 15691
rect 16215 15589 16249 15657
rect 19475 15521 19510 15555
rect 10241 14807 10275 15113
rect 10879 14807 10913 14875
rect 10879 14773 10885 14807
rect 20855 14433 20982 14467
rect 9965 13855 9999 13957
rect 17359 13345 17394 13379
rect 18245 13175 18279 13277
rect 10787 12631 10821 12699
rect 10787 12597 10793 12631
rect 7021 12087 7055 12393
rect 10787 11543 10821 11611
rect 10787 11509 10793 11543
rect 5451 11305 5457 11339
rect 5451 11237 5485 11305
rect 4537 10455 4571 10761
rect 15939 10217 15945 10251
rect 17687 10217 17693 10251
rect 15939 10149 15973 10217
rect 17687 10149 17721 10217
rect 9413 9435 9447 9537
rect 18739 8993 18774 9027
rect 14231 7905 14266 7939
rect 1443 6817 1478 6851
rect 8619 4641 8654 4675
rect 9355 4029 9390 4063
<< viali >>
rect 11437 25313 11471 25347
rect 13252 25313 13286 25347
rect 14264 25313 14298 25347
rect 10425 25245 10459 25279
rect 14335 25177 14369 25211
rect 11575 25109 11609 25143
rect 13323 25109 13357 25143
rect 10793 24905 10827 24939
rect 11069 24905 11103 24939
rect 14565 24905 14599 24939
rect 14933 24905 14967 24939
rect 10425 24837 10459 24871
rect 11897 24769 11931 24803
rect 13553 24769 13587 24803
rect 8928 24701 8962 24735
rect 9924 24701 9958 24735
rect 10885 24701 10919 24735
rect 11529 24701 11563 24735
rect 12725 24701 12759 24735
rect 12909 24701 12943 24735
rect 14080 24701 14114 24735
rect 10011 24633 10045 24667
rect 8999 24565 9033 24599
rect 9321 24565 9355 24599
rect 12173 24565 12207 24599
rect 12725 24565 12759 24599
rect 14151 24565 14185 24599
rect 9873 24361 9907 24395
rect 11437 24361 11471 24395
rect 14289 24361 14323 24395
rect 12633 24293 12667 24327
rect 12725 24293 12759 24327
rect 1444 24225 1478 24259
rect 8620 24225 8654 24259
rect 10149 24225 10183 24259
rect 14105 24225 14139 24259
rect 10793 24157 10827 24191
rect 12909 24157 12943 24191
rect 1547 24089 1581 24123
rect 10379 24089 10413 24123
rect 12357 24089 12391 24123
rect 8723 24021 8757 24055
rect 1869 23817 1903 23851
rect 8953 23817 8987 23851
rect 9873 23817 9907 23851
rect 10333 23817 10367 23851
rect 15761 23817 15795 23851
rect 16865 23817 16899 23851
rect 18705 23817 18739 23851
rect 21373 23817 21407 23851
rect 7205 23749 7239 23783
rect 11437 23749 11471 23783
rect 13553 23749 13587 23783
rect 13921 23749 13955 23783
rect 20269 23749 20303 23783
rect 10885 23681 10919 23715
rect 12541 23681 12575 23715
rect 14105 23681 14139 23715
rect 14381 23681 14415 23715
rect 1444 23613 1478 23647
rect 2237 23613 2271 23647
rect 2472 23613 2506 23647
rect 2881 23613 2915 23647
rect 3500 23613 3534 23647
rect 3893 23613 3927 23647
rect 4664 23613 4698 23647
rect 5089 23613 5123 23647
rect 7021 23613 7055 23647
rect 7573 23613 7607 23647
rect 8560 23613 8594 23647
rect 9413 23613 9447 23647
rect 9689 23613 9723 23647
rect 15577 23613 15611 23647
rect 16129 23613 16163 23647
rect 16681 23613 16715 23647
rect 17233 23613 17267 23647
rect 18521 23613 18555 23647
rect 19073 23613 19107 23647
rect 20085 23613 20119 23647
rect 20637 23613 20671 23647
rect 21189 23613 21223 23647
rect 2559 23545 2593 23579
rect 10977 23545 11011 23579
rect 11897 23545 11931 23579
rect 12633 23545 12667 23579
rect 13185 23545 13219 23579
rect 14197 23545 14231 23579
rect 21741 23545 21775 23579
rect 1547 23477 1581 23511
rect 3571 23477 3605 23511
rect 4767 23477 4801 23511
rect 8631 23477 8665 23511
rect 10701 23477 10735 23511
rect 12265 23477 12299 23511
rect 5319 23273 5353 23307
rect 7205 23273 7239 23307
rect 14105 23273 14139 23307
rect 14381 23273 14415 23307
rect 15439 23273 15473 23307
rect 6377 23205 6411 23239
rect 11345 23205 11379 23239
rect 11437 23205 11471 23239
rect 12909 23205 12943 23239
rect 13001 23205 13035 23239
rect 5216 23137 5250 23171
rect 8620 23137 8654 23171
rect 9781 23137 9815 23171
rect 10149 23137 10183 23171
rect 15368 23137 15402 23171
rect 6285 23069 6319 23103
rect 6929 23069 6963 23103
rect 10425 23069 10459 23103
rect 11989 23069 12023 23103
rect 13185 23069 13219 23103
rect 11069 23001 11103 23035
rect 8723 22933 8757 22967
rect 10793 22933 10827 22967
rect 12541 22933 12575 22967
rect 5641 22729 5675 22763
rect 6561 22729 6595 22763
rect 8493 22729 8527 22763
rect 11345 22729 11379 22763
rect 11621 22729 11655 22763
rect 12633 22729 12667 22763
rect 13369 22729 13403 22763
rect 16129 22729 16163 22763
rect 18705 22729 18739 22763
rect 6193 22661 6227 22695
rect 9781 22661 9815 22695
rect 14197 22661 14231 22695
rect 6929 22593 6963 22627
rect 7205 22593 7239 22627
rect 10333 22593 10367 22627
rect 13645 22593 13679 22627
rect 5800 22525 5834 22559
rect 8677 22525 8711 22559
rect 9229 22525 9263 22559
rect 12449 22525 12483 22559
rect 13001 22525 13035 22559
rect 15117 22525 15151 22559
rect 15577 22525 15611 22559
rect 18521 22525 18555 22559
rect 7021 22457 7055 22491
rect 8217 22457 8251 22491
rect 9413 22457 9447 22491
rect 10425 22457 10459 22491
rect 10977 22457 11011 22491
rect 13737 22457 13771 22491
rect 5181 22389 5215 22423
rect 5871 22389 5905 22423
rect 10057 22389 10091 22423
rect 14565 22389 14599 22423
rect 14933 22389 14967 22423
rect 15393 22389 15427 22423
rect 19165 22389 19199 22423
rect 6837 22185 6871 22219
rect 11897 22185 11931 22219
rect 12909 22185 12943 22219
rect 14381 22185 14415 22219
rect 19303 22185 19337 22219
rect 7297 22117 7331 22151
rect 10425 22117 10459 22151
rect 10977 22117 11011 22151
rect 13461 22117 13495 22151
rect 13553 22117 13587 22151
rect 14105 22117 14139 22151
rect 17785 22117 17819 22151
rect 2088 22049 2122 22083
rect 5156 22049 5190 22083
rect 6101 22049 6135 22083
rect 11805 22049 11839 22083
rect 12265 22049 12299 22083
rect 13277 22049 13311 22083
rect 15577 22049 15611 22083
rect 15853 22049 15887 22083
rect 18337 22049 18371 22083
rect 19200 22049 19234 22083
rect 7205 21981 7239 22015
rect 7849 21981 7883 22015
rect 10333 21981 10367 22015
rect 16037 21981 16071 22015
rect 17693 21981 17727 22015
rect 8677 21913 8711 21947
rect 2191 21845 2225 21879
rect 4353 21845 4387 21879
rect 5227 21845 5261 21879
rect 6239 21845 6273 21879
rect 16497 21845 16531 21879
rect 2053 21641 2087 21675
rect 5825 21641 5859 21675
rect 7757 21641 7791 21675
rect 8401 21641 8435 21675
rect 9781 21641 9815 21675
rect 11161 21641 11195 21675
rect 12725 21641 12759 21675
rect 14197 21641 14231 21675
rect 16221 21641 16255 21675
rect 20177 21641 20211 21675
rect 24225 21641 24259 21675
rect 5365 21573 5399 21607
rect 4353 21505 4387 21539
rect 8677 21505 8711 21539
rect 8953 21505 8987 21539
rect 12173 21505 12207 21539
rect 13277 21505 13311 21539
rect 13921 21505 13955 21539
rect 6837 21437 6871 21471
rect 10241 21437 10275 21471
rect 14933 21437 14967 21471
rect 15301 21437 15335 21471
rect 16405 21437 16439 21471
rect 16865 21437 16899 21471
rect 19692 21437 19726 21471
rect 23740 21437 23774 21471
rect 4445 21369 4479 21403
rect 4997 21369 5031 21403
rect 6653 21369 6687 21403
rect 7199 21369 7233 21403
rect 8125 21369 8159 21403
rect 8769 21369 8803 21403
rect 10562 21369 10596 21403
rect 13369 21369 13403 21403
rect 15577 21369 15611 21403
rect 15945 21369 15979 21403
rect 18153 21369 18187 21403
rect 18245 21369 18279 21403
rect 18797 21369 18831 21403
rect 19257 21369 19291 21403
rect 4077 21301 4111 21335
rect 6101 21301 6135 21335
rect 10149 21301 10183 21335
rect 11805 21301 11839 21335
rect 13093 21301 13127 21335
rect 14657 21301 14691 21335
rect 16497 21301 16531 21335
rect 17417 21301 17451 21335
rect 17785 21301 17819 21335
rect 19763 21301 19797 21335
rect 23811 21301 23845 21335
rect 1593 21097 1627 21131
rect 6929 21097 6963 21131
rect 7205 21097 7239 21131
rect 8861 21097 8895 21131
rect 9827 21097 9861 21131
rect 10701 21097 10735 21131
rect 11345 21097 11379 21131
rect 11897 21097 11931 21131
rect 14013 21097 14047 21131
rect 14933 21097 14967 21131
rect 15577 21097 15611 21131
rect 16037 21097 16071 21131
rect 16497 21097 16531 21131
rect 17049 21097 17083 21131
rect 19717 21097 19751 21131
rect 4261 21029 4295 21063
rect 6371 21029 6405 21063
rect 7757 21029 7791 21063
rect 7941 21029 7975 21063
rect 8033 21029 8067 21063
rect 13414 21029 13448 21063
rect 17693 21029 17727 21063
rect 18889 21029 18923 21063
rect 1409 20961 1443 20995
rect 9597 20961 9631 20995
rect 10977 20961 11011 20995
rect 13001 20961 13035 20995
rect 16129 20961 16163 20995
rect 2973 20893 3007 20927
rect 4169 20893 4203 20927
rect 4445 20893 4479 20927
rect 6009 20893 6043 20927
rect 8217 20893 8251 20927
rect 13093 20893 13127 20927
rect 18797 20893 18831 20927
rect 18521 20825 18555 20859
rect 19349 20825 19383 20859
rect 5089 20757 5123 20791
rect 10241 20757 10275 20791
rect 18153 20757 18187 20791
rect 2605 20553 2639 20587
rect 4261 20553 4295 20587
rect 4537 20553 4571 20587
rect 6101 20553 6135 20587
rect 6653 20553 6687 20587
rect 9689 20553 9723 20587
rect 11161 20553 11195 20587
rect 11897 20553 11931 20587
rect 13829 20553 13863 20587
rect 14105 20553 14139 20587
rect 25145 20485 25179 20519
rect 3249 20417 3283 20451
rect 3893 20417 3927 20451
rect 4813 20417 4847 20451
rect 5089 20417 5123 20451
rect 7021 20417 7055 20451
rect 7665 20417 7699 20451
rect 10241 20417 10275 20451
rect 12909 20417 12943 20451
rect 16129 20417 16163 20451
rect 17325 20417 17359 20451
rect 18429 20417 18463 20451
rect 19717 20417 19751 20451
rect 8401 20349 8435 20383
rect 8769 20349 8803 20383
rect 8953 20349 8987 20383
rect 14724 20349 14758 20383
rect 15117 20349 15151 20383
rect 24660 20349 24694 20383
rect 3341 20281 3375 20315
rect 4905 20281 4939 20315
rect 7113 20281 7147 20315
rect 10562 20281 10596 20315
rect 11437 20281 11471 20315
rect 12173 20281 12207 20315
rect 12725 20281 12759 20315
rect 13230 20281 13264 20315
rect 15577 20281 15611 20315
rect 15945 20281 15979 20315
rect 16450 20281 16484 20315
rect 18153 20281 18187 20315
rect 18245 20281 18279 20315
rect 19441 20281 19475 20315
rect 19809 20281 19843 20315
rect 20361 20281 20395 20315
rect 1685 20213 1719 20247
rect 2973 20213 3007 20247
rect 7941 20213 7975 20247
rect 8585 20213 8619 20247
rect 10057 20213 10091 20247
rect 14795 20213 14829 20247
rect 17049 20213 17083 20247
rect 17785 20213 17819 20247
rect 19073 20213 19107 20247
rect 24731 20213 24765 20247
rect 3801 20009 3835 20043
rect 6101 20009 6135 20043
rect 6837 20009 6871 20043
rect 7757 20009 7791 20043
rect 10701 20009 10735 20043
rect 13645 20009 13679 20043
rect 14013 20009 14047 20043
rect 16405 20009 16439 20043
rect 16957 20009 16991 20043
rect 19855 20009 19889 20043
rect 3157 19941 3191 19975
rect 4353 19941 4387 19975
rect 4905 19941 4939 19975
rect 7205 19941 7239 19975
rect 8211 19941 8245 19975
rect 11161 19941 11195 19975
rect 13087 19941 13121 19975
rect 18337 19941 18371 19975
rect 18889 19941 18923 19975
rect 19257 19941 19291 19975
rect 2973 19873 3007 19907
rect 6101 19873 6135 19907
rect 6377 19873 6411 19907
rect 9816 19873 9850 19907
rect 12725 19873 12759 19907
rect 16037 19873 16071 19907
rect 19717 19873 19751 19907
rect 4261 19805 4295 19839
rect 7849 19805 7883 19839
rect 9919 19805 9953 19839
rect 11069 19805 11103 19839
rect 11529 19805 11563 19839
rect 18245 19805 18279 19839
rect 20913 19805 20947 19839
rect 8769 19669 8803 19703
rect 10241 19669 10275 19703
rect 20177 19669 20211 19703
rect 6193 19465 6227 19499
rect 11069 19465 11103 19499
rect 11345 19465 11379 19499
rect 17877 19465 17911 19499
rect 19349 19465 19383 19499
rect 16497 19397 16531 19431
rect 4261 19329 4295 19363
rect 5917 19329 5951 19363
rect 7573 19329 7607 19363
rect 8493 19329 8527 19363
rect 9505 19329 9539 19363
rect 13553 19329 13587 19363
rect 15393 19329 15427 19363
rect 18797 19329 18831 19363
rect 19901 19329 19935 19363
rect 20177 19329 20211 19363
rect 5089 19261 5123 19295
rect 5457 19261 5491 19295
rect 5733 19261 5767 19295
rect 10241 19261 10275 19295
rect 10425 19261 10459 19295
rect 12909 19261 12943 19295
rect 13369 19261 13403 19295
rect 3065 19193 3099 19227
rect 3617 19193 3651 19227
rect 3709 19193 3743 19227
rect 6929 19193 6963 19227
rect 7021 19193 7055 19227
rect 8585 19193 8619 19227
rect 9137 19193 9171 19227
rect 14197 19261 14231 19295
rect 14473 19261 14507 19295
rect 15577 19261 15611 19295
rect 19717 19261 19751 19295
rect 14657 19193 14691 19227
rect 15898 19193 15932 19227
rect 17417 19193 17451 19227
rect 18337 19193 18371 19227
rect 18429 19193 18463 19227
rect 19993 19193 20027 19227
rect 2513 19125 2547 19159
rect 3433 19125 3467 19159
rect 4537 19125 4571 19159
rect 6653 19125 6687 19159
rect 7849 19125 7883 19159
rect 8309 19125 8343 19159
rect 9781 19125 9815 19159
rect 10057 19125 10091 19159
rect 12817 19125 12851 19159
rect 13093 19125 13127 19159
rect 13553 19125 13587 19159
rect 13737 19125 13771 19159
rect 16773 19125 16807 19159
rect 3893 18921 3927 18955
rect 8401 18921 8435 18955
rect 8769 18921 8803 18955
rect 12725 18921 12759 18955
rect 14749 18921 14783 18955
rect 16129 18921 16163 18955
rect 16589 18921 16623 18955
rect 17141 18921 17175 18955
rect 18981 18921 19015 18955
rect 19671 18921 19705 18955
rect 20085 18921 20119 18955
rect 3249 18853 3283 18887
rect 4077 18853 4111 18887
rect 6009 18853 6043 18887
rect 6929 18853 6963 18887
rect 7573 18853 7607 18887
rect 9873 18853 9907 18887
rect 11713 18853 11747 18887
rect 14381 18853 14415 18887
rect 15577 18853 15611 18887
rect 18153 18853 18187 18887
rect 1444 18785 1478 18819
rect 2881 18785 2915 18819
rect 4721 18785 4755 18819
rect 6561 18785 6595 18819
rect 13829 18785 13863 18819
rect 14105 18785 14139 18819
rect 19568 18785 19602 18819
rect 5917 18717 5951 18751
rect 7481 18717 7515 18751
rect 7757 18717 7791 18751
rect 9413 18717 9447 18751
rect 9781 18717 9815 18751
rect 10057 18717 10091 18751
rect 11621 18717 11655 18751
rect 12265 18717 12299 18751
rect 16221 18717 16255 18751
rect 17877 18717 17911 18751
rect 18061 18717 18095 18751
rect 18429 18717 18463 18751
rect 5641 18649 5675 18683
rect 1547 18581 1581 18615
rect 3525 18581 3559 18615
rect 5273 18581 5307 18615
rect 7297 18581 7331 18615
rect 11345 18581 11379 18615
rect 4353 18377 4387 18411
rect 6653 18377 6687 18411
rect 8677 18377 8711 18411
rect 17877 18377 17911 18411
rect 2605 18309 2639 18343
rect 6285 18309 6319 18343
rect 16221 18309 16255 18343
rect 19441 18309 19475 18343
rect 2237 18241 2271 18275
rect 9321 18241 9355 18275
rect 9597 18241 9631 18275
rect 12541 18241 12575 18275
rect 12817 18241 12851 18275
rect 14749 18241 14783 18275
rect 18429 18241 18463 18275
rect 20361 18241 20395 18275
rect 1476 18173 1510 18207
rect 2421 18173 2455 18207
rect 3433 18173 3467 18207
rect 5181 18173 5215 18207
rect 5733 18173 5767 18207
rect 7481 18173 7515 18207
rect 8401 18173 8435 18207
rect 9045 18173 9079 18207
rect 10701 18173 10735 18207
rect 11437 18173 11471 18207
rect 13737 18173 13771 18207
rect 16957 18173 16991 18207
rect 9413 18105 9447 18139
rect 11529 18105 11563 18139
rect 12633 18105 12667 18139
rect 16497 18105 16531 18139
rect 18153 18105 18187 18139
rect 18245 18105 18279 18139
rect 19165 18105 19199 18139
rect 19717 18105 19751 18139
rect 19809 18105 19843 18139
rect 1547 18037 1581 18071
rect 1961 18037 1995 18071
rect 3065 18037 3099 18071
rect 3801 18037 3835 18071
rect 4721 18037 4755 18071
rect 5089 18037 5123 18071
rect 5457 18037 5491 18071
rect 7297 18037 7331 18071
rect 7849 18037 7883 18071
rect 10241 18037 10275 18071
rect 11805 18037 11839 18071
rect 12265 18037 12299 18071
rect 14105 18037 14139 18071
rect 14657 18037 14691 18071
rect 15117 18037 15151 18071
rect 15669 18037 15703 18071
rect 17509 18037 17543 18071
rect 1685 17833 1719 17867
rect 5273 17833 5307 17867
rect 6469 17833 6503 17867
rect 6929 17833 6963 17867
rect 7757 17833 7791 17867
rect 8309 17833 8343 17867
rect 15853 17833 15887 17867
rect 17693 17833 17727 17867
rect 19303 17833 19337 17867
rect 19625 17833 19659 17867
rect 5911 17765 5945 17799
rect 9321 17765 9355 17799
rect 11621 17765 11655 17799
rect 13093 17765 13127 17799
rect 13185 17765 13219 17799
rect 13737 17765 13771 17799
rect 14565 17765 14599 17799
rect 16129 17765 16163 17799
rect 16221 17765 16255 17799
rect 16773 17765 16807 17799
rect 1961 17697 1995 17731
rect 2973 17697 3007 17731
rect 4604 17697 4638 17731
rect 9965 17697 9999 17731
rect 10149 17697 10183 17731
rect 17601 17697 17635 17731
rect 18061 17697 18095 17731
rect 19165 17697 19199 17731
rect 5549 17629 5583 17663
rect 7389 17629 7423 17663
rect 10241 17629 10275 17663
rect 11529 17629 11563 17663
rect 11897 17629 11931 17663
rect 2513 17561 2547 17595
rect 4675 17561 4709 17595
rect 12541 17561 12575 17595
rect 2145 17493 2179 17527
rect 3157 17493 3191 17527
rect 3433 17493 3467 17527
rect 4261 17493 4295 17527
rect 7205 17493 7239 17527
rect 8585 17493 8619 17527
rect 10701 17493 10735 17527
rect 12909 17493 12943 17527
rect 17417 17493 17451 17527
rect 18613 17493 18647 17527
rect 18981 17493 19015 17527
rect 2053 17289 2087 17323
rect 3341 17289 3375 17323
rect 4813 17289 4847 17323
rect 6193 17289 6227 17323
rect 6653 17289 6687 17323
rect 7113 17289 7147 17323
rect 9873 17289 9907 17323
rect 11529 17289 11563 17323
rect 13829 17289 13863 17323
rect 15669 17289 15703 17323
rect 20085 17289 20119 17323
rect 4905 17221 4939 17255
rect 5641 17221 5675 17255
rect 11253 17221 11287 17255
rect 13461 17221 13495 17255
rect 24777 17221 24811 17255
rect 1409 17085 1443 17119
rect 2789 17085 2823 17119
rect 2881 17085 2915 17119
rect 3893 17085 3927 17119
rect 5733 17153 5767 17187
rect 9505 17153 9539 17187
rect 10333 17153 10367 17187
rect 12541 17153 12575 17187
rect 12817 17153 12851 17187
rect 15301 17153 15335 17187
rect 18245 17153 18279 17187
rect 6745 17085 6779 17119
rect 7297 17085 7331 17119
rect 8033 17085 8067 17119
rect 8493 17085 8527 17119
rect 8953 17085 8987 17119
rect 9229 17085 9263 17119
rect 14565 17085 14599 17119
rect 15025 17085 15059 17119
rect 16129 17085 16163 17119
rect 18889 17085 18923 17119
rect 19876 17085 19910 17119
rect 20269 17085 20303 17119
rect 24593 17085 24627 17119
rect 25145 17085 25179 17119
rect 3709 17017 3743 17051
rect 4255 17017 4289 17051
rect 4905 17017 4939 17051
rect 5181 17017 5215 17051
rect 10695 17017 10729 17051
rect 12265 17017 12299 17051
rect 12633 17017 12667 17051
rect 16450 17017 16484 17051
rect 18337 17017 18371 17051
rect 1593 16949 1627 16983
rect 2421 16949 2455 16983
rect 3065 16949 3099 16983
rect 7757 16949 7791 16983
rect 10149 16949 10183 16983
rect 14473 16949 14507 16983
rect 15945 16949 15979 16983
rect 17049 16949 17083 16983
rect 17601 16949 17635 16983
rect 19165 16949 19199 16983
rect 3801 16745 3835 16779
rect 4169 16745 4203 16779
rect 8493 16745 8527 16779
rect 9505 16745 9539 16779
rect 10149 16745 10183 16779
rect 10701 16745 10735 16779
rect 11345 16745 11379 16779
rect 16773 16745 16807 16779
rect 17325 16745 17359 16779
rect 19717 16745 19751 16779
rect 9045 16677 9079 16711
rect 11713 16677 11747 16711
rect 12265 16677 12299 16711
rect 13093 16677 13127 16711
rect 18337 16677 18371 16711
rect 18889 16677 18923 16711
rect 1961 16609 1995 16643
rect 3008 16609 3042 16643
rect 4077 16609 4111 16643
rect 4721 16609 4755 16643
rect 4905 16609 4939 16643
rect 5457 16609 5491 16643
rect 7205 16609 7239 16643
rect 7389 16609 7423 16643
rect 8585 16609 8619 16643
rect 13461 16609 13495 16643
rect 15209 16609 15243 16643
rect 16405 16609 16439 16643
rect 24501 16609 24535 16643
rect 2145 16541 2179 16575
rect 7481 16541 7515 16575
rect 9781 16541 9815 16575
rect 10977 16541 11011 16575
rect 11621 16541 11655 16575
rect 18245 16541 18279 16575
rect 2789 16473 2823 16507
rect 3111 16473 3145 16507
rect 8769 16473 8803 16507
rect 15439 16473 15473 16507
rect 2421 16405 2455 16439
rect 3433 16405 3467 16439
rect 8033 16405 8067 16439
rect 14381 16405 14415 16439
rect 15853 16405 15887 16439
rect 16129 16405 16163 16439
rect 17693 16405 17727 16439
rect 18061 16405 18095 16439
rect 21373 16405 21407 16439
rect 24731 16405 24765 16439
rect 2973 16201 3007 16235
rect 7159 16201 7193 16235
rect 11805 16201 11839 16235
rect 13461 16201 13495 16235
rect 15301 16201 15335 16235
rect 16773 16201 16807 16235
rect 17785 16201 17819 16235
rect 19165 16201 19199 16235
rect 24685 16201 24719 16235
rect 5733 16133 5767 16167
rect 6653 16133 6687 16167
rect 9873 16133 9907 16167
rect 11345 16133 11379 16167
rect 17509 16133 17543 16167
rect 1685 16065 1719 16099
rect 2697 16065 2731 16099
rect 6929 16065 6963 16099
rect 9505 16065 9539 16099
rect 11069 16065 11103 16099
rect 18245 16065 18279 16099
rect 18889 16065 18923 16099
rect 20085 16065 20119 16099
rect 21373 16065 21407 16099
rect 21649 16065 21683 16099
rect 4077 15997 4111 16031
rect 4721 15997 4755 16031
rect 4905 15997 4939 16031
rect 5365 15997 5399 16031
rect 7481 15997 7515 16031
rect 8033 15997 8067 16031
rect 8493 15997 8527 16031
rect 8953 15997 8987 16031
rect 9229 15997 9263 16031
rect 10333 15997 10367 16031
rect 10425 15997 10459 16031
rect 10609 15997 10643 16031
rect 12541 15997 12575 16031
rect 14197 15997 14231 16031
rect 14565 15997 14599 16031
rect 14841 15997 14875 16031
rect 15853 15997 15887 16031
rect 1777 15929 1811 15963
rect 2329 15929 2363 15963
rect 3525 15929 3559 15963
rect 3801 15929 3835 15963
rect 6285 15929 6319 15963
rect 12449 15929 12483 15963
rect 15025 15929 15059 15963
rect 16174 15929 16208 15963
rect 17049 15929 17083 15963
rect 18337 15929 18371 15963
rect 19809 15929 19843 15963
rect 19901 15929 19935 15963
rect 21189 15929 21223 15963
rect 21465 15929 21499 15963
rect 4077 15861 4111 15895
rect 7849 15861 7883 15895
rect 10149 15861 10183 15895
rect 12265 15861 12299 15895
rect 15669 15861 15703 15895
rect 19533 15861 19567 15895
rect 3433 15657 3467 15691
rect 6469 15657 6503 15691
rect 8677 15657 8711 15691
rect 10149 15657 10183 15691
rect 11621 15657 11655 15691
rect 15669 15657 15703 15691
rect 16221 15657 16255 15691
rect 1777 15589 1811 15623
rect 1869 15589 1903 15623
rect 3893 15589 3927 15623
rect 4261 15589 4295 15623
rect 5825 15589 5859 15623
rect 12081 15589 12115 15623
rect 18061 15589 18095 15623
rect 5549 15521 5583 15555
rect 6009 15521 6043 15555
rect 6285 15521 6319 15555
rect 7389 15521 7423 15555
rect 7665 15521 7699 15555
rect 9689 15521 9723 15555
rect 9965 15521 9999 15555
rect 13553 15521 13587 15555
rect 15853 15521 15887 15555
rect 19441 15521 19475 15555
rect 4169 15453 4203 15487
rect 4445 15453 4479 15487
rect 5089 15453 5123 15487
rect 7573 15453 7607 15487
rect 11989 15453 12023 15487
rect 12357 15453 12391 15487
rect 13461 15453 13495 15487
rect 17969 15453 18003 15487
rect 20913 15453 20947 15487
rect 2329 15385 2363 15419
rect 3157 15385 3191 15419
rect 6101 15385 6135 15419
rect 9321 15385 9355 15419
rect 9781 15385 9815 15419
rect 18521 15385 18555 15419
rect 2697 15317 2731 15351
rect 7021 15317 7055 15351
rect 9045 15317 9079 15351
rect 10793 15317 10827 15351
rect 11069 15317 11103 15351
rect 12909 15317 12943 15351
rect 13277 15317 13311 15351
rect 16773 15317 16807 15351
rect 17785 15317 17819 15351
rect 18981 15317 19015 15351
rect 19579 15317 19613 15351
rect 6561 15113 6595 15147
rect 10241 15113 10275 15147
rect 10333 15113 10367 15147
rect 11989 15113 12023 15147
rect 17417 15113 17451 15147
rect 17877 15113 17911 15147
rect 2697 14977 2731 15011
rect 4537 14909 4571 14943
rect 4905 14909 4939 14943
rect 5457 14909 5491 14943
rect 5825 14909 5859 14943
rect 6837 14909 6871 14943
rect 7573 14909 7607 14943
rect 7941 14909 7975 14943
rect 8401 14909 8435 14943
rect 8769 14909 8803 14943
rect 9137 14909 9171 14943
rect 3018 14841 3052 14875
rect 9413 14841 9447 14875
rect 13093 15045 13127 15079
rect 21373 15045 21407 15079
rect 10517 14977 10551 15011
rect 12541 14977 12575 15011
rect 18153 14977 18187 15011
rect 18429 14977 18463 15011
rect 19165 14977 19199 15011
rect 19993 14977 20027 15011
rect 14473 14909 14507 14943
rect 14933 14909 14967 14943
rect 15209 14909 15243 14943
rect 16037 14909 16071 14943
rect 16957 14909 16991 14943
rect 21189 14909 21223 14943
rect 21649 14909 21683 14943
rect 1409 14773 1443 14807
rect 1961 14773 1995 14807
rect 2605 14773 2639 14807
rect 3617 14773 3651 14807
rect 4077 14773 4111 14807
rect 4537 14773 4571 14807
rect 6285 14773 6319 14807
rect 7021 14773 7055 14807
rect 9689 14773 9723 14807
rect 10241 14773 10275 14807
rect 12633 14841 12667 14875
rect 16358 14841 16392 14875
rect 18245 14841 18279 14875
rect 19717 14841 19751 14875
rect 19809 14841 19843 14875
rect 10885 14773 10919 14807
rect 11437 14773 11471 14807
rect 13553 14773 13587 14807
rect 14289 14773 14323 14807
rect 15485 14773 15519 14807
rect 15853 14773 15887 14807
rect 19441 14773 19475 14807
rect 2421 14569 2455 14603
rect 3249 14569 3283 14603
rect 4721 14569 4755 14603
rect 6193 14569 6227 14603
rect 10149 14569 10183 14603
rect 11897 14569 11931 14603
rect 14565 14569 14599 14603
rect 16497 14569 16531 14603
rect 18245 14569 18279 14603
rect 1863 14501 1897 14535
rect 2789 14501 2823 14535
rect 8585 14501 8619 14535
rect 11022 14501 11056 14535
rect 12633 14501 12667 14535
rect 13185 14501 13219 14535
rect 15622 14501 15656 14535
rect 17233 14501 17267 14535
rect 17325 14501 17359 14535
rect 17877 14501 17911 14535
rect 18797 14501 18831 14535
rect 18889 14501 18923 14535
rect 1501 14433 1535 14467
rect 4445 14433 4479 14467
rect 4905 14433 4939 14467
rect 5457 14433 5491 14467
rect 5825 14433 5859 14467
rect 6837 14433 6871 14467
rect 9137 14433 9171 14467
rect 9724 14433 9758 14467
rect 9827 14433 9861 14467
rect 14064 14433 14098 14467
rect 20821 14433 20855 14467
rect 24593 14433 24627 14467
rect 4353 14365 4387 14399
rect 6745 14365 6779 14399
rect 8309 14365 8343 14399
rect 10701 14365 10735 14399
rect 12541 14365 12575 14399
rect 13461 14365 13495 14399
rect 14151 14365 14185 14399
rect 15301 14365 15335 14399
rect 18521 14365 18555 14399
rect 19073 14365 19107 14399
rect 11621 14297 11655 14331
rect 24777 14297 24811 14331
rect 3893 14229 3927 14263
rect 6653 14229 6687 14263
rect 7941 14229 7975 14263
rect 9413 14229 9447 14263
rect 10517 14229 10551 14263
rect 12357 14229 12391 14263
rect 16221 14229 16255 14263
rect 19809 14229 19843 14263
rect 21051 14229 21085 14263
rect 2973 14025 3007 14059
rect 4537 14025 4571 14059
rect 4905 14025 4939 14059
rect 6285 14025 6319 14059
rect 9689 14025 9723 14059
rect 11621 14025 11655 14059
rect 12265 14025 12299 14059
rect 13737 14025 13771 14059
rect 17233 14025 17267 14059
rect 17877 14025 17911 14059
rect 19073 14025 19107 14059
rect 24731 14025 24765 14059
rect 25053 14025 25087 14059
rect 6653 13957 6687 13991
rect 9965 13957 9999 13991
rect 10333 13957 10367 13991
rect 11253 13957 11287 13991
rect 14013 13957 14047 13991
rect 21465 13957 21499 13991
rect 1685 13889 1719 13923
rect 9413 13889 9447 13923
rect 13185 13889 13219 13923
rect 15117 13889 15151 13923
rect 15853 13889 15887 13923
rect 18429 13889 18463 13923
rect 4721 13821 4755 13855
rect 5549 13821 5583 13855
rect 5733 13821 5767 13855
rect 7757 13821 7791 13855
rect 7941 13821 7975 13855
rect 8401 13821 8435 13855
rect 8769 13821 8803 13855
rect 9137 13821 9171 13855
rect 9965 13821 9999 13855
rect 10057 13821 10091 13855
rect 10241 13821 10275 13855
rect 10517 13821 10551 13855
rect 14473 13821 14507 13855
rect 14933 13821 14967 13855
rect 15945 13821 15979 13855
rect 16497 13821 16531 13855
rect 19692 13821 19726 13855
rect 20085 13821 20119 13855
rect 20672 13821 20706 13855
rect 21097 13821 21131 13855
rect 24660 13821 24694 13855
rect 1777 13753 1811 13787
rect 2329 13753 2363 13787
rect 3249 13753 3283 13787
rect 3341 13753 3375 13787
rect 3893 13753 3927 13787
rect 7389 13753 7423 13787
rect 10977 13753 11011 13787
rect 12541 13753 12575 13787
rect 12633 13753 12667 13787
rect 18153 13753 18187 13787
rect 18245 13753 18279 13787
rect 25513 13753 25547 13787
rect 2605 13685 2639 13719
rect 5181 13685 5215 13719
rect 5917 13685 5951 13719
rect 6929 13685 6963 13719
rect 15393 13685 15427 13719
rect 16037 13685 16071 13719
rect 19441 13685 19475 13719
rect 19763 13685 19797 13719
rect 20775 13685 20809 13719
rect 3249 13481 3283 13515
rect 5825 13481 5859 13515
rect 7573 13481 7607 13515
rect 10241 13481 10275 13515
rect 10563 13481 10597 13515
rect 12541 13481 12575 13515
rect 14381 13481 14415 13515
rect 15117 13481 15151 13515
rect 16313 13481 16347 13515
rect 17233 13481 17267 13515
rect 17463 13481 17497 13515
rect 1685 13413 1719 13447
rect 2237 13413 2271 13447
rect 4077 13413 4111 13447
rect 5089 13413 5123 13447
rect 9413 13413 9447 13447
rect 11621 13413 11655 13447
rect 13093 13413 13127 13447
rect 13185 13413 13219 13447
rect 16037 13413 16071 13447
rect 18521 13413 18555 13447
rect 19073 13413 19107 13447
rect 4169 13345 4203 13379
rect 6193 13345 6227 13379
rect 6469 13345 6503 13379
rect 8033 13345 8067 13379
rect 8309 13345 8343 13379
rect 10460 13345 10494 13379
rect 15301 13345 15335 13379
rect 15853 13345 15887 13379
rect 17325 13345 17359 13379
rect 20948 13345 20982 13379
rect 23648 13345 23682 13379
rect 1593 13277 1627 13311
rect 2881 13277 2915 13311
rect 3893 13277 3927 13311
rect 6929 13277 6963 13311
rect 8493 13277 8527 13311
rect 9873 13277 9907 13311
rect 11529 13277 11563 13311
rect 13369 13277 13403 13311
rect 18245 13277 18279 13311
rect 18429 13277 18463 13311
rect 2605 13209 2639 13243
rect 5457 13209 5491 13243
rect 6285 13209 6319 13243
rect 8125 13209 8159 13243
rect 12081 13209 12115 13243
rect 16773 13209 16807 13243
rect 21051 13209 21085 13243
rect 7849 13141 7883 13175
rect 9137 13141 9171 13175
rect 10885 13141 10919 13175
rect 12817 13141 12851 13175
rect 18153 13141 18187 13175
rect 18245 13141 18279 13175
rect 23719 13141 23753 13175
rect 2421 12937 2455 12971
rect 6561 12937 6595 12971
rect 10333 12937 10367 12971
rect 13829 12937 13863 12971
rect 14289 12937 14323 12971
rect 15945 12937 15979 12971
rect 19073 12937 19107 12971
rect 19441 12937 19475 12971
rect 19763 12937 19797 12971
rect 21097 12937 21131 12971
rect 23857 12937 23891 12971
rect 1501 12869 1535 12903
rect 3985 12869 4019 12903
rect 4629 12869 4663 12903
rect 5917 12869 5951 12903
rect 9965 12869 9999 12903
rect 11345 12869 11379 12903
rect 13093 12869 13127 12903
rect 14657 12869 14691 12903
rect 9597 12801 9631 12835
rect 10425 12801 10459 12835
rect 11713 12801 11747 12835
rect 14933 12801 14967 12835
rect 16497 12801 16531 12835
rect 18153 12801 18187 12835
rect 20775 12801 20809 12835
rect 1409 12733 1443 12767
rect 1685 12733 1719 12767
rect 4537 12733 4571 12767
rect 4813 12733 4847 12767
rect 8217 12733 8251 12767
rect 8585 12733 8619 12767
rect 9045 12733 9079 12767
rect 9321 12733 9355 12767
rect 17141 12733 17175 12767
rect 19692 12733 19726 12767
rect 20688 12733 20722 12767
rect 21465 12733 21499 12767
rect 2145 12665 2179 12699
rect 3065 12665 3099 12699
rect 3157 12665 3191 12699
rect 3709 12665 3743 12699
rect 7573 12665 7607 12699
rect 12541 12665 12575 12699
rect 12633 12665 12667 12699
rect 15025 12665 15059 12699
rect 15577 12665 15611 12699
rect 16589 12665 16623 12699
rect 18245 12665 18279 12699
rect 18797 12665 18831 12699
rect 2881 12597 2915 12631
rect 4353 12597 4387 12631
rect 4997 12597 5031 12631
rect 6193 12597 6227 12631
rect 6837 12597 6871 12631
rect 7941 12597 7975 12631
rect 10793 12597 10827 12631
rect 12265 12597 12299 12631
rect 13553 12597 13587 12631
rect 16221 12597 16255 12631
rect 17417 12597 17451 12631
rect 17785 12597 17819 12631
rect 20177 12597 20211 12631
rect 1869 12393 1903 12427
rect 2881 12393 2915 12427
rect 3525 12393 3559 12427
rect 3801 12393 3835 12427
rect 4169 12393 4203 12427
rect 7021 12393 7055 12427
rect 9413 12393 9447 12427
rect 9781 12393 9815 12427
rect 11897 12393 11931 12427
rect 13093 12393 13127 12427
rect 14933 12393 14967 12427
rect 1409 12257 1443 12291
rect 2881 12257 2915 12291
rect 4353 12257 4387 12291
rect 4813 12257 4847 12291
rect 4997 12257 5031 12291
rect 5273 12257 5307 12291
rect 6837 12257 6871 12291
rect 1593 12121 1627 12155
rect 5917 12121 5951 12155
rect 12173 12325 12207 12359
rect 16266 12325 16300 12359
rect 17785 12325 17819 12359
rect 17877 12325 17911 12359
rect 7573 12257 7607 12291
rect 7757 12257 7791 12291
rect 8309 12257 8343 12291
rect 8585 12257 8619 12291
rect 9965 12257 9999 12291
rect 10149 12257 10183 12291
rect 10517 12257 10551 12291
rect 10885 12257 10919 12291
rect 13645 12257 13679 12291
rect 19257 12257 19291 12291
rect 19717 12257 19751 12291
rect 20980 12257 21014 12291
rect 23648 12257 23682 12291
rect 12081 12189 12115 12223
rect 13553 12189 13587 12223
rect 15945 12189 15979 12223
rect 19809 12189 19843 12223
rect 8677 12121 8711 12155
rect 12633 12121 12667 12155
rect 18337 12121 18371 12155
rect 2237 12053 2271 12087
rect 6193 12053 6227 12087
rect 7021 12053 7055 12087
rect 7113 12053 7147 12087
rect 9045 12053 9079 12087
rect 11437 12053 11471 12087
rect 16865 12053 16899 12087
rect 17233 12053 17267 12087
rect 18797 12053 18831 12087
rect 21051 12053 21085 12087
rect 23719 12053 23753 12087
rect 6193 11849 6227 11883
rect 7021 11849 7055 11883
rect 9873 11849 9907 11883
rect 10333 11849 10367 11883
rect 13645 11849 13679 11883
rect 15393 11849 15427 11883
rect 20775 11849 20809 11883
rect 23857 11849 23891 11883
rect 24777 11849 24811 11883
rect 6653 11781 6687 11815
rect 14289 11781 14323 11815
rect 19763 11781 19797 11815
rect 1547 11713 1581 11747
rect 7389 11713 7423 11747
rect 9597 11713 9631 11747
rect 10425 11713 10459 11747
rect 12265 11713 12299 11747
rect 12541 11713 12575 11747
rect 13185 11713 13219 11747
rect 16497 11713 16531 11747
rect 18153 11713 18187 11747
rect 19257 11713 19291 11747
rect 1444 11645 1478 11679
rect 1869 11645 1903 11679
rect 2697 11645 2731 11679
rect 4721 11645 4755 11679
rect 4905 11645 4939 11679
rect 5457 11645 5491 11679
rect 5825 11645 5859 11679
rect 6837 11645 6871 11679
rect 7665 11645 7699 11679
rect 8217 11645 8251 11679
rect 8585 11645 8619 11679
rect 8953 11645 8987 11679
rect 9413 11645 9447 11679
rect 14473 11645 14507 11679
rect 15945 11645 15979 11679
rect 19660 11645 19694 11679
rect 20085 11645 20119 11679
rect 20704 11645 20738 11679
rect 24593 11645 24627 11679
rect 25145 11645 25179 11679
rect 2605 11577 2639 11611
rect 3018 11577 3052 11611
rect 5917 11577 5951 11611
rect 12633 11577 12667 11611
rect 14835 11577 14869 11611
rect 16589 11577 16623 11611
rect 17141 11577 17175 11611
rect 18245 11577 18279 11611
rect 18797 11577 18831 11611
rect 21189 11577 21223 11611
rect 3617 11509 3651 11543
rect 4169 11509 4203 11543
rect 10793 11509 10827 11543
rect 11345 11509 11379 11543
rect 11805 11509 11839 11543
rect 13921 11509 13955 11543
rect 17693 11509 17727 11543
rect 21465 11509 21499 11543
rect 2421 11305 2455 11339
rect 2881 11305 2915 11339
rect 3157 11305 3191 11339
rect 3893 11305 3927 11339
rect 4997 11305 5031 11339
rect 5457 11305 5491 11339
rect 9413 11305 9447 11339
rect 10977 11305 11011 11339
rect 11437 11305 11471 11339
rect 12541 11305 12575 11339
rect 16589 11305 16623 11339
rect 18153 11305 18187 11339
rect 19625 11305 19659 11339
rect 24777 11305 24811 11339
rect 3525 11237 3559 11271
rect 6653 11237 6687 11271
rect 7021 11237 7055 11271
rect 7573 11237 7607 11271
rect 8217 11237 8251 11271
rect 11713 11237 11747 11271
rect 15663 11237 15697 11271
rect 17233 11237 17267 11271
rect 18429 11237 18463 11271
rect 18797 11237 18831 11271
rect 1777 11169 1811 11203
rect 2973 11169 3007 11203
rect 4123 11169 4157 11203
rect 4537 11169 4571 11203
rect 8620 11169 8654 11203
rect 9965 11169 9999 11203
rect 10425 11169 10459 11203
rect 13921 11169 13955 11203
rect 14105 11169 14139 11203
rect 21373 11169 21407 11203
rect 24593 11169 24627 11203
rect 5089 11101 5123 11135
rect 6929 11101 6963 11135
rect 10701 11101 10735 11135
rect 11621 11101 11655 11135
rect 11897 11101 11931 11135
rect 14381 11101 14415 11135
rect 15301 11101 15335 11135
rect 17141 11101 17175 11135
rect 18705 11101 18739 11135
rect 18981 11101 19015 11135
rect 4215 11033 4249 11067
rect 6285 11033 6319 11067
rect 17693 11033 17727 11067
rect 1685 10965 1719 10999
rect 6009 10965 6043 10999
rect 8723 10965 8757 10999
rect 9137 10965 9171 10999
rect 12909 10965 12943 10999
rect 14933 10965 14967 10999
rect 16221 10965 16255 10999
rect 16865 10965 16899 10999
rect 21557 10965 21591 10999
rect 2513 10761 2547 10795
rect 4537 10761 4571 10795
rect 5089 10761 5123 10795
rect 6285 10761 6319 10795
rect 8217 10761 8251 10795
rect 8585 10761 8619 10795
rect 11805 10761 11839 10795
rect 14381 10761 14415 10795
rect 15945 10761 15979 10795
rect 16865 10761 16899 10795
rect 19441 10761 19475 10795
rect 19809 10761 19843 10795
rect 21373 10761 21407 10795
rect 24685 10761 24719 10795
rect 1593 10625 1627 10659
rect 2881 10625 2915 10659
rect 3709 10625 3743 10659
rect 3985 10625 4019 10659
rect 1501 10557 1535 10591
rect 1777 10557 1811 10591
rect 3249 10557 3283 10591
rect 2237 10489 2271 10523
rect 3801 10489 3835 10523
rect 4721 10693 4755 10727
rect 5825 10693 5859 10727
rect 13645 10693 13679 10727
rect 19073 10693 19107 10727
rect 6653 10625 6687 10659
rect 6837 10625 6871 10659
rect 11529 10625 11563 10659
rect 12541 10625 12575 10659
rect 15025 10625 15059 10659
rect 15669 10625 15703 10659
rect 18153 10625 18187 10659
rect 18429 10625 18463 10659
rect 6929 10557 6963 10591
rect 8953 10557 8987 10591
rect 9413 10557 9447 10591
rect 10333 10557 10367 10591
rect 11345 10557 11379 10591
rect 13185 10557 13219 10591
rect 19625 10557 19659 10591
rect 20085 10557 20119 10591
rect 5273 10489 5307 10523
rect 5365 10489 5399 10523
rect 9689 10489 9723 10523
rect 12633 10489 12667 10523
rect 14841 10489 14875 10523
rect 15117 10489 15151 10523
rect 16957 10489 16991 10523
rect 17785 10489 17819 10523
rect 18245 10489 18279 10523
rect 4537 10421 4571 10455
rect 9965 10421 9999 10455
rect 12173 10421 12207 10455
rect 14013 10421 14047 10455
rect 17509 10421 17543 10455
rect 2421 10217 2455 10251
rect 2789 10217 2823 10251
rect 3157 10217 3191 10251
rect 3433 10217 3467 10251
rect 4261 10217 4295 10251
rect 4629 10217 4663 10251
rect 6101 10217 6135 10251
rect 7113 10217 7147 10251
rect 9045 10217 9079 10251
rect 9873 10217 9907 10251
rect 11437 10217 11471 10251
rect 11805 10217 11839 10251
rect 13921 10217 13955 10251
rect 15945 10217 15979 10251
rect 16497 10217 16531 10251
rect 17141 10217 17175 10251
rect 17693 10217 17727 10251
rect 18245 10217 18279 10251
rect 2145 10149 2179 10183
rect 6469 10149 6503 10183
rect 10241 10149 10275 10183
rect 10517 10149 10551 10183
rect 10609 10149 10643 10183
rect 12173 10149 12207 10183
rect 19211 10149 19245 10183
rect 1501 10081 1535 10115
rect 2973 10081 3007 10115
rect 4077 10081 4111 10115
rect 5089 10081 5123 10115
rect 5365 10081 5399 10115
rect 5825 10081 5859 10115
rect 6653 10081 6687 10115
rect 8125 10081 8159 10115
rect 8493 10081 8527 10115
rect 13921 10081 13955 10115
rect 14105 10081 14139 10115
rect 19124 10081 19158 10115
rect 8769 10013 8803 10047
rect 12081 10013 12115 10047
rect 12725 10013 12759 10047
rect 15577 10013 15611 10047
rect 17325 10013 17359 10047
rect 3893 9945 3927 9979
rect 5181 9945 5215 9979
rect 11069 9945 11103 9979
rect 4997 9877 5031 9911
rect 6837 9877 6871 9911
rect 7849 9877 7883 9911
rect 14657 9877 14691 9911
rect 2421 9673 2455 9707
rect 11253 9673 11287 9707
rect 13737 9673 13771 9707
rect 15301 9673 15335 9707
rect 15577 9673 15611 9707
rect 17877 9673 17911 9707
rect 19257 9673 19291 9707
rect 2789 9605 2823 9639
rect 3157 9605 3191 9639
rect 7021 9605 7055 9639
rect 9137 9605 9171 9639
rect 1501 9537 1535 9571
rect 1869 9537 1903 9571
rect 4353 9537 4387 9571
rect 7941 9537 7975 9571
rect 9413 9537 9447 9571
rect 9505 9537 9539 9571
rect 9689 9537 9723 9571
rect 14381 9537 14415 9571
rect 18521 9537 18555 9571
rect 1409 9469 1443 9503
rect 1685 9469 1719 9503
rect 3893 9469 3927 9503
rect 4077 9469 4111 9503
rect 4721 9469 4755 9503
rect 5181 9469 5215 9503
rect 5273 9469 5307 9503
rect 5457 9469 5491 9503
rect 6561 9469 6595 9503
rect 6837 9469 6871 9503
rect 11989 9469 12023 9503
rect 15945 9469 15979 9503
rect 17325 9469 17359 9503
rect 5917 9401 5951 9435
rect 7757 9401 7791 9435
rect 8262 9401 8296 9435
rect 9413 9401 9447 9435
rect 10010 9401 10044 9435
rect 11713 9401 11747 9435
rect 12541 9401 12575 9435
rect 12633 9401 12667 9435
rect 13185 9401 13219 9435
rect 14105 9401 14139 9435
rect 14197 9401 14231 9435
rect 16266 9401 16300 9435
rect 18245 9401 18279 9435
rect 18337 9401 18371 9435
rect 4997 9333 5031 9367
rect 6193 9333 6227 9367
rect 7297 9333 7331 9367
rect 8861 9333 8895 9367
rect 10609 9333 10643 9367
rect 10977 9333 11011 9367
rect 16865 9333 16899 9367
rect 2881 9129 2915 9163
rect 3157 9129 3191 9163
rect 3709 9129 3743 9163
rect 7113 9129 7147 9163
rect 7849 9129 7883 9163
rect 9873 9129 9907 9163
rect 11989 9129 12023 9163
rect 12449 9129 12483 9163
rect 13737 9129 13771 9163
rect 14381 9129 14415 9163
rect 16681 9129 16715 9163
rect 18521 9129 18555 9163
rect 18843 9129 18877 9163
rect 1409 9061 1443 9095
rect 2421 9061 2455 9095
rect 5273 9061 5307 9095
rect 11390 9061 11424 9095
rect 13138 9061 13172 9095
rect 14105 9061 14139 9095
rect 17325 9061 17359 9095
rect 17877 9061 17911 9095
rect 1501 8993 1535 9027
rect 2973 8993 3007 9027
rect 4629 8993 4663 9027
rect 6101 8993 6135 9027
rect 6377 8993 6411 9027
rect 8309 8993 8343 9027
rect 8493 8993 8527 9027
rect 9689 8993 9723 9027
rect 11069 8993 11103 9027
rect 15301 8993 15335 9027
rect 15853 8993 15887 9027
rect 18705 8993 18739 9027
rect 4353 8925 4387 8959
rect 6561 8925 6595 8959
rect 8585 8925 8619 8959
rect 12817 8925 12851 8959
rect 16037 8925 16071 8959
rect 17233 8925 17267 8959
rect 18153 8925 18187 8959
rect 6193 8857 6227 8891
rect 5549 8789 5583 8823
rect 6009 8789 6043 8823
rect 10609 8789 10643 8823
rect 10977 8789 11011 8823
rect 15117 8789 15151 8823
rect 16313 8789 16347 8823
rect 3341 8585 3375 8619
rect 6101 8585 6135 8619
rect 9781 8585 9815 8619
rect 13737 8585 13771 8619
rect 15301 8585 15335 8619
rect 17141 8585 17175 8619
rect 4261 8517 4295 8551
rect 7849 8517 7883 8551
rect 9413 8517 9447 8551
rect 12173 8517 12207 8551
rect 18199 8517 18233 8551
rect 3065 8449 3099 8483
rect 5825 8449 5859 8483
rect 6929 8449 6963 8483
rect 7297 8449 7331 8483
rect 8401 8449 8435 8483
rect 8493 8449 8527 8483
rect 10885 8449 10919 8483
rect 11529 8449 11563 8483
rect 14565 8449 14599 8483
rect 16865 8449 16899 8483
rect 4077 8381 4111 8415
rect 5181 8381 5215 8415
rect 6561 8381 6595 8415
rect 6837 8381 6871 8415
rect 7113 8381 7147 8415
rect 10057 8381 10091 8415
rect 15761 8381 15795 8415
rect 16313 8381 16347 8415
rect 17877 8381 17911 8415
rect 18096 8381 18130 8415
rect 8814 8313 8848 8347
rect 10609 8313 10643 8347
rect 10701 8313 10735 8347
rect 12725 8313 12759 8347
rect 12817 8313 12851 8347
rect 13369 8313 13403 8347
rect 14289 8313 14323 8347
rect 14381 8313 14415 8347
rect 1593 8245 1627 8279
rect 3985 8245 4019 8279
rect 4537 8245 4571 8279
rect 4997 8245 5031 8279
rect 14013 8245 14047 8279
rect 16037 8245 16071 8279
rect 18797 8245 18831 8279
rect 6837 8041 6871 8075
rect 7941 8041 7975 8075
rect 9045 8041 9079 8075
rect 11253 8041 11287 8075
rect 13645 8041 13679 8075
rect 15393 8041 15427 8075
rect 16313 8041 16347 8075
rect 17233 8041 17267 8075
rect 6285 7973 6319 8007
rect 8217 7973 8251 8007
rect 10378 7973 10412 8007
rect 12817 7973 12851 8007
rect 13369 7973 13403 8007
rect 4537 7905 4571 7939
rect 5549 7905 5583 7939
rect 5825 7905 5859 7939
rect 7205 7905 7239 7939
rect 14197 7905 14231 7939
rect 15577 7905 15611 7939
rect 15853 7905 15887 7939
rect 8125 7837 8159 7871
rect 8769 7837 8803 7871
rect 10057 7837 10091 7871
rect 12725 7837 12759 7871
rect 14335 7837 14369 7871
rect 5641 7769 5675 7803
rect 4721 7701 4755 7735
rect 10977 7701 11011 7735
rect 12541 7701 12575 7735
rect 14657 7701 14691 7735
rect 6101 7497 6135 7531
rect 7021 7497 7055 7531
rect 7941 7497 7975 7531
rect 8309 7497 8343 7531
rect 9597 7497 9631 7531
rect 11897 7497 11931 7531
rect 12265 7497 12299 7531
rect 12587 7497 12621 7531
rect 13599 7497 13633 7531
rect 15393 7497 15427 7531
rect 9965 7429 9999 7463
rect 13001 7429 13035 7463
rect 10517 7361 10551 7395
rect 14289 7361 14323 7395
rect 1460 7293 1494 7327
rect 1869 7293 1903 7327
rect 5181 7293 5215 7327
rect 6837 7293 6871 7327
rect 7297 7293 7331 7327
rect 8401 7293 8435 7327
rect 12516 7293 12550 7327
rect 13496 7293 13530 7327
rect 1547 7225 1581 7259
rect 5825 7225 5859 7259
rect 6469 7225 6503 7259
rect 8722 7225 8756 7259
rect 10241 7225 10275 7259
rect 10333 7225 10367 7259
rect 13277 7225 13311 7259
rect 4537 7157 4571 7191
rect 4997 7157 5031 7191
rect 9321 7157 9355 7191
rect 11161 7157 11195 7191
rect 15669 7157 15703 7191
rect 6101 6953 6135 6987
rect 9137 6953 9171 6987
rect 10149 6953 10183 6987
rect 13875 6953 13909 6987
rect 7849 6885 7883 6919
rect 8769 6885 8803 6919
rect 10609 6885 10643 6919
rect 11345 6885 11379 6919
rect 11897 6885 11931 6919
rect 1409 6817 1443 6851
rect 5641 6817 5675 6851
rect 5733 6817 5767 6851
rect 5917 6817 5951 6851
rect 8033 6817 8067 6851
rect 8493 6817 8527 6851
rect 12792 6817 12826 6851
rect 13804 6817 13838 6851
rect 11253 6749 11287 6783
rect 1547 6681 1581 6715
rect 5089 6613 5123 6647
rect 12863 6613 12897 6647
rect 1593 6409 1627 6443
rect 6009 6409 6043 6443
rect 8033 6409 8067 6443
rect 8401 6409 8435 6443
rect 11345 6409 11379 6443
rect 11713 6409 11747 6443
rect 12817 6409 12851 6443
rect 13829 6409 13863 6443
rect 6377 6341 6411 6375
rect 13277 6341 13311 6375
rect 7757 6273 7791 6307
rect 8585 6273 8619 6307
rect 10241 6273 10275 6307
rect 10885 6273 10919 6307
rect 9505 6205 9539 6239
rect 13093 6205 13127 6239
rect 8906 6137 8940 6171
rect 9873 6137 9907 6171
rect 10425 6137 10459 6171
rect 10517 6137 10551 6171
rect 5641 6069 5675 6103
rect 8953 5865 8987 5899
rect 10057 5865 10091 5899
rect 12863 5865 12897 5899
rect 13185 5865 13219 5899
rect 10333 5797 10367 5831
rect 10885 5797 10919 5831
rect 8493 5729 8527 5763
rect 12760 5729 12794 5763
rect 10241 5661 10275 5695
rect 11713 5661 11747 5695
rect 8677 5593 8711 5627
rect 8309 5321 8343 5355
rect 9505 5321 9539 5355
rect 12725 5321 12759 5355
rect 10057 5185 10091 5219
rect 10333 5185 10367 5219
rect 7941 5049 7975 5083
rect 8493 5049 8527 5083
rect 8585 5049 8619 5083
rect 9137 5049 9171 5083
rect 10149 5049 10183 5083
rect 9781 4981 9815 5015
rect 11069 4981 11103 5015
rect 8723 4777 8757 4811
rect 10057 4709 10091 4743
rect 11437 4709 11471 4743
rect 8585 4641 8619 4675
rect 11529 4641 11563 4675
rect 8493 4573 8527 4607
rect 9965 4573 9999 4607
rect 10241 4573 10275 4607
rect 8677 4233 8711 4267
rect 9229 4233 9263 4267
rect 10241 4233 10275 4267
rect 11529 4233 11563 4267
rect 9781 4097 9815 4131
rect 10425 4097 10459 4131
rect 10885 4097 10919 4131
rect 9321 4029 9355 4063
rect 20244 4029 20278 4063
rect 10517 3961 10551 3995
rect 9459 3893 9493 3927
rect 20315 3893 20349 3927
rect 20729 3893 20763 3927
rect 9413 3689 9447 3723
rect 10793 3689 10827 3723
rect 9689 3621 9723 3655
rect 9781 3553 9815 3587
rect 8769 3145 8803 3179
rect 9781 3145 9815 3179
rect 11437 3145 11471 3179
rect 8861 2941 8895 2975
rect 11044 2941 11078 2975
rect 9045 2805 9079 2839
rect 11115 2805 11149 2839
rect 4491 2601 4525 2635
rect 5503 2601 5537 2635
rect 10977 2601 11011 2635
rect 12771 2601 12805 2635
rect 19395 2601 19429 2635
rect 4420 2465 4454 2499
rect 4813 2465 4847 2499
rect 5432 2465 5466 2499
rect 10333 2465 10367 2499
rect 12700 2465 12734 2499
rect 13829 2465 13863 2499
rect 14381 2465 14415 2499
rect 15761 2465 15795 2499
rect 16865 2465 16899 2499
rect 17417 2465 17451 2499
rect 19324 2465 19358 2499
rect 22753 2465 22787 2499
rect 23305 2465 23339 2499
rect 24593 2465 24627 2499
rect 25145 2465 25179 2499
rect 16405 2397 16439 2431
rect 19809 2397 19843 2431
rect 14013 2329 14047 2363
rect 15945 2329 15979 2363
rect 22937 2329 22971 2363
rect 5917 2261 5951 2295
rect 10517 2261 10551 2295
rect 13185 2261 13219 2295
rect 17049 2261 17083 2295
rect 24777 2261 24811 2295
<< metal1 >>
rect 13446 27480 13452 27532
rect 13504 27520 13510 27532
rect 14734 27520 14740 27532
rect 13504 27492 14740 27520
rect 13504 27480 13510 27492
rect 14734 27480 14740 27492
rect 14792 27480 14798 27532
rect 15286 27480 15292 27532
rect 15344 27520 15350 27532
rect 26418 27520 26424 27532
rect 15344 27492 26424 27520
rect 15344 27480 15350 27492
rect 26418 27480 26424 27492
rect 26476 27480 26482 27532
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 11422 25344 11428 25356
rect 11383 25316 11428 25344
rect 11422 25304 11428 25316
rect 11480 25304 11486 25356
rect 13240 25347 13298 25353
rect 13240 25313 13252 25347
rect 13286 25344 13298 25347
rect 13538 25344 13544 25356
rect 13286 25316 13544 25344
rect 13286 25313 13298 25316
rect 13240 25307 13298 25313
rect 13538 25304 13544 25316
rect 13596 25304 13602 25356
rect 14252 25347 14310 25353
rect 14252 25313 14264 25347
rect 14298 25344 14310 25347
rect 14550 25344 14556 25356
rect 14298 25316 14556 25344
rect 14298 25313 14310 25316
rect 14252 25307 14310 25313
rect 14550 25304 14556 25316
rect 14608 25344 14614 25356
rect 15378 25344 15384 25356
rect 14608 25316 15384 25344
rect 14608 25304 14614 25316
rect 15378 25304 15384 25316
rect 15436 25304 15442 25356
rect 10413 25279 10471 25285
rect 10413 25245 10425 25279
rect 10459 25276 10471 25279
rect 11330 25276 11336 25288
rect 10459 25248 11336 25276
rect 10459 25245 10471 25248
rect 10413 25239 10471 25245
rect 11330 25236 11336 25248
rect 11388 25236 11394 25288
rect 12986 25168 12992 25220
rect 13044 25208 13050 25220
rect 14323 25211 14381 25217
rect 14323 25208 14335 25211
rect 13044 25180 14335 25208
rect 13044 25168 13050 25180
rect 14323 25177 14335 25180
rect 14369 25177 14381 25211
rect 14323 25171 14381 25177
rect 10778 25100 10784 25152
rect 10836 25140 10842 25152
rect 11563 25143 11621 25149
rect 11563 25140 11575 25143
rect 10836 25112 11575 25140
rect 10836 25100 10842 25112
rect 11563 25109 11575 25112
rect 11609 25109 11621 25143
rect 11563 25103 11621 25109
rect 12618 25100 12624 25152
rect 12676 25140 12682 25152
rect 13311 25143 13369 25149
rect 13311 25140 13323 25143
rect 12676 25112 13323 25140
rect 12676 25100 12682 25112
rect 13311 25109 13323 25112
rect 13357 25109 13369 25143
rect 13311 25103 13369 25109
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 10778 24936 10784 24948
rect 10739 24908 10784 24936
rect 10778 24896 10784 24908
rect 10836 24896 10842 24948
rect 11054 24936 11060 24948
rect 11015 24908 11060 24936
rect 11054 24896 11060 24908
rect 11112 24896 11118 24948
rect 14550 24936 14556 24948
rect 14511 24908 14556 24936
rect 14550 24896 14556 24908
rect 14608 24896 14614 24948
rect 14921 24939 14979 24945
rect 14921 24905 14933 24939
rect 14967 24936 14979 24939
rect 15286 24936 15292 24948
rect 14967 24908 15292 24936
rect 14967 24905 14979 24908
rect 14921 24899 14979 24905
rect 10413 24871 10471 24877
rect 10413 24837 10425 24871
rect 10459 24868 10471 24871
rect 11698 24868 11704 24880
rect 10459 24840 11704 24868
rect 10459 24837 10471 24840
rect 10413 24831 10471 24837
rect 8916 24735 8974 24741
rect 8916 24701 8928 24735
rect 8962 24732 8974 24735
rect 9912 24735 9970 24741
rect 8962 24704 9352 24732
rect 8962 24701 8974 24704
rect 8916 24695 8974 24701
rect 9324 24608 9352 24704
rect 9912 24701 9924 24735
rect 9958 24732 9970 24735
rect 10428 24732 10456 24831
rect 11698 24828 11704 24840
rect 11756 24868 11762 24880
rect 14090 24868 14096 24880
rect 11756 24840 14096 24868
rect 11756 24828 11762 24840
rect 14090 24828 14096 24840
rect 14148 24868 14154 24880
rect 14458 24868 14464 24880
rect 14148 24840 14464 24868
rect 14148 24828 14154 24840
rect 14458 24828 14464 24840
rect 14516 24828 14522 24880
rect 11885 24803 11943 24809
rect 11885 24769 11897 24803
rect 11931 24800 11943 24803
rect 13078 24800 13084 24812
rect 11931 24772 13084 24800
rect 11931 24769 11943 24772
rect 11885 24763 11943 24769
rect 9958 24704 10456 24732
rect 9958 24701 9970 24704
rect 9912 24695 9970 24701
rect 10778 24692 10784 24744
rect 10836 24732 10842 24744
rect 10873 24735 10931 24741
rect 10873 24732 10885 24735
rect 10836 24704 10885 24732
rect 10836 24692 10842 24704
rect 10873 24701 10885 24704
rect 10919 24701 10931 24735
rect 10873 24695 10931 24701
rect 11422 24692 11428 24744
rect 11480 24732 11486 24744
rect 11517 24735 11575 24741
rect 11517 24732 11529 24735
rect 11480 24704 11529 24732
rect 11480 24692 11486 24704
rect 11517 24701 11529 24704
rect 11563 24732 11575 24735
rect 12342 24732 12348 24744
rect 11563 24704 12348 24732
rect 11563 24701 11575 24704
rect 11517 24695 11575 24701
rect 12342 24692 12348 24704
rect 12400 24692 12406 24744
rect 12728 24741 12756 24772
rect 13078 24760 13084 24772
rect 13136 24760 13142 24812
rect 13538 24800 13544 24812
rect 13499 24772 13544 24800
rect 13538 24760 13544 24772
rect 13596 24760 13602 24812
rect 12713 24735 12771 24741
rect 12713 24701 12725 24735
rect 12759 24701 12771 24735
rect 12713 24695 12771 24701
rect 12897 24735 12955 24741
rect 12897 24701 12909 24735
rect 12943 24701 12955 24735
rect 12897 24695 12955 24701
rect 14068 24735 14126 24741
rect 14068 24701 14080 24735
rect 14114 24732 14126 24735
rect 14936 24732 14964 24899
rect 15286 24896 15292 24908
rect 15344 24896 15350 24948
rect 14114 24704 14964 24732
rect 14114 24701 14126 24704
rect 14068 24695 14126 24701
rect 9999 24667 10057 24673
rect 9999 24633 10011 24667
rect 10045 24664 10057 24667
rect 11238 24664 11244 24676
rect 10045 24636 11244 24664
rect 10045 24633 10057 24636
rect 9999 24627 10057 24633
rect 11238 24624 11244 24636
rect 11296 24624 11302 24676
rect 12912 24664 12940 24695
rect 12176 24636 12940 24664
rect 8987 24599 9045 24605
rect 8987 24565 8999 24599
rect 9033 24596 9045 24599
rect 9214 24596 9220 24608
rect 9033 24568 9220 24596
rect 9033 24565 9045 24568
rect 8987 24559 9045 24565
rect 9214 24556 9220 24568
rect 9272 24556 9278 24608
rect 9306 24556 9312 24608
rect 9364 24596 9370 24608
rect 9364 24568 9409 24596
rect 9364 24556 9370 24568
rect 12066 24556 12072 24608
rect 12124 24596 12130 24608
rect 12176 24605 12204 24636
rect 12161 24599 12219 24605
rect 12161 24596 12173 24599
rect 12124 24568 12173 24596
rect 12124 24556 12130 24568
rect 12161 24565 12173 24568
rect 12207 24565 12219 24599
rect 12710 24596 12716 24608
rect 12671 24568 12716 24596
rect 12161 24559 12219 24565
rect 12710 24556 12716 24568
rect 12768 24556 12774 24608
rect 14139 24599 14197 24605
rect 14139 24565 14151 24599
rect 14185 24596 14197 24599
rect 14274 24596 14280 24608
rect 14185 24568 14280 24596
rect 14185 24565 14197 24568
rect 14139 24559 14197 24565
rect 14274 24556 14280 24568
rect 14332 24556 14338 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 5442 24352 5448 24404
rect 5500 24392 5506 24404
rect 6454 24392 6460 24404
rect 5500 24364 6460 24392
rect 5500 24352 5506 24364
rect 6454 24352 6460 24364
rect 6512 24352 6518 24404
rect 9214 24352 9220 24404
rect 9272 24392 9278 24404
rect 9674 24392 9680 24404
rect 9272 24364 9680 24392
rect 9272 24352 9278 24364
rect 9674 24352 9680 24364
rect 9732 24392 9738 24404
rect 9861 24395 9919 24401
rect 9861 24392 9873 24395
rect 9732 24364 9873 24392
rect 9732 24352 9738 24364
rect 9861 24361 9873 24364
rect 9907 24361 9919 24395
rect 9861 24355 9919 24361
rect 11425 24395 11483 24401
rect 11425 24361 11437 24395
rect 11471 24392 11483 24395
rect 12434 24392 12440 24404
rect 11471 24364 12440 24392
rect 11471 24361 11483 24364
rect 11425 24355 11483 24361
rect 12434 24352 12440 24364
rect 12492 24352 12498 24404
rect 14277 24395 14335 24401
rect 14277 24361 14289 24395
rect 14323 24392 14335 24395
rect 23382 24392 23388 24404
rect 14323 24364 23388 24392
rect 14323 24361 14335 24364
rect 14277 24355 14335 24361
rect 23382 24352 23388 24364
rect 23440 24352 23446 24404
rect 12618 24324 12624 24336
rect 12579 24296 12624 24324
rect 12618 24284 12624 24296
rect 12676 24284 12682 24336
rect 12713 24327 12771 24333
rect 12713 24293 12725 24327
rect 12759 24324 12771 24327
rect 12802 24324 12808 24336
rect 12759 24296 12808 24324
rect 12759 24293 12771 24296
rect 12713 24287 12771 24293
rect 12802 24284 12808 24296
rect 12860 24284 12866 24336
rect 1210 24216 1216 24268
rect 1268 24256 1274 24268
rect 1432 24259 1490 24265
rect 1432 24256 1444 24259
rect 1268 24228 1444 24256
rect 1268 24216 1274 24228
rect 1432 24225 1444 24228
rect 1478 24225 1490 24259
rect 1432 24219 1490 24225
rect 5350 24216 5356 24268
rect 5408 24256 5414 24268
rect 8608 24259 8666 24265
rect 8608 24256 8620 24259
rect 5408 24228 8620 24256
rect 5408 24216 5414 24228
rect 8608 24225 8620 24228
rect 8654 24256 8666 24259
rect 8938 24256 8944 24268
rect 8654 24228 8944 24256
rect 8654 24225 8666 24228
rect 8608 24219 8666 24225
rect 8938 24216 8944 24228
rect 8996 24216 9002 24268
rect 10137 24259 10195 24265
rect 10137 24225 10149 24259
rect 10183 24256 10195 24259
rect 10318 24256 10324 24268
rect 10183 24228 10324 24256
rect 10183 24225 10195 24228
rect 10137 24219 10195 24225
rect 10318 24216 10324 24228
rect 10376 24216 10382 24268
rect 14090 24256 14096 24268
rect 14051 24228 14096 24256
rect 14090 24216 14096 24228
rect 14148 24216 14154 24268
rect 10781 24191 10839 24197
rect 10781 24188 10793 24191
rect 4126 24160 10793 24188
rect 1535 24123 1593 24129
rect 1535 24089 1547 24123
rect 1581 24120 1593 24123
rect 4126 24120 4154 24160
rect 10781 24157 10793 24160
rect 10827 24188 10839 24191
rect 10870 24188 10876 24200
rect 10827 24160 10876 24188
rect 10827 24157 10839 24160
rect 10781 24151 10839 24157
rect 10870 24148 10876 24160
rect 10928 24148 10934 24200
rect 12894 24188 12900 24200
rect 12855 24160 12900 24188
rect 12894 24148 12900 24160
rect 12952 24148 12958 24200
rect 1581 24092 4154 24120
rect 10367 24123 10425 24129
rect 1581 24089 1593 24092
rect 1535 24083 1593 24089
rect 10367 24089 10379 24123
rect 10413 24120 10425 24123
rect 12345 24123 12403 24129
rect 12345 24120 12357 24123
rect 10413 24092 12357 24120
rect 10413 24089 10425 24092
rect 10367 24083 10425 24089
rect 12345 24089 12357 24092
rect 12391 24120 12403 24123
rect 12526 24120 12532 24132
rect 12391 24092 12532 24120
rect 12391 24089 12403 24092
rect 12345 24083 12403 24089
rect 12526 24080 12532 24092
rect 12584 24080 12590 24132
rect 8386 24012 8392 24064
rect 8444 24052 8450 24064
rect 8711 24055 8769 24061
rect 8711 24052 8723 24055
rect 8444 24024 8723 24052
rect 8444 24012 8450 24024
rect 8711 24021 8723 24024
rect 8757 24021 8769 24055
rect 8711 24015 8769 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1210 23808 1216 23860
rect 1268 23848 1274 23860
rect 1857 23851 1915 23857
rect 1857 23848 1869 23851
rect 1268 23820 1869 23848
rect 1268 23808 1274 23820
rect 1857 23817 1869 23820
rect 1903 23817 1915 23851
rect 8938 23848 8944 23860
rect 8899 23820 8944 23848
rect 1857 23811 1915 23817
rect 8938 23808 8944 23820
rect 8996 23808 9002 23860
rect 9861 23851 9919 23857
rect 9861 23817 9873 23851
rect 9907 23848 9919 23851
rect 10134 23848 10140 23860
rect 9907 23820 10140 23848
rect 9907 23817 9919 23820
rect 9861 23811 9919 23817
rect 10134 23808 10140 23820
rect 10192 23808 10198 23860
rect 10318 23848 10324 23860
rect 10231 23820 10324 23848
rect 10318 23808 10324 23820
rect 10376 23848 10382 23860
rect 11974 23848 11980 23860
rect 10376 23820 11980 23848
rect 10376 23808 10382 23820
rect 11974 23808 11980 23820
rect 12032 23808 12038 23860
rect 15749 23851 15807 23857
rect 12912 23820 14412 23848
rect 12912 23792 12940 23820
rect 7193 23783 7251 23789
rect 7193 23749 7205 23783
rect 7239 23780 7251 23783
rect 9030 23780 9036 23792
rect 7239 23752 9036 23780
rect 7239 23749 7251 23752
rect 7193 23743 7251 23749
rect 9030 23740 9036 23752
rect 9088 23740 9094 23792
rect 11425 23783 11483 23789
rect 11425 23749 11437 23783
rect 11471 23780 11483 23783
rect 12894 23780 12900 23792
rect 11471 23752 12900 23780
rect 11471 23749 11483 23752
rect 11425 23743 11483 23749
rect 12894 23740 12900 23752
rect 12952 23740 12958 23792
rect 13541 23783 13599 23789
rect 13541 23749 13553 23783
rect 13587 23780 13599 23783
rect 13909 23783 13967 23789
rect 13587 23752 13814 23780
rect 13587 23749 13599 23752
rect 13541 23743 13599 23749
rect 10870 23712 10876 23724
rect 10831 23684 10876 23712
rect 10870 23672 10876 23684
rect 10928 23672 10934 23724
rect 12526 23712 12532 23724
rect 12487 23684 12532 23712
rect 12526 23672 12532 23684
rect 12584 23672 12590 23724
rect 13786 23712 13814 23752
rect 13909 23749 13921 23783
rect 13955 23780 13967 23783
rect 13998 23780 14004 23792
rect 13955 23752 14004 23780
rect 13955 23749 13967 23752
rect 13909 23743 13967 23749
rect 13998 23740 14004 23752
rect 14056 23740 14062 23792
rect 14384 23724 14412 23820
rect 15749 23817 15761 23851
rect 15795 23848 15807 23851
rect 16390 23848 16396 23860
rect 15795 23820 16396 23848
rect 15795 23817 15807 23820
rect 15749 23811 15807 23817
rect 16390 23808 16396 23820
rect 16448 23808 16454 23860
rect 16853 23851 16911 23857
rect 16853 23817 16865 23851
rect 16899 23848 16911 23851
rect 17402 23848 17408 23860
rect 16899 23820 17408 23848
rect 16899 23817 16911 23820
rect 16853 23811 16911 23817
rect 17402 23808 17408 23820
rect 17460 23808 17466 23860
rect 18693 23851 18751 23857
rect 18693 23817 18705 23851
rect 18739 23848 18751 23851
rect 20438 23848 20444 23860
rect 18739 23820 20444 23848
rect 18739 23817 18751 23820
rect 18693 23811 18751 23817
rect 20438 23808 20444 23820
rect 20496 23808 20502 23860
rect 21361 23851 21419 23857
rect 21361 23817 21373 23851
rect 21407 23848 21419 23851
rect 24210 23848 24216 23860
rect 21407 23820 24216 23848
rect 21407 23817 21419 23820
rect 21361 23811 21419 23817
rect 24210 23808 24216 23820
rect 24268 23808 24274 23860
rect 20257 23783 20315 23789
rect 20257 23749 20269 23783
rect 20303 23780 20315 23783
rect 22370 23780 22376 23792
rect 20303 23752 22376 23780
rect 20303 23749 20315 23752
rect 20257 23743 20315 23749
rect 22370 23740 22376 23752
rect 22428 23740 22434 23792
rect 14093 23715 14151 23721
rect 14093 23712 14105 23715
rect 13786 23684 14105 23712
rect 14093 23681 14105 23684
rect 14139 23712 14151 23715
rect 14274 23712 14280 23724
rect 14139 23684 14280 23712
rect 14139 23681 14151 23684
rect 14093 23675 14151 23681
rect 14274 23672 14280 23684
rect 14332 23672 14338 23724
rect 14366 23672 14372 23724
rect 14424 23712 14430 23724
rect 14424 23684 14469 23712
rect 14424 23672 14430 23684
rect 14550 23672 14556 23724
rect 14608 23712 14614 23724
rect 14608 23684 15608 23712
rect 14608 23672 14614 23684
rect 1118 23604 1124 23656
rect 1176 23644 1182 23656
rect 1432 23647 1490 23653
rect 1432 23644 1444 23647
rect 1176 23616 1444 23644
rect 1176 23604 1182 23616
rect 1432 23613 1444 23616
rect 1478 23644 1490 23647
rect 2225 23647 2283 23653
rect 2225 23644 2237 23647
rect 1478 23616 2237 23644
rect 1478 23613 1490 23616
rect 1432 23607 1490 23613
rect 2225 23613 2237 23616
rect 2271 23613 2283 23647
rect 2225 23607 2283 23613
rect 2460 23647 2518 23653
rect 2460 23613 2472 23647
rect 2506 23644 2518 23647
rect 2682 23644 2688 23656
rect 2506 23616 2688 23644
rect 2506 23613 2518 23616
rect 2460 23607 2518 23613
rect 2682 23604 2688 23616
rect 2740 23644 2746 23656
rect 2869 23647 2927 23653
rect 2869 23644 2881 23647
rect 2740 23616 2881 23644
rect 2740 23604 2746 23616
rect 2869 23613 2881 23616
rect 2915 23613 2927 23647
rect 2869 23607 2927 23613
rect 3488 23647 3546 23653
rect 3488 23613 3500 23647
rect 3534 23644 3546 23647
rect 3694 23644 3700 23656
rect 3534 23616 3700 23644
rect 3534 23613 3546 23616
rect 3488 23607 3546 23613
rect 3694 23604 3700 23616
rect 3752 23644 3758 23656
rect 3881 23647 3939 23653
rect 3881 23644 3893 23647
rect 3752 23616 3893 23644
rect 3752 23604 3758 23616
rect 3881 23613 3893 23616
rect 3927 23613 3939 23647
rect 3881 23607 3939 23613
rect 4430 23604 4436 23656
rect 4488 23644 4494 23656
rect 4652 23647 4710 23653
rect 4652 23644 4664 23647
rect 4488 23616 4664 23644
rect 4488 23604 4494 23616
rect 4652 23613 4664 23616
rect 4698 23644 4710 23647
rect 5077 23647 5135 23653
rect 5077 23644 5089 23647
rect 4698 23616 5089 23644
rect 4698 23613 4710 23616
rect 4652 23607 4710 23613
rect 5077 23613 5089 23616
rect 5123 23613 5135 23647
rect 7006 23644 7012 23656
rect 6919 23616 7012 23644
rect 5077 23607 5135 23613
rect 7006 23604 7012 23616
rect 7064 23644 7070 23656
rect 7561 23647 7619 23653
rect 7561 23644 7573 23647
rect 7064 23616 7573 23644
rect 7064 23604 7070 23616
rect 7561 23613 7573 23616
rect 7607 23613 7619 23647
rect 7561 23607 7619 23613
rect 8548 23647 8606 23653
rect 8548 23613 8560 23647
rect 8594 23644 8606 23647
rect 9398 23644 9404 23656
rect 8594 23616 9404 23644
rect 8594 23613 8606 23616
rect 8548 23607 8606 23613
rect 9398 23604 9404 23616
rect 9456 23604 9462 23656
rect 9674 23644 9680 23656
rect 9635 23616 9680 23644
rect 9674 23604 9680 23616
rect 9732 23604 9738 23656
rect 15580 23653 15608 23684
rect 18598 23672 18604 23724
rect 18656 23712 18662 23724
rect 18656 23684 20116 23712
rect 18656 23672 18662 23684
rect 15565 23647 15623 23653
rect 15565 23613 15577 23647
rect 15611 23644 15623 23647
rect 16117 23647 16175 23653
rect 16117 23644 16129 23647
rect 15611 23616 16129 23644
rect 15611 23613 15623 23616
rect 15565 23607 15623 23613
rect 16117 23613 16129 23616
rect 16163 23613 16175 23647
rect 16117 23607 16175 23613
rect 16669 23647 16727 23653
rect 16669 23613 16681 23647
rect 16715 23644 16727 23647
rect 17221 23647 17279 23653
rect 17221 23644 17233 23647
rect 16715 23616 17233 23644
rect 16715 23613 16727 23616
rect 16669 23607 16727 23613
rect 17221 23613 17233 23616
rect 17267 23644 17279 23647
rect 17310 23644 17316 23656
rect 17267 23616 17316 23644
rect 17267 23613 17279 23616
rect 17221 23607 17279 23613
rect 17310 23604 17316 23616
rect 17368 23604 17374 23656
rect 18506 23644 18512 23656
rect 18419 23616 18512 23644
rect 18506 23604 18512 23616
rect 18564 23644 18570 23656
rect 20088 23653 20116 23684
rect 19061 23647 19119 23653
rect 19061 23644 19073 23647
rect 18564 23616 19073 23644
rect 18564 23604 18570 23616
rect 19061 23613 19073 23616
rect 19107 23613 19119 23647
rect 19061 23607 19119 23613
rect 20073 23647 20131 23653
rect 20073 23613 20085 23647
rect 20119 23644 20131 23647
rect 20625 23647 20683 23653
rect 20625 23644 20637 23647
rect 20119 23616 20637 23644
rect 20119 23613 20131 23616
rect 20073 23607 20131 23613
rect 20625 23613 20637 23616
rect 20671 23613 20683 23647
rect 20625 23607 20683 23613
rect 21177 23647 21235 23653
rect 21177 23613 21189 23647
rect 21223 23613 21235 23647
rect 21177 23607 21235 23613
rect 2547 23579 2605 23585
rect 2547 23545 2559 23579
rect 2593 23576 2605 23579
rect 10965 23579 11023 23585
rect 2593 23548 3464 23576
rect 2593 23545 2605 23548
rect 2547 23539 2605 23545
rect 3436 23520 3464 23548
rect 10965 23545 10977 23579
rect 11011 23545 11023 23579
rect 10965 23539 11023 23545
rect 11885 23579 11943 23585
rect 11885 23545 11897 23579
rect 11931 23576 11943 23579
rect 12526 23576 12532 23588
rect 11931 23548 12532 23576
rect 11931 23545 11943 23548
rect 11885 23539 11943 23545
rect 1535 23511 1593 23517
rect 1535 23477 1547 23511
rect 1581 23508 1593 23511
rect 1670 23508 1676 23520
rect 1581 23480 1676 23508
rect 1581 23477 1593 23480
rect 1535 23471 1593 23477
rect 1670 23468 1676 23480
rect 1728 23468 1734 23520
rect 3418 23468 3424 23520
rect 3476 23468 3482 23520
rect 3559 23511 3617 23517
rect 3559 23477 3571 23511
rect 3605 23508 3617 23511
rect 3694 23508 3700 23520
rect 3605 23480 3700 23508
rect 3605 23477 3617 23480
rect 3559 23471 3617 23477
rect 3694 23468 3700 23480
rect 3752 23468 3758 23520
rect 4755 23511 4813 23517
rect 4755 23477 4767 23511
rect 4801 23508 4813 23511
rect 7098 23508 7104 23520
rect 4801 23480 7104 23508
rect 4801 23477 4813 23480
rect 4755 23471 4813 23477
rect 7098 23468 7104 23480
rect 7156 23468 7162 23520
rect 7926 23468 7932 23520
rect 7984 23508 7990 23520
rect 8619 23511 8677 23517
rect 8619 23508 8631 23511
rect 7984 23480 8631 23508
rect 7984 23468 7990 23480
rect 8619 23477 8631 23480
rect 8665 23477 8677 23511
rect 8619 23471 8677 23477
rect 10689 23511 10747 23517
rect 10689 23477 10701 23511
rect 10735 23508 10747 23511
rect 10980 23508 11008 23539
rect 12526 23536 12532 23548
rect 12584 23536 12590 23588
rect 12621 23579 12679 23585
rect 12621 23545 12633 23579
rect 12667 23545 12679 23579
rect 13170 23576 13176 23588
rect 13131 23548 13176 23576
rect 12621 23539 12679 23545
rect 11422 23508 11428 23520
rect 10735 23480 11428 23508
rect 10735 23477 10747 23480
rect 10689 23471 10747 23477
rect 11422 23468 11428 23480
rect 11480 23468 11486 23520
rect 12158 23468 12164 23520
rect 12216 23508 12222 23520
rect 12253 23511 12311 23517
rect 12253 23508 12265 23511
rect 12216 23480 12265 23508
rect 12216 23468 12222 23480
rect 12253 23477 12265 23480
rect 12299 23508 12311 23511
rect 12636 23508 12664 23539
rect 13170 23536 13176 23548
rect 13228 23536 13234 23588
rect 13786 23548 13952 23576
rect 13786 23508 13814 23548
rect 12299 23480 13814 23508
rect 13924 23508 13952 23548
rect 14182 23536 14188 23588
rect 14240 23576 14246 23588
rect 14240 23548 14285 23576
rect 14240 23536 14246 23548
rect 19978 23536 19984 23588
rect 20036 23576 20042 23588
rect 21192 23576 21220 23607
rect 21729 23579 21787 23585
rect 21729 23576 21741 23579
rect 20036 23548 21741 23576
rect 20036 23536 20042 23548
rect 21729 23545 21741 23548
rect 21775 23545 21787 23579
rect 21729 23539 21787 23545
rect 14200 23508 14228 23536
rect 13924 23480 14228 23508
rect 12299 23477 12311 23480
rect 12253 23471 12311 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 5307 23307 5365 23313
rect 5307 23273 5319 23307
rect 5353 23304 5365 23307
rect 7006 23304 7012 23316
rect 5353 23276 7012 23304
rect 5353 23273 5365 23276
rect 5307 23267 5365 23273
rect 7006 23264 7012 23276
rect 7064 23264 7070 23316
rect 7098 23264 7104 23316
rect 7156 23304 7162 23316
rect 7193 23307 7251 23313
rect 7193 23304 7205 23307
rect 7156 23276 7205 23304
rect 7156 23264 7162 23276
rect 7193 23273 7205 23276
rect 7239 23273 7251 23307
rect 7193 23267 7251 23273
rect 11238 23264 11244 23316
rect 11296 23304 11302 23316
rect 14090 23304 14096 23316
rect 11296 23276 12940 23304
rect 14051 23276 14096 23304
rect 11296 23264 11302 23276
rect 12912 23248 12940 23276
rect 14090 23264 14096 23276
rect 14148 23264 14154 23316
rect 14366 23304 14372 23316
rect 14327 23276 14372 23304
rect 14366 23264 14372 23276
rect 14424 23264 14430 23316
rect 15427 23307 15485 23313
rect 15427 23273 15439 23307
rect 15473 23304 15485 23307
rect 18598 23304 18604 23316
rect 15473 23276 18604 23304
rect 15473 23273 15485 23276
rect 15427 23267 15485 23273
rect 18598 23264 18604 23276
rect 18656 23264 18662 23316
rect 6362 23236 6368 23248
rect 6323 23208 6368 23236
rect 6362 23196 6368 23208
rect 6420 23196 6426 23248
rect 11330 23236 11336 23248
rect 11291 23208 11336 23236
rect 11330 23196 11336 23208
rect 11388 23196 11394 23248
rect 11422 23196 11428 23248
rect 11480 23236 11486 23248
rect 12894 23236 12900 23248
rect 11480 23208 11525 23236
rect 12807 23208 12900 23236
rect 11480 23196 11486 23208
rect 12894 23196 12900 23208
rect 12952 23196 12958 23248
rect 12989 23239 13047 23245
rect 12989 23205 13001 23239
rect 13035 23236 13047 23239
rect 13262 23236 13268 23248
rect 13035 23208 13268 23236
rect 13035 23205 13047 23208
rect 12989 23199 13047 23205
rect 13262 23196 13268 23208
rect 13320 23196 13326 23248
rect 4982 23128 4988 23180
rect 5040 23168 5046 23180
rect 5204 23171 5262 23177
rect 5204 23168 5216 23171
rect 5040 23140 5216 23168
rect 5040 23128 5046 23140
rect 5204 23137 5216 23140
rect 5250 23137 5262 23171
rect 5204 23131 5262 23137
rect 8478 23128 8484 23180
rect 8536 23168 8542 23180
rect 8608 23171 8666 23177
rect 8608 23168 8620 23171
rect 8536 23140 8620 23168
rect 8536 23128 8542 23140
rect 8608 23137 8620 23140
rect 8654 23137 8666 23171
rect 9766 23168 9772 23180
rect 9727 23140 9772 23168
rect 8608 23131 8666 23137
rect 9766 23128 9772 23140
rect 9824 23128 9830 23180
rect 9950 23128 9956 23180
rect 10008 23168 10014 23180
rect 10137 23171 10195 23177
rect 10137 23168 10149 23171
rect 10008 23140 10149 23168
rect 10008 23128 10014 23140
rect 10137 23137 10149 23140
rect 10183 23137 10195 23171
rect 10137 23131 10195 23137
rect 15356 23171 15414 23177
rect 15356 23137 15368 23171
rect 15402 23168 15414 23171
rect 16114 23168 16120 23180
rect 15402 23140 16120 23168
rect 15402 23137 15414 23140
rect 15356 23131 15414 23137
rect 16114 23128 16120 23140
rect 16172 23128 16178 23180
rect 6270 23100 6276 23112
rect 6231 23072 6276 23100
rect 6270 23060 6276 23072
rect 6328 23060 6334 23112
rect 6917 23103 6975 23109
rect 6917 23069 6929 23103
rect 6963 23100 6975 23103
rect 7190 23100 7196 23112
rect 6963 23072 7196 23100
rect 6963 23069 6975 23072
rect 6917 23063 6975 23069
rect 7190 23060 7196 23072
rect 7248 23060 7254 23112
rect 10413 23103 10471 23109
rect 10413 23069 10425 23103
rect 10459 23100 10471 23103
rect 11790 23100 11796 23112
rect 10459 23072 11796 23100
rect 10459 23069 10471 23072
rect 10413 23063 10471 23069
rect 11790 23060 11796 23072
rect 11848 23060 11854 23112
rect 11977 23103 12035 23109
rect 11977 23069 11989 23103
rect 12023 23100 12035 23103
rect 13170 23100 13176 23112
rect 12023 23072 13176 23100
rect 12023 23069 12035 23072
rect 11977 23063 12035 23069
rect 13170 23060 13176 23072
rect 13228 23060 13234 23112
rect 11057 23035 11115 23041
rect 11057 23032 11069 23035
rect 10336 23004 11069 23032
rect 10336 22976 10364 23004
rect 11057 23001 11069 23004
rect 11103 23001 11115 23035
rect 11057 22995 11115 23001
rect 8711 22967 8769 22973
rect 8711 22933 8723 22967
rect 8757 22964 8769 22967
rect 10318 22964 10324 22976
rect 8757 22936 10324 22964
rect 8757 22933 8769 22936
rect 8711 22927 8769 22933
rect 10318 22924 10324 22936
rect 10376 22924 10382 22976
rect 10778 22964 10784 22976
rect 10739 22936 10784 22964
rect 10778 22924 10784 22936
rect 10836 22964 10842 22976
rect 12529 22967 12587 22973
rect 12529 22964 12541 22967
rect 10836 22936 12541 22964
rect 10836 22924 10842 22936
rect 12529 22933 12541 22936
rect 12575 22964 12587 22967
rect 12802 22964 12808 22976
rect 12575 22936 12808 22964
rect 12575 22933 12587 22936
rect 12529 22927 12587 22933
rect 12802 22924 12808 22936
rect 12860 22964 12866 22976
rect 13262 22964 13268 22976
rect 12860 22936 13268 22964
rect 12860 22924 12866 22936
rect 13262 22924 13268 22936
rect 13320 22924 13326 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 3418 22720 3424 22772
rect 3476 22760 3482 22772
rect 5629 22763 5687 22769
rect 5629 22760 5641 22763
rect 3476 22732 5641 22760
rect 3476 22720 3482 22732
rect 5629 22729 5641 22732
rect 5675 22760 5687 22763
rect 6270 22760 6276 22772
rect 5675 22732 6276 22760
rect 5675 22729 5687 22732
rect 5629 22723 5687 22729
rect 6270 22720 6276 22732
rect 6328 22720 6334 22772
rect 6362 22720 6368 22772
rect 6420 22760 6426 22772
rect 6549 22763 6607 22769
rect 6549 22760 6561 22763
rect 6420 22732 6561 22760
rect 6420 22720 6426 22732
rect 6549 22729 6561 22732
rect 6595 22729 6607 22763
rect 8478 22760 8484 22772
rect 8439 22732 8484 22760
rect 6549 22723 6607 22729
rect 8478 22720 8484 22732
rect 8536 22720 8542 22772
rect 11330 22760 11336 22772
rect 11291 22732 11336 22760
rect 11330 22720 11336 22732
rect 11388 22720 11394 22772
rect 11422 22720 11428 22772
rect 11480 22760 11486 22772
rect 11609 22763 11667 22769
rect 11609 22760 11621 22763
rect 11480 22732 11621 22760
rect 11480 22720 11486 22732
rect 11609 22729 11621 22732
rect 11655 22729 11667 22763
rect 12618 22760 12624 22772
rect 12579 22732 12624 22760
rect 11609 22723 11667 22729
rect 12618 22720 12624 22732
rect 12676 22720 12682 22772
rect 13262 22720 13268 22772
rect 13320 22760 13326 22772
rect 13357 22763 13415 22769
rect 13357 22760 13369 22763
rect 13320 22732 13369 22760
rect 13320 22720 13326 22732
rect 13357 22729 13369 22732
rect 13403 22729 13415 22763
rect 16114 22760 16120 22772
rect 13357 22723 13415 22729
rect 14200 22732 16120 22760
rect 6181 22695 6239 22701
rect 6181 22661 6193 22695
rect 6227 22692 6239 22695
rect 8496 22692 8524 22720
rect 9766 22692 9772 22704
rect 6227 22664 8524 22692
rect 9679 22664 9772 22692
rect 6227 22661 6239 22664
rect 6181 22655 6239 22661
rect 5788 22559 5846 22565
rect 5788 22525 5800 22559
rect 5834 22556 5846 22559
rect 6196 22556 6224 22655
rect 9766 22652 9772 22664
rect 9824 22692 9830 22704
rect 11146 22692 11152 22704
rect 9824 22664 11152 22692
rect 9824 22652 9830 22664
rect 11146 22652 11152 22664
rect 11204 22652 11210 22704
rect 14090 22652 14096 22704
rect 14148 22692 14154 22704
rect 14200 22701 14228 22732
rect 16114 22720 16120 22732
rect 16172 22720 16178 22772
rect 18693 22763 18751 22769
rect 18693 22729 18705 22763
rect 18739 22760 18751 22763
rect 19426 22760 19432 22772
rect 18739 22732 19432 22760
rect 18739 22729 18751 22732
rect 18693 22723 18751 22729
rect 19426 22720 19432 22732
rect 19484 22720 19490 22772
rect 14185 22695 14243 22701
rect 14185 22692 14197 22695
rect 14148 22664 14197 22692
rect 14148 22652 14154 22664
rect 14185 22661 14197 22664
rect 14231 22661 14243 22695
rect 14185 22655 14243 22661
rect 6917 22627 6975 22633
rect 6917 22593 6929 22627
rect 6963 22624 6975 22627
rect 7098 22624 7104 22636
rect 6963 22596 7104 22624
rect 6963 22593 6975 22596
rect 6917 22587 6975 22593
rect 7098 22584 7104 22596
rect 7156 22584 7162 22636
rect 7190 22584 7196 22636
rect 7248 22624 7254 22636
rect 10318 22624 10324 22636
rect 7248 22596 7293 22624
rect 10279 22596 10324 22624
rect 7248 22584 7254 22596
rect 10318 22584 10324 22596
rect 10376 22584 10382 22636
rect 13633 22627 13691 22633
rect 13633 22593 13645 22627
rect 13679 22624 13691 22627
rect 14366 22624 14372 22636
rect 13679 22596 14372 22624
rect 13679 22593 13691 22596
rect 13633 22587 13691 22593
rect 14366 22584 14372 22596
rect 14424 22584 14430 22636
rect 8662 22556 8668 22568
rect 5834 22528 6224 22556
rect 8623 22528 8668 22556
rect 5834 22525 5846 22528
rect 5788 22519 5846 22525
rect 8662 22516 8668 22528
rect 8720 22516 8726 22568
rect 9217 22559 9275 22565
rect 9217 22525 9229 22559
rect 9263 22556 9275 22559
rect 9263 22528 9996 22556
rect 9263 22525 9275 22528
rect 9217 22519 9275 22525
rect 7006 22488 7012 22500
rect 6967 22460 7012 22488
rect 7006 22448 7012 22460
rect 7064 22448 7070 22500
rect 8205 22491 8263 22497
rect 8205 22457 8217 22491
rect 8251 22488 8263 22491
rect 9232 22488 9260 22519
rect 9398 22488 9404 22500
rect 8251 22460 9260 22488
rect 9359 22460 9404 22488
rect 8251 22457 8263 22460
rect 8205 22451 8263 22457
rect 9398 22448 9404 22460
rect 9456 22448 9462 22500
rect 9968 22432 9996 22528
rect 11974 22516 11980 22568
rect 12032 22556 12038 22568
rect 12437 22559 12495 22565
rect 12437 22556 12449 22559
rect 12032 22528 12449 22556
rect 12032 22516 12038 22528
rect 12437 22525 12449 22528
rect 12483 22556 12495 22559
rect 12989 22559 13047 22565
rect 12989 22556 13001 22559
rect 12483 22528 13001 22556
rect 12483 22525 12495 22528
rect 12437 22519 12495 22525
rect 12989 22525 13001 22528
rect 13035 22525 13047 22559
rect 15105 22559 15163 22565
rect 15105 22556 15117 22559
rect 12989 22519 13047 22525
rect 14568 22528 15117 22556
rect 10413 22491 10471 22497
rect 10413 22457 10425 22491
rect 10459 22488 10471 22491
rect 10778 22488 10784 22500
rect 10459 22460 10784 22488
rect 10459 22457 10471 22460
rect 10413 22451 10471 22457
rect 10778 22448 10784 22460
rect 10836 22448 10842 22500
rect 10962 22488 10968 22500
rect 10923 22460 10968 22488
rect 10962 22448 10968 22460
rect 11020 22448 11026 22500
rect 13722 22488 13728 22500
rect 13683 22460 13728 22488
rect 13722 22448 13728 22460
rect 13780 22448 13786 22500
rect 4982 22380 4988 22432
rect 5040 22420 5046 22432
rect 5169 22423 5227 22429
rect 5169 22420 5181 22423
rect 5040 22392 5181 22420
rect 5040 22380 5046 22392
rect 5169 22389 5181 22392
rect 5215 22389 5227 22423
rect 5169 22383 5227 22389
rect 5859 22423 5917 22429
rect 5859 22389 5871 22423
rect 5905 22420 5917 22423
rect 5994 22420 6000 22432
rect 5905 22392 6000 22420
rect 5905 22389 5917 22392
rect 5859 22383 5917 22389
rect 5994 22380 6000 22392
rect 6052 22380 6058 22432
rect 9950 22380 9956 22432
rect 10008 22420 10014 22432
rect 10045 22423 10103 22429
rect 10045 22420 10057 22423
rect 10008 22392 10057 22420
rect 10008 22380 10014 22392
rect 10045 22389 10057 22392
rect 10091 22389 10103 22423
rect 10045 22383 10103 22389
rect 13998 22380 14004 22432
rect 14056 22420 14062 22432
rect 14568 22429 14596 22528
rect 15105 22525 15117 22528
rect 15151 22556 15163 22559
rect 15470 22556 15476 22568
rect 15151 22528 15476 22556
rect 15151 22525 15163 22528
rect 15105 22519 15163 22525
rect 15470 22516 15476 22528
rect 15528 22516 15534 22568
rect 15565 22559 15623 22565
rect 15565 22525 15577 22559
rect 15611 22525 15623 22559
rect 15565 22519 15623 22525
rect 18509 22559 18567 22565
rect 18509 22525 18521 22559
rect 18555 22556 18567 22559
rect 18555 22528 19196 22556
rect 18555 22525 18567 22528
rect 18509 22519 18567 22525
rect 15580 22488 15608 22519
rect 14936 22460 15608 22488
rect 14936 22432 14964 22460
rect 19168 22432 19196 22528
rect 14553 22423 14611 22429
rect 14553 22420 14565 22423
rect 14056 22392 14565 22420
rect 14056 22380 14062 22392
rect 14553 22389 14565 22392
rect 14599 22389 14611 22423
rect 14918 22420 14924 22432
rect 14879 22392 14924 22420
rect 14553 22383 14611 22389
rect 14918 22380 14924 22392
rect 14976 22380 14982 22432
rect 15378 22420 15384 22432
rect 15339 22392 15384 22420
rect 15378 22380 15384 22392
rect 15436 22380 15442 22432
rect 19150 22420 19156 22432
rect 19111 22392 19156 22420
rect 19150 22380 19156 22392
rect 19208 22380 19214 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 6825 22219 6883 22225
rect 6825 22185 6837 22219
rect 6871 22216 6883 22219
rect 7006 22216 7012 22228
rect 6871 22188 7012 22216
rect 6871 22185 6883 22188
rect 6825 22179 6883 22185
rect 7006 22176 7012 22188
rect 7064 22176 7070 22228
rect 11422 22216 11428 22228
rect 10428 22188 11428 22216
rect 6362 22108 6368 22160
rect 6420 22148 6426 22160
rect 6914 22148 6920 22160
rect 6420 22120 6920 22148
rect 6420 22108 6426 22120
rect 6914 22108 6920 22120
rect 6972 22148 6978 22160
rect 7285 22151 7343 22157
rect 7285 22148 7297 22151
rect 6972 22120 7297 22148
rect 6972 22108 6978 22120
rect 7285 22117 7297 22120
rect 7331 22117 7343 22151
rect 7285 22111 7343 22117
rect 9766 22108 9772 22160
rect 9824 22148 9830 22160
rect 10428 22157 10456 22188
rect 11422 22176 11428 22188
rect 11480 22176 11486 22228
rect 11882 22216 11888 22228
rect 11843 22188 11888 22216
rect 11882 22176 11888 22188
rect 11940 22176 11946 22228
rect 12894 22216 12900 22228
rect 12855 22188 12900 22216
rect 12894 22176 12900 22188
rect 12952 22176 12958 22228
rect 13722 22176 13728 22228
rect 13780 22216 13786 22228
rect 14369 22219 14427 22225
rect 14369 22216 14381 22219
rect 13780 22188 14381 22216
rect 13780 22176 13786 22188
rect 14369 22185 14381 22188
rect 14415 22185 14427 22219
rect 14369 22179 14427 22185
rect 19150 22176 19156 22228
rect 19208 22216 19214 22228
rect 19291 22219 19349 22225
rect 19291 22216 19303 22219
rect 19208 22188 19303 22216
rect 19208 22176 19214 22188
rect 19291 22185 19303 22188
rect 19337 22185 19349 22219
rect 19291 22179 19349 22185
rect 10413 22151 10471 22157
rect 10413 22148 10425 22151
rect 9824 22120 10425 22148
rect 9824 22108 9830 22120
rect 10413 22117 10425 22120
rect 10459 22117 10471 22151
rect 10962 22148 10968 22160
rect 10923 22120 10968 22148
rect 10413 22111 10471 22117
rect 10962 22108 10968 22120
rect 11020 22148 11026 22160
rect 11514 22148 11520 22160
rect 11020 22120 11520 22148
rect 11020 22108 11026 22120
rect 11514 22108 11520 22120
rect 11572 22148 11578 22160
rect 11572 22120 12388 22148
rect 11572 22108 11578 22120
rect 14 22040 20 22092
rect 72 22080 78 22092
rect 2038 22080 2044 22092
rect 2096 22089 2102 22092
rect 2096 22083 2134 22089
rect 72 22052 2044 22080
rect 72 22040 78 22052
rect 2038 22040 2044 22052
rect 2122 22049 2134 22083
rect 2096 22043 2134 22049
rect 5144 22083 5202 22089
rect 5144 22049 5156 22083
rect 5190 22080 5202 22083
rect 5350 22080 5356 22092
rect 5190 22052 5356 22080
rect 5190 22049 5202 22052
rect 5144 22043 5202 22049
rect 2096 22040 2102 22043
rect 5350 22040 5356 22052
rect 5408 22040 5414 22092
rect 6089 22083 6147 22089
rect 6089 22049 6101 22083
rect 6135 22080 6147 22083
rect 6178 22080 6184 22092
rect 6135 22052 6184 22080
rect 6135 22049 6147 22052
rect 6089 22043 6147 22049
rect 6178 22040 6184 22052
rect 6236 22040 6242 22092
rect 11606 22040 11612 22092
rect 11664 22080 11670 22092
rect 11793 22083 11851 22089
rect 11793 22080 11805 22083
rect 11664 22052 11805 22080
rect 11664 22040 11670 22052
rect 11793 22049 11805 22052
rect 11839 22049 11851 22083
rect 11793 22043 11851 22049
rect 12066 22040 12072 22092
rect 12124 22080 12130 22092
rect 12250 22080 12256 22092
rect 12124 22052 12256 22080
rect 12124 22040 12130 22052
rect 12250 22040 12256 22052
rect 12308 22040 12314 22092
rect 12360 22080 12388 22120
rect 13170 22108 13176 22160
rect 13228 22148 13234 22160
rect 13449 22151 13507 22157
rect 13449 22148 13461 22151
rect 13228 22120 13461 22148
rect 13228 22108 13234 22120
rect 13449 22117 13461 22120
rect 13495 22117 13507 22151
rect 13449 22111 13507 22117
rect 13541 22151 13599 22157
rect 13541 22117 13553 22151
rect 13587 22148 13599 22151
rect 13630 22148 13636 22160
rect 13587 22120 13636 22148
rect 13587 22117 13599 22120
rect 13541 22111 13599 22117
rect 13630 22108 13636 22120
rect 13688 22108 13694 22160
rect 14090 22148 14096 22160
rect 14051 22120 14096 22148
rect 14090 22108 14096 22120
rect 14148 22108 14154 22160
rect 17402 22108 17408 22160
rect 17460 22148 17466 22160
rect 17773 22151 17831 22157
rect 17773 22148 17785 22151
rect 17460 22120 17785 22148
rect 17460 22108 17466 22120
rect 17773 22117 17785 22120
rect 17819 22117 17831 22151
rect 17773 22111 17831 22117
rect 13262 22080 13268 22092
rect 12360 22052 13268 22080
rect 13262 22040 13268 22052
rect 13320 22040 13326 22092
rect 15565 22083 15623 22089
rect 15565 22049 15577 22083
rect 15611 22080 15623 22083
rect 15838 22080 15844 22092
rect 15611 22052 15700 22080
rect 15799 22052 15844 22080
rect 15611 22049 15623 22052
rect 15565 22043 15623 22049
rect 5994 21972 6000 22024
rect 6052 22012 6058 22024
rect 7193 22015 7251 22021
rect 7193 22012 7205 22015
rect 6052 21984 7205 22012
rect 6052 21972 6058 21984
rect 7193 21981 7205 21984
rect 7239 21981 7251 22015
rect 7193 21975 7251 21981
rect 7282 21972 7288 22024
rect 7340 22012 7346 22024
rect 7837 22015 7895 22021
rect 7837 22012 7849 22015
rect 7340 21984 7849 22012
rect 7340 21972 7346 21984
rect 7837 21981 7849 21984
rect 7883 22012 7895 22015
rect 8938 22012 8944 22024
rect 7883 21984 8944 22012
rect 7883 21981 7895 21984
rect 7837 21975 7895 21981
rect 8938 21972 8944 21984
rect 8996 21972 9002 22024
rect 10321 22015 10379 22021
rect 10321 21981 10333 22015
rect 10367 22012 10379 22015
rect 10686 22012 10692 22024
rect 10367 21984 10692 22012
rect 10367 21981 10379 21984
rect 10321 21975 10379 21981
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 14918 22012 14924 22024
rect 13786 21984 14924 22012
rect 5534 21904 5540 21956
rect 5592 21944 5598 21956
rect 8662 21944 8668 21956
rect 5592 21916 8668 21944
rect 5592 21904 5598 21916
rect 8662 21904 8668 21916
rect 8720 21904 8726 21956
rect 12250 21904 12256 21956
rect 12308 21944 12314 21956
rect 13786 21944 13814 21984
rect 14918 21972 14924 21984
rect 14976 21972 14982 22024
rect 15672 21956 15700 22052
rect 15838 22040 15844 22052
rect 15896 22040 15902 22092
rect 18322 22040 18328 22092
rect 18380 22080 18386 22092
rect 19188 22083 19246 22089
rect 19188 22080 19200 22083
rect 18380 22052 19200 22080
rect 18380 22040 18386 22052
rect 19188 22049 19200 22052
rect 19234 22049 19246 22083
rect 19188 22043 19246 22049
rect 16022 22012 16028 22024
rect 15983 21984 16028 22012
rect 16022 21972 16028 21984
rect 16080 21972 16086 22024
rect 17678 22012 17684 22024
rect 17639 21984 17684 22012
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 15654 21944 15660 21956
rect 12308 21916 13814 21944
rect 15567 21916 15660 21944
rect 12308 21904 12314 21916
rect 15654 21904 15660 21916
rect 15712 21944 15718 21956
rect 15712 21916 16528 21944
rect 15712 21904 15718 21916
rect 16500 21888 16528 21916
rect 2179 21879 2237 21885
rect 2179 21845 2191 21879
rect 2225 21876 2237 21879
rect 2590 21876 2596 21888
rect 2225 21848 2596 21876
rect 2225 21845 2237 21848
rect 2179 21839 2237 21845
rect 2590 21836 2596 21848
rect 2648 21836 2654 21888
rect 4338 21876 4344 21888
rect 4299 21848 4344 21876
rect 4338 21836 4344 21848
rect 4396 21836 4402 21888
rect 5215 21879 5273 21885
rect 5215 21845 5227 21879
rect 5261 21876 5273 21879
rect 6086 21876 6092 21888
rect 5261 21848 6092 21876
rect 5261 21845 5273 21848
rect 5215 21839 5273 21845
rect 6086 21836 6092 21848
rect 6144 21836 6150 21888
rect 6227 21879 6285 21885
rect 6227 21845 6239 21879
rect 6273 21876 6285 21879
rect 6730 21876 6736 21888
rect 6273 21848 6736 21876
rect 6273 21845 6285 21848
rect 6227 21839 6285 21845
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 16482 21876 16488 21888
rect 16443 21848 16488 21876
rect 16482 21836 16488 21848
rect 16540 21836 16546 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2038 21672 2044 21684
rect 1999 21644 2044 21672
rect 2038 21632 2044 21644
rect 2096 21632 2102 21684
rect 5813 21675 5871 21681
rect 5813 21641 5825 21675
rect 5859 21672 5871 21675
rect 5994 21672 6000 21684
rect 5859 21644 6000 21672
rect 5859 21641 5871 21644
rect 5813 21635 5871 21641
rect 5994 21632 6000 21644
rect 6052 21632 6058 21684
rect 7006 21632 7012 21684
rect 7064 21672 7070 21684
rect 7745 21675 7803 21681
rect 7745 21672 7757 21675
rect 7064 21644 7757 21672
rect 7064 21632 7070 21644
rect 7745 21641 7757 21644
rect 7791 21672 7803 21675
rect 8018 21672 8024 21684
rect 7791 21644 8024 21672
rect 7791 21641 7803 21644
rect 7745 21635 7803 21641
rect 8018 21632 8024 21644
rect 8076 21672 8082 21684
rect 8389 21675 8447 21681
rect 8389 21672 8401 21675
rect 8076 21644 8401 21672
rect 8076 21632 8082 21644
rect 8389 21641 8401 21644
rect 8435 21641 8447 21675
rect 9766 21672 9772 21684
rect 9727 21644 9772 21672
rect 8389 21635 8447 21641
rect 9766 21632 9772 21644
rect 9824 21632 9830 21684
rect 10778 21632 10784 21684
rect 10836 21672 10842 21684
rect 11149 21675 11207 21681
rect 11149 21672 11161 21675
rect 10836 21644 11161 21672
rect 10836 21632 10842 21644
rect 11149 21641 11161 21644
rect 11195 21641 11207 21675
rect 11149 21635 11207 21641
rect 12713 21675 12771 21681
rect 12713 21641 12725 21675
rect 12759 21672 12771 21675
rect 13170 21672 13176 21684
rect 12759 21644 13176 21672
rect 12759 21641 12771 21644
rect 12713 21635 12771 21641
rect 13170 21632 13176 21644
rect 13228 21632 13234 21684
rect 13630 21632 13636 21684
rect 13688 21672 13694 21684
rect 14185 21675 14243 21681
rect 14185 21672 14197 21675
rect 13688 21644 14197 21672
rect 13688 21632 13694 21644
rect 14185 21641 14197 21644
rect 14231 21641 14243 21675
rect 14185 21635 14243 21641
rect 15470 21632 15476 21684
rect 15528 21672 15534 21684
rect 16209 21675 16267 21681
rect 16209 21672 16221 21675
rect 15528 21644 16221 21672
rect 15528 21632 15534 21644
rect 16209 21641 16221 21644
rect 16255 21641 16267 21675
rect 20162 21672 20168 21684
rect 20123 21644 20168 21672
rect 16209 21635 16267 21641
rect 5350 21604 5356 21616
rect 4126 21576 5356 21604
rect 2682 21496 2688 21548
rect 2740 21536 2746 21548
rect 4126 21536 4154 21576
rect 5350 21564 5356 21576
rect 5408 21604 5414 21616
rect 9674 21604 9680 21616
rect 5408 21576 9680 21604
rect 5408 21564 5414 21576
rect 9674 21564 9680 21576
rect 9732 21564 9738 21616
rect 11606 21564 11612 21616
rect 11664 21604 11670 21616
rect 14274 21604 14280 21616
rect 11664 21576 14280 21604
rect 11664 21564 11670 21576
rect 14274 21564 14280 21576
rect 14332 21564 14338 21616
rect 4338 21536 4344 21548
rect 2740 21508 4154 21536
rect 4299 21508 4344 21536
rect 2740 21496 2746 21508
rect 4338 21496 4344 21508
rect 4396 21496 4402 21548
rect 6086 21496 6092 21548
rect 6144 21536 6150 21548
rect 8665 21539 8723 21545
rect 8665 21536 8677 21539
rect 6144 21508 8677 21536
rect 6144 21496 6150 21508
rect 8665 21505 8677 21508
rect 8711 21536 8723 21539
rect 8846 21536 8852 21548
rect 8711 21508 8852 21536
rect 8711 21505 8723 21508
rect 8665 21499 8723 21505
rect 8846 21496 8852 21508
rect 8904 21496 8910 21548
rect 8938 21496 8944 21548
rect 8996 21536 9002 21548
rect 8996 21508 9041 21536
rect 8996 21496 9002 21508
rect 9950 21496 9956 21548
rect 10008 21536 10014 21548
rect 12161 21539 12219 21545
rect 12161 21536 12173 21539
rect 10008 21508 12173 21536
rect 10008 21496 10014 21508
rect 12161 21505 12173 21508
rect 12207 21536 12219 21539
rect 12250 21536 12256 21548
rect 12207 21508 12256 21536
rect 12207 21505 12219 21508
rect 12161 21499 12219 21505
rect 12250 21496 12256 21508
rect 12308 21496 12314 21548
rect 13262 21536 13268 21548
rect 13223 21508 13268 21536
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 13909 21539 13967 21545
rect 13909 21505 13921 21539
rect 13955 21536 13967 21539
rect 14090 21536 14096 21548
rect 13955 21508 14096 21536
rect 13955 21505 13967 21508
rect 13909 21499 13967 21505
rect 14090 21496 14096 21508
rect 14148 21496 14154 21548
rect 6825 21471 6883 21477
rect 6825 21437 6837 21471
rect 6871 21468 6883 21471
rect 6871 21440 8156 21468
rect 6871 21437 6883 21440
rect 6825 21431 6883 21437
rect 4433 21403 4491 21409
rect 4433 21369 4445 21403
rect 4479 21369 4491 21403
rect 4982 21400 4988 21412
rect 4943 21372 4988 21400
rect 4433 21363 4491 21369
rect 3970 21292 3976 21344
rect 4028 21332 4034 21344
rect 4065 21335 4123 21341
rect 4065 21332 4077 21335
rect 4028 21304 4077 21332
rect 4028 21292 4034 21304
rect 4065 21301 4077 21304
rect 4111 21332 4123 21335
rect 4448 21332 4476 21363
rect 4982 21360 4988 21372
rect 5040 21360 5046 21412
rect 6638 21400 6644 21412
rect 6551 21372 6644 21400
rect 6638 21360 6644 21372
rect 6696 21400 6702 21412
rect 7187 21403 7245 21409
rect 7187 21400 7199 21403
rect 6696 21372 7199 21400
rect 6696 21360 6702 21372
rect 7187 21369 7199 21372
rect 7233 21400 7245 21403
rect 7742 21400 7748 21412
rect 7233 21372 7748 21400
rect 7233 21369 7245 21372
rect 7187 21363 7245 21369
rect 7742 21360 7748 21372
rect 7800 21360 7806 21412
rect 8128 21409 8156 21440
rect 10042 21428 10048 21480
rect 10100 21468 10106 21480
rect 10229 21471 10287 21477
rect 10229 21468 10241 21471
rect 10100 21440 10241 21468
rect 10100 21428 10106 21440
rect 10229 21437 10241 21440
rect 10275 21437 10287 21471
rect 14918 21468 14924 21480
rect 14879 21440 14924 21468
rect 10229 21431 10287 21437
rect 14918 21428 14924 21440
rect 14976 21428 14982 21480
rect 15289 21471 15347 21477
rect 15289 21437 15301 21471
rect 15335 21437 15347 21471
rect 16224 21468 16252 21635
rect 20162 21632 20168 21644
rect 20220 21632 20226 21684
rect 24213 21675 24271 21681
rect 24213 21641 24225 21675
rect 24259 21672 24271 21675
rect 25406 21672 25412 21684
rect 24259 21644 25412 21672
rect 24259 21641 24271 21644
rect 24213 21635 24271 21641
rect 16393 21471 16451 21477
rect 16393 21468 16405 21471
rect 16224 21440 16405 21468
rect 15289 21431 15347 21437
rect 16393 21437 16405 21440
rect 16439 21437 16451 21471
rect 16393 21431 16451 21437
rect 8113 21403 8171 21409
rect 8113 21369 8125 21403
rect 8159 21400 8171 21403
rect 8478 21400 8484 21412
rect 8159 21372 8484 21400
rect 8159 21369 8171 21372
rect 8113 21363 8171 21369
rect 8478 21360 8484 21372
rect 8536 21360 8542 21412
rect 8757 21403 8815 21409
rect 8757 21369 8769 21403
rect 8803 21369 8815 21403
rect 10550 21403 10608 21409
rect 10550 21400 10562 21403
rect 8757 21363 8815 21369
rect 10152 21372 10562 21400
rect 4111 21304 4476 21332
rect 4111 21301 4123 21304
rect 4065 21295 4123 21301
rect 5074 21292 5080 21344
rect 5132 21332 5138 21344
rect 6089 21335 6147 21341
rect 6089 21332 6101 21335
rect 5132 21304 6101 21332
rect 5132 21292 5138 21304
rect 6089 21301 6101 21304
rect 6135 21332 6147 21335
rect 6178 21332 6184 21344
rect 6135 21304 6184 21332
rect 6135 21301 6147 21304
rect 6089 21295 6147 21301
rect 6178 21292 6184 21304
rect 6236 21292 6242 21344
rect 8018 21292 8024 21344
rect 8076 21332 8082 21344
rect 8772 21332 8800 21363
rect 10152 21344 10180 21372
rect 10550 21369 10562 21372
rect 10596 21369 10608 21403
rect 10550 21363 10608 21369
rect 13354 21360 13360 21412
rect 13412 21400 13418 21412
rect 15304 21400 15332 21431
rect 16482 21428 16488 21480
rect 16540 21468 16546 21480
rect 16853 21471 16911 21477
rect 16853 21468 16865 21471
rect 16540 21440 16865 21468
rect 16540 21428 16546 21440
rect 16853 21437 16865 21440
rect 16899 21437 16911 21471
rect 16853 21431 16911 21437
rect 19680 21471 19738 21477
rect 19680 21437 19692 21471
rect 19726 21468 19738 21471
rect 20162 21468 20168 21480
rect 19726 21440 20168 21468
rect 19726 21437 19738 21440
rect 19680 21431 19738 21437
rect 20162 21428 20168 21440
rect 20220 21428 20226 21480
rect 23728 21471 23786 21477
rect 23728 21437 23740 21471
rect 23774 21468 23786 21471
rect 24228 21468 24256 21635
rect 25406 21632 25412 21644
rect 25464 21632 25470 21684
rect 23774 21440 24256 21468
rect 23774 21437 23786 21440
rect 23728 21431 23786 21437
rect 15562 21400 15568 21412
rect 13412 21372 13457 21400
rect 14660 21372 15332 21400
rect 15523 21372 15568 21400
rect 13412 21360 13418 21372
rect 10134 21332 10140 21344
rect 8076 21304 8800 21332
rect 10095 21304 10140 21332
rect 8076 21292 8082 21304
rect 10134 21292 10140 21304
rect 10192 21292 10198 21344
rect 11606 21292 11612 21344
rect 11664 21332 11670 21344
rect 11793 21335 11851 21341
rect 11793 21332 11805 21335
rect 11664 21304 11805 21332
rect 11664 21292 11670 21304
rect 11793 21301 11805 21304
rect 11839 21301 11851 21335
rect 11793 21295 11851 21301
rect 13081 21335 13139 21341
rect 13081 21301 13093 21335
rect 13127 21332 13139 21335
rect 13372 21332 13400 21360
rect 13127 21304 13400 21332
rect 13127 21301 13139 21304
rect 13081 21295 13139 21301
rect 14274 21292 14280 21344
rect 14332 21332 14338 21344
rect 14660 21341 14688 21372
rect 15562 21360 15568 21372
rect 15620 21360 15626 21412
rect 15838 21360 15844 21412
rect 15896 21400 15902 21412
rect 15933 21403 15991 21409
rect 15933 21400 15945 21403
rect 15896 21372 15945 21400
rect 15896 21360 15902 21372
rect 15933 21369 15945 21372
rect 15979 21400 15991 21403
rect 17586 21400 17592 21412
rect 15979 21372 17592 21400
rect 15979 21369 15991 21372
rect 15933 21363 15991 21369
rect 17586 21360 17592 21372
rect 17644 21360 17650 21412
rect 18138 21400 18144 21412
rect 18099 21372 18144 21400
rect 18138 21360 18144 21372
rect 18196 21360 18202 21412
rect 18233 21403 18291 21409
rect 18233 21369 18245 21403
rect 18279 21369 18291 21403
rect 18233 21363 18291 21369
rect 14645 21335 14703 21341
rect 14645 21332 14657 21335
rect 14332 21304 14657 21332
rect 14332 21292 14338 21304
rect 14645 21301 14657 21304
rect 14691 21301 14703 21335
rect 16482 21332 16488 21344
rect 16443 21304 16488 21332
rect 14645 21295 14703 21301
rect 16482 21292 16488 21304
rect 16540 21292 16546 21344
rect 16942 21292 16948 21344
rect 17000 21332 17006 21344
rect 17402 21332 17408 21344
rect 17000 21304 17408 21332
rect 17000 21292 17006 21304
rect 17402 21292 17408 21304
rect 17460 21292 17466 21344
rect 17770 21332 17776 21344
rect 17731 21304 17776 21332
rect 17770 21292 17776 21304
rect 17828 21332 17834 21344
rect 18248 21332 18276 21363
rect 18322 21360 18328 21412
rect 18380 21400 18386 21412
rect 18785 21403 18843 21409
rect 18785 21400 18797 21403
rect 18380 21372 18797 21400
rect 18380 21360 18386 21372
rect 18785 21369 18797 21372
rect 18831 21400 18843 21403
rect 19245 21403 19303 21409
rect 19245 21400 19257 21403
rect 18831 21372 19257 21400
rect 18831 21369 18843 21372
rect 18785 21363 18843 21369
rect 19245 21369 19257 21372
rect 19291 21400 19303 21403
rect 20070 21400 20076 21412
rect 19291 21372 20076 21400
rect 19291 21369 19303 21372
rect 19245 21363 19303 21369
rect 20070 21360 20076 21372
rect 20128 21360 20134 21412
rect 17828 21304 18276 21332
rect 17828 21292 17834 21304
rect 19518 21292 19524 21344
rect 19576 21332 19582 21344
rect 19751 21335 19809 21341
rect 19751 21332 19763 21335
rect 19576 21304 19763 21332
rect 19576 21292 19582 21304
rect 19751 21301 19763 21304
rect 19797 21301 19809 21335
rect 19751 21295 19809 21301
rect 20530 21292 20536 21344
rect 20588 21332 20594 21344
rect 23799 21335 23857 21341
rect 23799 21332 23811 21335
rect 20588 21304 23811 21332
rect 20588 21292 20594 21304
rect 23799 21301 23811 21304
rect 23845 21301 23857 21335
rect 23799 21295 23857 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1578 21128 1584 21140
rect 1539 21100 1584 21128
rect 1578 21088 1584 21100
rect 1636 21088 1642 21140
rect 6914 21128 6920 21140
rect 6875 21100 6920 21128
rect 6914 21088 6920 21100
rect 6972 21128 6978 21140
rect 7193 21131 7251 21137
rect 7193 21128 7205 21131
rect 6972 21100 7205 21128
rect 6972 21088 6978 21100
rect 7193 21097 7205 21100
rect 7239 21097 7251 21131
rect 8846 21128 8852 21140
rect 8807 21100 8852 21128
rect 7193 21091 7251 21097
rect 8846 21088 8852 21100
rect 8904 21088 8910 21140
rect 9815 21131 9873 21137
rect 9815 21097 9827 21131
rect 9861 21128 9873 21131
rect 10686 21128 10692 21140
rect 9861 21100 10692 21128
rect 9861 21097 9873 21100
rect 9815 21091 9873 21097
rect 10686 21088 10692 21100
rect 10744 21088 10750 21140
rect 11330 21128 11336 21140
rect 11291 21100 11336 21128
rect 11330 21088 11336 21100
rect 11388 21088 11394 21140
rect 11885 21131 11943 21137
rect 11885 21097 11897 21131
rect 11931 21128 11943 21131
rect 12158 21128 12164 21140
rect 11931 21100 12164 21128
rect 11931 21097 11943 21100
rect 11885 21091 11943 21097
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 13722 21088 13728 21140
rect 13780 21128 13786 21140
rect 14001 21131 14059 21137
rect 14001 21128 14013 21131
rect 13780 21100 14013 21128
rect 13780 21088 13786 21100
rect 14001 21097 14013 21100
rect 14047 21097 14059 21131
rect 14918 21128 14924 21140
rect 14831 21100 14924 21128
rect 14001 21091 14059 21097
rect 14918 21088 14924 21100
rect 14976 21128 14982 21140
rect 15565 21131 15623 21137
rect 15565 21128 15577 21131
rect 14976 21100 15577 21128
rect 14976 21088 14982 21100
rect 15565 21097 15577 21100
rect 15611 21128 15623 21131
rect 15654 21128 15660 21140
rect 15611 21100 15660 21128
rect 15611 21097 15623 21100
rect 15565 21091 15623 21097
rect 15654 21088 15660 21100
rect 15712 21088 15718 21140
rect 16022 21128 16028 21140
rect 15983 21100 16028 21128
rect 16022 21088 16028 21100
rect 16080 21128 16086 21140
rect 16080 21100 16160 21128
rect 16080 21088 16086 21100
rect 4246 21060 4252 21072
rect 4207 21032 4252 21060
rect 4246 21020 4252 21032
rect 4304 21020 4310 21072
rect 6086 21020 6092 21072
rect 6144 21060 6150 21072
rect 6359 21063 6417 21069
rect 6359 21060 6371 21063
rect 6144 21032 6371 21060
rect 6144 21020 6150 21032
rect 6359 21029 6371 21032
rect 6405 21060 6417 21063
rect 6638 21060 6644 21072
rect 6405 21032 6644 21060
rect 6405 21029 6417 21032
rect 6359 21023 6417 21029
rect 6638 21020 6644 21032
rect 6696 21020 6702 21072
rect 7745 21063 7803 21069
rect 7745 21029 7757 21063
rect 7791 21060 7803 21063
rect 7926 21060 7932 21072
rect 7791 21032 7932 21060
rect 7791 21029 7803 21032
rect 7745 21023 7803 21029
rect 7926 21020 7932 21032
rect 7984 21020 7990 21072
rect 8018 21020 8024 21072
rect 8076 21060 8082 21072
rect 8076 21032 8121 21060
rect 8076 21020 8082 21032
rect 13170 21020 13176 21072
rect 13228 21060 13234 21072
rect 13402 21063 13460 21069
rect 13402 21060 13414 21063
rect 13228 21032 13414 21060
rect 13228 21020 13234 21032
rect 13402 21029 13414 21032
rect 13448 21029 13460 21063
rect 13402 21023 13460 21029
rect 1397 20995 1455 21001
rect 1397 20961 1409 20995
rect 1443 20992 1455 20995
rect 1762 20992 1768 21004
rect 1443 20964 1768 20992
rect 1443 20961 1455 20964
rect 1397 20955 1455 20961
rect 1762 20952 1768 20964
rect 1820 20952 1826 21004
rect 9585 20995 9643 21001
rect 9585 20961 9597 20995
rect 9631 20992 9643 20995
rect 9674 20992 9680 21004
rect 9631 20964 9680 20992
rect 9631 20961 9643 20964
rect 9585 20955 9643 20961
rect 9674 20952 9680 20964
rect 9732 20952 9738 21004
rect 10965 20995 11023 21001
rect 10965 20961 10977 20995
rect 11011 20992 11023 20995
rect 11882 20992 11888 21004
rect 11011 20964 11888 20992
rect 11011 20961 11023 20964
rect 10965 20955 11023 20961
rect 11882 20952 11888 20964
rect 11940 20952 11946 21004
rect 12894 20952 12900 21004
rect 12952 20992 12958 21004
rect 12989 20995 13047 21001
rect 12989 20992 13001 20995
rect 12952 20964 13001 20992
rect 12952 20952 12958 20964
rect 12989 20961 13001 20964
rect 13035 20992 13047 20995
rect 15378 20992 15384 21004
rect 13035 20964 15384 20992
rect 13035 20961 13047 20964
rect 12989 20955 13047 20961
rect 15378 20952 15384 20964
rect 15436 20952 15442 21004
rect 16132 21001 16160 21100
rect 16390 21088 16396 21140
rect 16448 21128 16454 21140
rect 16485 21131 16543 21137
rect 16485 21128 16497 21131
rect 16448 21100 16497 21128
rect 16448 21088 16454 21100
rect 16485 21097 16497 21100
rect 16531 21097 16543 21131
rect 16485 21091 16543 21097
rect 17037 21131 17095 21137
rect 17037 21097 17049 21131
rect 17083 21128 17095 21131
rect 17770 21128 17776 21140
rect 17083 21100 17776 21128
rect 17083 21097 17095 21100
rect 17037 21091 17095 21097
rect 17770 21088 17776 21100
rect 17828 21088 17834 21140
rect 19518 21088 19524 21140
rect 19576 21128 19582 21140
rect 19705 21131 19763 21137
rect 19705 21128 19717 21131
rect 19576 21100 19717 21128
rect 19576 21088 19582 21100
rect 19705 21097 19717 21100
rect 19751 21097 19763 21131
rect 19705 21091 19763 21097
rect 17678 21060 17684 21072
rect 17639 21032 17684 21060
rect 17678 21020 17684 21032
rect 17736 21020 17742 21072
rect 18877 21063 18935 21069
rect 18877 21029 18889 21063
rect 18923 21060 18935 21063
rect 18966 21060 18972 21072
rect 18923 21032 18972 21060
rect 18923 21029 18935 21032
rect 18877 21023 18935 21029
rect 18966 21020 18972 21032
rect 19024 21020 19030 21072
rect 16117 20995 16175 21001
rect 16117 20961 16129 20995
rect 16163 20961 16175 20995
rect 16117 20955 16175 20961
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20924 3019 20927
rect 3786 20924 3792 20936
rect 3007 20896 3792 20924
rect 3007 20893 3019 20896
rect 2961 20887 3019 20893
rect 3786 20884 3792 20896
rect 3844 20924 3850 20936
rect 4157 20927 4215 20933
rect 4157 20924 4169 20927
rect 3844 20896 4169 20924
rect 3844 20884 3850 20896
rect 4157 20893 4169 20896
rect 4203 20893 4215 20927
rect 4430 20924 4436 20936
rect 4391 20896 4436 20924
rect 4157 20887 4215 20893
rect 4430 20884 4436 20896
rect 4488 20884 4494 20936
rect 5994 20924 6000 20936
rect 5955 20896 6000 20924
rect 5994 20884 6000 20896
rect 6052 20884 6058 20936
rect 7650 20884 7656 20936
rect 7708 20924 7714 20936
rect 8205 20927 8263 20933
rect 8205 20924 8217 20927
rect 7708 20896 8217 20924
rect 7708 20884 7714 20896
rect 8205 20893 8217 20896
rect 8251 20893 8263 20927
rect 8205 20887 8263 20893
rect 11790 20884 11796 20936
rect 11848 20924 11854 20936
rect 13081 20927 13139 20933
rect 13081 20924 13093 20927
rect 11848 20896 13093 20924
rect 11848 20884 11854 20896
rect 13081 20893 13093 20896
rect 13127 20924 13139 20927
rect 14090 20924 14096 20936
rect 13127 20896 14096 20924
rect 13127 20893 13139 20896
rect 13081 20887 13139 20893
rect 14090 20884 14096 20896
rect 14148 20884 14154 20936
rect 18138 20884 18144 20936
rect 18196 20924 18202 20936
rect 18785 20927 18843 20933
rect 18196 20896 18552 20924
rect 18196 20884 18202 20896
rect 6178 20816 6184 20868
rect 6236 20856 6242 20868
rect 11606 20856 11612 20868
rect 6236 20828 11612 20856
rect 6236 20816 6242 20828
rect 11606 20816 11612 20828
rect 11664 20816 11670 20868
rect 18524 20865 18552 20896
rect 18785 20893 18797 20927
rect 18831 20924 18843 20927
rect 19242 20924 19248 20936
rect 18831 20896 19248 20924
rect 18831 20893 18843 20896
rect 18785 20887 18843 20893
rect 19242 20884 19248 20896
rect 19300 20924 19306 20936
rect 20530 20924 20536 20936
rect 19300 20896 20536 20924
rect 19300 20884 19306 20896
rect 20530 20884 20536 20896
rect 20588 20884 20594 20936
rect 18509 20859 18567 20865
rect 18509 20825 18521 20859
rect 18555 20856 18567 20859
rect 19337 20859 19395 20865
rect 19337 20856 19349 20859
rect 18555 20828 19349 20856
rect 18555 20825 18567 20828
rect 18509 20819 18567 20825
rect 19337 20825 19349 20828
rect 19383 20856 19395 20859
rect 20346 20856 20352 20868
rect 19383 20828 20352 20856
rect 19383 20825 19395 20828
rect 19337 20819 19395 20825
rect 20346 20816 20352 20828
rect 20404 20816 20410 20868
rect 4798 20748 4804 20800
rect 4856 20788 4862 20800
rect 5077 20791 5135 20797
rect 5077 20788 5089 20791
rect 4856 20760 5089 20788
rect 4856 20748 4862 20760
rect 5077 20757 5089 20760
rect 5123 20757 5135 20791
rect 5077 20751 5135 20757
rect 10042 20748 10048 20800
rect 10100 20788 10106 20800
rect 10229 20791 10287 20797
rect 10229 20788 10241 20791
rect 10100 20760 10241 20788
rect 10100 20748 10106 20760
rect 10229 20757 10241 20760
rect 10275 20757 10287 20791
rect 18138 20788 18144 20800
rect 18099 20760 18144 20788
rect 10229 20751 10287 20757
rect 18138 20748 18144 20760
rect 18196 20748 18202 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2590 20584 2596 20596
rect 2551 20556 2596 20584
rect 2590 20544 2596 20556
rect 2648 20584 2654 20596
rect 4246 20584 4252 20596
rect 2648 20556 3280 20584
rect 4207 20556 4252 20584
rect 2648 20544 2654 20556
rect 3252 20457 3280 20556
rect 4246 20544 4252 20556
rect 4304 20584 4310 20596
rect 4525 20587 4583 20593
rect 4525 20584 4537 20587
rect 4304 20556 4537 20584
rect 4304 20544 4310 20556
rect 4525 20553 4537 20556
rect 4571 20553 4583 20587
rect 6086 20584 6092 20596
rect 6047 20556 6092 20584
rect 4525 20547 4583 20553
rect 6086 20544 6092 20556
rect 6144 20544 6150 20596
rect 6641 20587 6699 20593
rect 6641 20553 6653 20587
rect 6687 20584 6699 20587
rect 6914 20584 6920 20596
rect 6687 20556 6920 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 6914 20544 6920 20556
rect 6972 20544 6978 20596
rect 9674 20584 9680 20596
rect 9635 20556 9680 20584
rect 9674 20544 9680 20556
rect 9732 20544 9738 20596
rect 11149 20587 11207 20593
rect 11149 20553 11161 20587
rect 11195 20584 11207 20587
rect 11422 20584 11428 20596
rect 11195 20556 11428 20584
rect 11195 20553 11207 20556
rect 11149 20547 11207 20553
rect 11422 20544 11428 20556
rect 11480 20544 11486 20596
rect 11882 20584 11888 20596
rect 11843 20556 11888 20584
rect 11882 20544 11888 20556
rect 11940 20544 11946 20596
rect 13630 20544 13636 20596
rect 13688 20584 13694 20596
rect 13817 20587 13875 20593
rect 13817 20584 13829 20587
rect 13688 20556 13829 20584
rect 13688 20544 13694 20556
rect 13817 20553 13829 20556
rect 13863 20553 13875 20587
rect 14090 20584 14096 20596
rect 14051 20556 14096 20584
rect 13817 20547 13875 20553
rect 14090 20544 14096 20556
rect 14148 20544 14154 20596
rect 4338 20476 4344 20528
rect 4396 20516 4402 20528
rect 4396 20488 5120 20516
rect 4396 20476 4402 20488
rect 3237 20451 3295 20457
rect 3237 20417 3249 20451
rect 3283 20417 3295 20451
rect 3237 20411 3295 20417
rect 3881 20451 3939 20457
rect 3881 20417 3893 20451
rect 3927 20448 3939 20451
rect 4430 20448 4436 20460
rect 3927 20420 4436 20448
rect 3927 20417 3939 20420
rect 3881 20411 3939 20417
rect 4430 20408 4436 20420
rect 4488 20408 4494 20460
rect 4798 20448 4804 20460
rect 4759 20420 4804 20448
rect 4798 20408 4804 20420
rect 4856 20408 4862 20460
rect 5092 20457 5120 20488
rect 17862 20476 17868 20528
rect 17920 20516 17926 20528
rect 20806 20516 20812 20528
rect 17920 20488 20812 20516
rect 17920 20476 17926 20488
rect 20806 20476 20812 20488
rect 20864 20476 20870 20528
rect 25130 20516 25136 20528
rect 25091 20488 25136 20516
rect 25130 20476 25136 20488
rect 25188 20476 25194 20528
rect 5077 20451 5135 20457
rect 5077 20417 5089 20451
rect 5123 20417 5135 20451
rect 5077 20411 5135 20417
rect 6730 20408 6736 20460
rect 6788 20448 6794 20460
rect 7009 20451 7067 20457
rect 7009 20448 7021 20451
rect 6788 20420 7021 20448
rect 6788 20408 6794 20420
rect 7009 20417 7021 20420
rect 7055 20417 7067 20451
rect 7650 20448 7656 20460
rect 7611 20420 7656 20448
rect 7009 20411 7067 20417
rect 7650 20408 7656 20420
rect 7708 20408 7714 20460
rect 9398 20408 9404 20460
rect 9456 20448 9462 20460
rect 10229 20451 10287 20457
rect 10229 20448 10241 20451
rect 9456 20420 10241 20448
rect 9456 20408 9462 20420
rect 10229 20417 10241 20420
rect 10275 20448 10287 20451
rect 10686 20448 10692 20460
rect 10275 20420 10692 20448
rect 10275 20417 10287 20420
rect 10229 20411 10287 20417
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 12894 20448 12900 20460
rect 12855 20420 12900 20448
rect 12894 20408 12900 20420
rect 12952 20408 12958 20460
rect 15562 20408 15568 20460
rect 15620 20448 15626 20460
rect 16117 20451 16175 20457
rect 16117 20448 16129 20451
rect 15620 20420 16129 20448
rect 15620 20408 15626 20420
rect 16117 20417 16129 20420
rect 16163 20448 16175 20451
rect 17313 20451 17371 20457
rect 17313 20448 17325 20451
rect 16163 20420 17325 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 17313 20417 17325 20420
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 17678 20408 17684 20460
rect 17736 20448 17742 20460
rect 18417 20451 18475 20457
rect 18417 20448 18429 20451
rect 17736 20420 18429 20448
rect 17736 20408 17742 20420
rect 18417 20417 18429 20420
rect 18463 20448 18475 20451
rect 18874 20448 18880 20460
rect 18463 20420 18880 20448
rect 18463 20417 18475 20420
rect 18417 20411 18475 20417
rect 18874 20408 18880 20420
rect 18932 20408 18938 20460
rect 19518 20408 19524 20460
rect 19576 20448 19582 20460
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 19576 20420 19717 20448
rect 19576 20408 19582 20420
rect 19705 20417 19717 20420
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 8389 20383 8447 20389
rect 8389 20349 8401 20383
rect 8435 20380 8447 20383
rect 8757 20383 8815 20389
rect 8757 20380 8769 20383
rect 8435 20352 8769 20380
rect 8435 20349 8447 20352
rect 8389 20343 8447 20349
rect 8757 20349 8769 20352
rect 8803 20380 8815 20383
rect 8846 20380 8852 20392
rect 8803 20352 8852 20380
rect 8803 20349 8815 20352
rect 8757 20343 8815 20349
rect 8846 20340 8852 20352
rect 8904 20340 8910 20392
rect 8941 20383 8999 20389
rect 8941 20349 8953 20383
rect 8987 20349 8999 20383
rect 8941 20343 8999 20349
rect 14712 20383 14770 20389
rect 14712 20349 14724 20383
rect 14758 20380 14770 20383
rect 15102 20380 15108 20392
rect 14758 20352 15108 20380
rect 14758 20349 14770 20352
rect 14712 20343 14770 20349
rect 3329 20315 3387 20321
rect 3329 20312 3341 20315
rect 2976 20284 3341 20312
rect 2976 20256 3004 20284
rect 3329 20281 3341 20284
rect 3375 20281 3387 20315
rect 3329 20275 3387 20281
rect 4893 20315 4951 20321
rect 4893 20281 4905 20315
rect 4939 20281 4951 20315
rect 4893 20275 4951 20281
rect 1673 20247 1731 20253
rect 1673 20213 1685 20247
rect 1719 20244 1731 20247
rect 1762 20244 1768 20256
rect 1719 20216 1768 20244
rect 1719 20213 1731 20216
rect 1673 20207 1731 20213
rect 1762 20204 1768 20216
rect 1820 20204 1826 20256
rect 2958 20244 2964 20256
rect 2919 20216 2964 20244
rect 2958 20204 2964 20216
rect 3016 20204 3022 20256
rect 3142 20204 3148 20256
rect 3200 20244 3206 20256
rect 4246 20244 4252 20256
rect 3200 20216 4252 20244
rect 3200 20204 3206 20216
rect 4246 20204 4252 20216
rect 4304 20244 4310 20256
rect 4908 20244 4936 20275
rect 7006 20272 7012 20324
rect 7064 20312 7070 20324
rect 7101 20315 7159 20321
rect 7101 20312 7113 20315
rect 7064 20284 7113 20312
rect 7064 20272 7070 20284
rect 7101 20281 7113 20284
rect 7147 20281 7159 20315
rect 8956 20312 8984 20343
rect 15102 20340 15108 20352
rect 15160 20340 15166 20392
rect 24648 20383 24706 20389
rect 24648 20349 24660 20383
rect 24694 20380 24706 20383
rect 25148 20380 25176 20476
rect 24694 20352 25176 20380
rect 24694 20349 24706 20352
rect 24648 20343 24706 20349
rect 10134 20312 10140 20324
rect 7101 20275 7159 20281
rect 7944 20284 8984 20312
rect 10047 20284 10140 20312
rect 4304 20216 4936 20244
rect 4304 20204 4310 20216
rect 6362 20204 6368 20256
rect 6420 20244 6426 20256
rect 7944 20253 7972 20284
rect 7929 20247 7987 20253
rect 7929 20244 7941 20247
rect 6420 20216 7941 20244
rect 6420 20204 6426 20216
rect 7929 20213 7941 20216
rect 7975 20213 7987 20247
rect 7929 20207 7987 20213
rect 8478 20204 8484 20256
rect 8536 20244 8542 20256
rect 8573 20247 8631 20253
rect 8573 20244 8585 20247
rect 8536 20216 8585 20244
rect 8536 20204 8542 20216
rect 8573 20213 8585 20216
rect 8619 20213 8631 20247
rect 8573 20207 8631 20213
rect 9674 20204 9680 20256
rect 9732 20244 9738 20256
rect 10060 20253 10088 20284
rect 10134 20272 10140 20284
rect 10192 20312 10198 20324
rect 10550 20315 10608 20321
rect 10550 20312 10562 20315
rect 10192 20284 10562 20312
rect 10192 20272 10198 20284
rect 10550 20281 10562 20284
rect 10596 20312 10608 20315
rect 11330 20312 11336 20324
rect 10596 20284 11336 20312
rect 10596 20281 10608 20284
rect 10550 20275 10608 20281
rect 11330 20272 11336 20284
rect 11388 20312 11394 20324
rect 11425 20315 11483 20321
rect 11425 20312 11437 20315
rect 11388 20284 11437 20312
rect 11388 20272 11394 20284
rect 11425 20281 11437 20284
rect 11471 20312 11483 20315
rect 12161 20315 12219 20321
rect 12161 20312 12173 20315
rect 11471 20284 12173 20312
rect 11471 20281 11483 20284
rect 11425 20275 11483 20281
rect 12161 20281 12173 20284
rect 12207 20312 12219 20315
rect 12713 20315 12771 20321
rect 12713 20312 12725 20315
rect 12207 20284 12725 20312
rect 12207 20281 12219 20284
rect 12161 20275 12219 20281
rect 12713 20281 12725 20284
rect 12759 20312 12771 20315
rect 13170 20312 13176 20324
rect 12759 20284 13176 20312
rect 12759 20281 12771 20284
rect 12713 20275 12771 20281
rect 13170 20272 13176 20284
rect 13228 20321 13234 20324
rect 13228 20315 13276 20321
rect 13228 20281 13230 20315
rect 13264 20281 13276 20315
rect 13228 20275 13276 20281
rect 13228 20272 13234 20275
rect 15378 20272 15384 20324
rect 15436 20312 15442 20324
rect 15565 20315 15623 20321
rect 15565 20312 15577 20315
rect 15436 20284 15577 20312
rect 15436 20272 15442 20284
rect 15565 20281 15577 20284
rect 15611 20312 15623 20315
rect 15933 20315 15991 20321
rect 15933 20312 15945 20315
rect 15611 20284 15945 20312
rect 15611 20281 15623 20284
rect 15565 20275 15623 20281
rect 15933 20281 15945 20284
rect 15979 20312 15991 20315
rect 16390 20312 16396 20324
rect 15979 20284 16396 20312
rect 15979 20281 15991 20284
rect 15933 20275 15991 20281
rect 16390 20272 16396 20284
rect 16448 20321 16454 20324
rect 16448 20315 16496 20321
rect 16448 20281 16450 20315
rect 16484 20281 16496 20315
rect 18138 20312 18144 20324
rect 18099 20284 18144 20312
rect 16448 20275 16496 20281
rect 16448 20272 16454 20275
rect 18138 20272 18144 20284
rect 18196 20272 18202 20324
rect 18233 20315 18291 20321
rect 18233 20281 18245 20315
rect 18279 20281 18291 20315
rect 18233 20275 18291 20281
rect 10045 20247 10103 20253
rect 10045 20244 10057 20247
rect 9732 20216 10057 20244
rect 9732 20204 9738 20216
rect 10045 20213 10057 20216
rect 10091 20213 10103 20247
rect 10045 20207 10103 20213
rect 14783 20247 14841 20253
rect 14783 20213 14795 20247
rect 14829 20244 14841 20247
rect 15470 20244 15476 20256
rect 14829 20216 15476 20244
rect 14829 20213 14841 20216
rect 14783 20207 14841 20213
rect 15470 20204 15476 20216
rect 15528 20204 15534 20256
rect 17037 20247 17095 20253
rect 17037 20213 17049 20247
rect 17083 20244 17095 20247
rect 17770 20244 17776 20256
rect 17083 20216 17776 20244
rect 17083 20213 17095 20216
rect 17037 20207 17095 20213
rect 17770 20204 17776 20216
rect 17828 20244 17834 20256
rect 18248 20244 18276 20275
rect 18322 20272 18328 20324
rect 18380 20312 18386 20324
rect 19334 20312 19340 20324
rect 18380 20284 19340 20312
rect 18380 20272 18386 20284
rect 19334 20272 19340 20284
rect 19392 20312 19398 20324
rect 19429 20315 19487 20321
rect 19429 20312 19441 20315
rect 19392 20284 19441 20312
rect 19392 20272 19398 20284
rect 19429 20281 19441 20284
rect 19475 20312 19487 20315
rect 19797 20315 19855 20321
rect 19797 20312 19809 20315
rect 19475 20284 19809 20312
rect 19475 20281 19487 20284
rect 19429 20275 19487 20281
rect 19797 20281 19809 20284
rect 19843 20281 19855 20315
rect 20346 20312 20352 20324
rect 20307 20284 20352 20312
rect 19797 20275 19855 20281
rect 20346 20272 20352 20284
rect 20404 20272 20410 20324
rect 18966 20244 18972 20256
rect 17828 20216 18972 20244
rect 17828 20204 17834 20216
rect 18966 20204 18972 20216
rect 19024 20244 19030 20256
rect 19061 20247 19119 20253
rect 19061 20244 19073 20247
rect 19024 20216 19073 20244
rect 19024 20204 19030 20216
rect 19061 20213 19073 20216
rect 19107 20213 19119 20247
rect 19061 20207 19119 20213
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 24719 20247 24777 20253
rect 24719 20244 24731 20247
rect 19576 20216 24731 20244
rect 19576 20204 19582 20216
rect 24719 20213 24731 20216
rect 24765 20213 24777 20247
rect 24719 20207 24777 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 3786 20040 3792 20052
rect 3747 20012 3792 20040
rect 3786 20000 3792 20012
rect 3844 20000 3850 20052
rect 5994 20000 6000 20052
rect 6052 20040 6058 20052
rect 6089 20043 6147 20049
rect 6089 20040 6101 20043
rect 6052 20012 6101 20040
rect 6052 20000 6058 20012
rect 6089 20009 6101 20012
rect 6135 20040 6147 20043
rect 6825 20043 6883 20049
rect 6825 20040 6837 20043
rect 6135 20012 6837 20040
rect 6135 20009 6147 20012
rect 6089 20003 6147 20009
rect 6825 20009 6837 20012
rect 6871 20009 6883 20043
rect 6825 20003 6883 20009
rect 7745 20043 7803 20049
rect 7745 20009 7757 20043
rect 7791 20040 7803 20043
rect 8018 20040 8024 20052
rect 7791 20012 8024 20040
rect 7791 20009 7803 20012
rect 7745 20003 7803 20009
rect 8018 20000 8024 20012
rect 8076 20000 8082 20052
rect 10686 20040 10692 20052
rect 10647 20012 10692 20040
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 13354 20000 13360 20052
rect 13412 20040 13418 20052
rect 13633 20043 13691 20049
rect 13633 20040 13645 20043
rect 13412 20012 13645 20040
rect 13412 20000 13418 20012
rect 13633 20009 13645 20012
rect 13679 20009 13691 20043
rect 13633 20003 13691 20009
rect 14001 20043 14059 20049
rect 14001 20009 14013 20043
rect 14047 20040 14059 20043
rect 14182 20040 14188 20052
rect 14047 20012 14188 20040
rect 14047 20009 14059 20012
rect 14001 20003 14059 20009
rect 14182 20000 14188 20012
rect 14240 20040 14246 20052
rect 14826 20040 14832 20052
rect 14240 20012 14832 20040
rect 14240 20000 14246 20012
rect 14826 20000 14832 20012
rect 14884 20000 14890 20052
rect 16390 20040 16396 20052
rect 16351 20012 16396 20040
rect 16390 20000 16396 20012
rect 16448 20000 16454 20052
rect 16942 20040 16948 20052
rect 16903 20012 16948 20040
rect 16942 20000 16948 20012
rect 17000 20000 17006 20052
rect 18138 20000 18144 20052
rect 18196 20040 18202 20052
rect 19843 20043 19901 20049
rect 19843 20040 19855 20043
rect 18196 20012 19855 20040
rect 18196 20000 18202 20012
rect 19843 20009 19855 20012
rect 19889 20009 19901 20043
rect 19843 20003 19901 20009
rect 3142 19972 3148 19984
rect 3103 19944 3148 19972
rect 3142 19932 3148 19944
rect 3200 19932 3206 19984
rect 4062 19932 4068 19984
rect 4120 19972 4126 19984
rect 4341 19975 4399 19981
rect 4341 19972 4353 19975
rect 4120 19944 4353 19972
rect 4120 19932 4126 19944
rect 4341 19941 4353 19944
rect 4387 19941 4399 19975
rect 4341 19935 4399 19941
rect 4893 19975 4951 19981
rect 4893 19941 4905 19975
rect 4939 19972 4951 19975
rect 4982 19972 4988 19984
rect 4939 19944 4988 19972
rect 4939 19941 4951 19944
rect 4893 19935 4951 19941
rect 4982 19932 4988 19944
rect 5040 19932 5046 19984
rect 6730 19932 6736 19984
rect 6788 19972 6794 19984
rect 7193 19975 7251 19981
rect 7193 19972 7205 19975
rect 6788 19944 7205 19972
rect 6788 19932 6794 19944
rect 7193 19941 7205 19944
rect 7239 19941 7251 19975
rect 7193 19935 7251 19941
rect 8199 19975 8257 19981
rect 8199 19941 8211 19975
rect 8245 19972 8257 19975
rect 9674 19972 9680 19984
rect 8245 19944 9680 19972
rect 8245 19941 8257 19944
rect 8199 19935 8257 19941
rect 2958 19904 2964 19916
rect 2919 19876 2964 19904
rect 2958 19864 2964 19876
rect 3016 19864 3022 19916
rect 6089 19907 6147 19913
rect 6089 19873 6101 19907
rect 6135 19904 6147 19907
rect 6178 19904 6184 19916
rect 6135 19876 6184 19904
rect 6135 19873 6147 19876
rect 6089 19867 6147 19873
rect 6178 19864 6184 19876
rect 6236 19864 6242 19916
rect 6362 19904 6368 19916
rect 6323 19876 6368 19904
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 7742 19864 7748 19916
rect 7800 19904 7806 19916
rect 8214 19904 8242 19935
rect 9674 19932 9680 19944
rect 9732 19932 9738 19984
rect 11054 19932 11060 19984
rect 11112 19972 11118 19984
rect 11149 19975 11207 19981
rect 11149 19972 11161 19975
rect 11112 19944 11161 19972
rect 11112 19932 11118 19944
rect 11149 19941 11161 19944
rect 11195 19972 11207 19975
rect 12158 19972 12164 19984
rect 11195 19944 12164 19972
rect 11195 19941 11207 19944
rect 11149 19935 11207 19941
rect 12158 19932 12164 19944
rect 12216 19932 12222 19984
rect 13075 19975 13133 19981
rect 13075 19941 13087 19975
rect 13121 19972 13133 19975
rect 13170 19972 13176 19984
rect 13121 19944 13176 19972
rect 13121 19941 13133 19944
rect 13075 19935 13133 19941
rect 13170 19932 13176 19944
rect 13228 19972 13234 19984
rect 13906 19972 13912 19984
rect 13228 19944 13912 19972
rect 13228 19932 13234 19944
rect 13906 19932 13912 19944
rect 13964 19932 13970 19984
rect 18322 19972 18328 19984
rect 18283 19944 18328 19972
rect 18322 19932 18328 19944
rect 18380 19932 18386 19984
rect 18874 19972 18880 19984
rect 18835 19944 18880 19972
rect 18874 19932 18880 19944
rect 18932 19932 18938 19984
rect 19242 19972 19248 19984
rect 19203 19944 19248 19972
rect 19242 19932 19248 19944
rect 19300 19932 19306 19984
rect 7800 19876 8242 19904
rect 7800 19864 7806 19876
rect 9398 19864 9404 19916
rect 9456 19904 9462 19916
rect 9804 19907 9862 19913
rect 9804 19904 9816 19907
rect 9456 19876 9816 19904
rect 9456 19864 9462 19876
rect 9804 19873 9816 19876
rect 9850 19873 9862 19907
rect 12710 19904 12716 19916
rect 12671 19876 12716 19904
rect 9804 19867 9862 19873
rect 12710 19864 12716 19876
rect 12768 19864 12774 19916
rect 16025 19907 16083 19913
rect 16025 19873 16037 19907
rect 16071 19904 16083 19907
rect 16114 19904 16120 19916
rect 16071 19876 16120 19904
rect 16071 19873 16083 19876
rect 16025 19867 16083 19873
rect 16114 19864 16120 19876
rect 16172 19904 16178 19916
rect 16482 19904 16488 19916
rect 16172 19876 16488 19904
rect 16172 19864 16178 19876
rect 16482 19864 16488 19876
rect 16540 19864 16546 19916
rect 19702 19904 19708 19916
rect 19663 19876 19708 19904
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 3878 19796 3884 19848
rect 3936 19836 3942 19848
rect 4249 19839 4307 19845
rect 4249 19836 4261 19839
rect 3936 19808 4261 19836
rect 3936 19796 3942 19808
rect 4249 19805 4261 19808
rect 4295 19836 4307 19839
rect 4430 19836 4436 19848
rect 4295 19808 4436 19836
rect 4295 19805 4307 19808
rect 4249 19799 4307 19805
rect 4430 19796 4436 19808
rect 4488 19796 4494 19848
rect 7374 19796 7380 19848
rect 7432 19836 7438 19848
rect 7837 19839 7895 19845
rect 7837 19836 7849 19839
rect 7432 19808 7849 19836
rect 7432 19796 7438 19808
rect 7837 19805 7849 19808
rect 7883 19805 7895 19839
rect 7837 19799 7895 19805
rect 9907 19839 9965 19845
rect 9907 19805 9919 19839
rect 9953 19836 9965 19839
rect 11057 19839 11115 19845
rect 11057 19836 11069 19839
rect 9953 19808 11069 19836
rect 9953 19805 9965 19808
rect 9907 19799 9965 19805
rect 11057 19805 11069 19808
rect 11103 19836 11115 19839
rect 11330 19836 11336 19848
rect 11103 19808 11336 19836
rect 11103 19805 11115 19808
rect 11057 19799 11115 19805
rect 11330 19796 11336 19808
rect 11388 19796 11394 19848
rect 11514 19836 11520 19848
rect 11475 19808 11520 19836
rect 11514 19796 11520 19808
rect 11572 19796 11578 19848
rect 17862 19796 17868 19848
rect 17920 19836 17926 19848
rect 18233 19839 18291 19845
rect 18233 19836 18245 19839
rect 17920 19808 18245 19836
rect 17920 19796 17926 19808
rect 18233 19805 18245 19808
rect 18279 19836 18291 19839
rect 20901 19839 20959 19845
rect 20901 19836 20913 19839
rect 18279 19808 20913 19836
rect 18279 19805 18291 19808
rect 18233 19799 18291 19805
rect 20901 19805 20913 19808
rect 20947 19805 20959 19839
rect 20901 19799 20959 19805
rect 14 19660 20 19712
rect 72 19700 78 19712
rect 4982 19700 4988 19712
rect 72 19672 4988 19700
rect 72 19660 78 19672
rect 4982 19660 4988 19672
rect 5040 19660 5046 19712
rect 8754 19700 8760 19712
rect 8715 19672 8760 19700
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 9950 19660 9956 19712
rect 10008 19700 10014 19712
rect 10229 19703 10287 19709
rect 10229 19700 10241 19703
rect 10008 19672 10241 19700
rect 10008 19660 10014 19672
rect 10229 19669 10241 19672
rect 10275 19669 10287 19703
rect 10229 19663 10287 19669
rect 19426 19660 19432 19712
rect 19484 19700 19490 19712
rect 20165 19703 20223 19709
rect 20165 19700 20177 19703
rect 19484 19672 20177 19700
rect 19484 19660 19490 19672
rect 20165 19669 20177 19672
rect 20211 19669 20223 19703
rect 20165 19663 20223 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 6178 19496 6184 19508
rect 6139 19468 6184 19496
rect 6178 19456 6184 19468
rect 6236 19456 6242 19508
rect 11054 19496 11060 19508
rect 6288 19468 10594 19496
rect 11015 19468 11060 19496
rect 6288 19428 6316 19468
rect 5644 19400 6316 19428
rect 4249 19363 4307 19369
rect 4249 19329 4261 19363
rect 4295 19360 4307 19363
rect 4338 19360 4344 19372
rect 4295 19332 4344 19360
rect 4295 19329 4307 19332
rect 4249 19323 4307 19329
rect 4338 19320 4344 19332
rect 4396 19320 4402 19372
rect 5077 19295 5135 19301
rect 5077 19261 5089 19295
rect 5123 19292 5135 19295
rect 5445 19295 5503 19301
rect 5445 19292 5457 19295
rect 5123 19264 5457 19292
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 5445 19261 5457 19264
rect 5491 19292 5503 19295
rect 5644 19292 5672 19400
rect 7466 19388 7472 19440
rect 7524 19428 7530 19440
rect 8202 19428 8208 19440
rect 7524 19400 8208 19428
rect 7524 19388 7530 19400
rect 8202 19388 8208 19400
rect 8260 19388 8266 19440
rect 10566 19428 10594 19468
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 11330 19496 11336 19508
rect 11291 19468 11336 19496
rect 11330 19456 11336 19468
rect 11388 19456 11394 19508
rect 14090 19496 14096 19508
rect 14003 19468 14096 19496
rect 14090 19456 14096 19468
rect 14148 19496 14154 19508
rect 17586 19496 17592 19508
rect 14148 19468 17592 19496
rect 14148 19456 14154 19468
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 17862 19496 17868 19508
rect 17823 19468 17868 19496
rect 17862 19456 17868 19468
rect 17920 19456 17926 19508
rect 19334 19496 19340 19508
rect 19295 19468 19340 19496
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 19426 19456 19432 19508
rect 19484 19496 19490 19508
rect 19484 19468 19702 19496
rect 19484 19456 19490 19468
rect 11146 19428 11152 19440
rect 10566 19400 11152 19428
rect 11146 19388 11152 19400
rect 11204 19388 11210 19440
rect 16485 19431 16543 19437
rect 16485 19397 16497 19431
rect 16531 19428 16543 19431
rect 16531 19400 19610 19428
rect 16531 19397 16543 19400
rect 16485 19391 16543 19397
rect 5905 19363 5963 19369
rect 5905 19329 5917 19363
rect 5951 19360 5963 19363
rect 7374 19360 7380 19372
rect 5951 19332 7380 19360
rect 5951 19329 5963 19332
rect 5905 19323 5963 19329
rect 7374 19320 7380 19332
rect 7432 19320 7438 19372
rect 7561 19363 7619 19369
rect 7561 19329 7573 19363
rect 7607 19360 7619 19363
rect 7650 19360 7656 19372
rect 7607 19332 7656 19360
rect 7607 19329 7619 19332
rect 7561 19323 7619 19329
rect 7650 19320 7656 19332
rect 7708 19360 7714 19372
rect 8481 19363 8539 19369
rect 8481 19360 8493 19363
rect 7708 19332 8493 19360
rect 7708 19320 7714 19332
rect 8481 19329 8493 19332
rect 8527 19360 8539 19363
rect 8662 19360 8668 19372
rect 8527 19332 8668 19360
rect 8527 19329 8539 19332
rect 8481 19323 8539 19329
rect 8662 19320 8668 19332
rect 8720 19320 8726 19372
rect 8846 19320 8852 19372
rect 8904 19360 8910 19372
rect 9493 19363 9551 19369
rect 9493 19360 9505 19363
rect 8904 19332 9505 19360
rect 8904 19320 8910 19332
rect 9493 19329 9505 19332
rect 9539 19360 9551 19363
rect 13541 19363 13599 19369
rect 13541 19360 13553 19363
rect 9539 19332 13553 19360
rect 9539 19329 9551 19332
rect 9493 19323 9551 19329
rect 5491 19264 5672 19292
rect 5721 19295 5779 19301
rect 5491 19261 5503 19264
rect 5445 19255 5503 19261
rect 5721 19261 5733 19295
rect 5767 19292 5779 19295
rect 6362 19292 6368 19304
rect 5767 19264 6368 19292
rect 5767 19261 5779 19264
rect 5721 19255 5779 19261
rect 6362 19252 6368 19264
rect 6420 19292 6426 19304
rect 10244 19301 10272 19332
rect 13541 19329 13553 19332
rect 13587 19329 13599 19363
rect 13541 19323 13599 19329
rect 13906 19320 13912 19372
rect 13964 19360 13970 19372
rect 15378 19360 15384 19372
rect 13964 19332 15384 19360
rect 13964 19320 13970 19332
rect 15378 19320 15384 19332
rect 15436 19320 15442 19372
rect 18782 19360 18788 19372
rect 18743 19332 18788 19360
rect 18782 19320 18788 19332
rect 18840 19320 18846 19372
rect 19582 19334 19610 19400
rect 10229 19295 10287 19301
rect 6420 19264 6684 19292
rect 6420 19252 6426 19264
rect 3053 19227 3111 19233
rect 3053 19193 3065 19227
rect 3099 19224 3111 19227
rect 3234 19224 3240 19236
rect 3099 19196 3240 19224
rect 3099 19193 3111 19196
rect 3053 19187 3111 19193
rect 3234 19184 3240 19196
rect 3292 19224 3298 19236
rect 3605 19227 3663 19233
rect 3605 19224 3617 19227
rect 3292 19196 3617 19224
rect 3292 19184 3298 19196
rect 3605 19193 3617 19196
rect 3651 19193 3663 19227
rect 3605 19187 3663 19193
rect 3697 19227 3755 19233
rect 3697 19193 3709 19227
rect 3743 19224 3755 19227
rect 3743 19196 4154 19224
rect 3743 19193 3755 19196
rect 3697 19187 3755 19193
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2958 19156 2964 19168
rect 2547 19128 2964 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2958 19116 2964 19128
rect 3016 19156 3022 19168
rect 3421 19159 3479 19165
rect 3421 19156 3433 19159
rect 3016 19128 3433 19156
rect 3016 19116 3022 19128
rect 3421 19125 3433 19128
rect 3467 19156 3479 19159
rect 3712 19156 3740 19187
rect 3467 19128 3740 19156
rect 4126 19156 4154 19196
rect 4338 19156 4344 19168
rect 4126 19128 4344 19156
rect 3467 19125 3479 19128
rect 3421 19119 3479 19125
rect 4338 19116 4344 19128
rect 4396 19116 4402 19168
rect 4522 19156 4528 19168
rect 4483 19128 4528 19156
rect 4522 19116 4528 19128
rect 4580 19116 4586 19168
rect 6656 19165 6684 19264
rect 10229 19261 10241 19295
rect 10275 19261 10287 19295
rect 10229 19255 10287 19261
rect 10413 19295 10471 19301
rect 10413 19261 10425 19295
rect 10459 19261 10471 19295
rect 10413 19255 10471 19261
rect 6914 19224 6920 19236
rect 6875 19196 6920 19224
rect 6914 19184 6920 19196
rect 6972 19184 6978 19236
rect 7006 19184 7012 19236
rect 7064 19224 7070 19236
rect 8573 19227 8631 19233
rect 7064 19196 7109 19224
rect 7064 19184 7070 19196
rect 8573 19193 8585 19227
rect 8619 19224 8631 19227
rect 8754 19224 8760 19236
rect 8619 19196 8760 19224
rect 8619 19193 8631 19196
rect 8573 19187 8631 19193
rect 6641 19159 6699 19165
rect 6641 19125 6653 19159
rect 6687 19156 6699 19159
rect 6730 19156 6736 19168
rect 6687 19128 6736 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 6730 19116 6736 19128
rect 6788 19116 6794 19168
rect 7742 19116 7748 19168
rect 7800 19156 7806 19168
rect 7837 19159 7895 19165
rect 7837 19156 7849 19159
rect 7800 19128 7849 19156
rect 7800 19116 7806 19128
rect 7837 19125 7849 19128
rect 7883 19125 7895 19159
rect 7837 19119 7895 19125
rect 8297 19159 8355 19165
rect 8297 19125 8309 19159
rect 8343 19156 8355 19159
rect 8588 19156 8616 19187
rect 8754 19184 8760 19196
rect 8812 19184 8818 19236
rect 9125 19227 9183 19233
rect 9125 19193 9137 19227
rect 9171 19224 9183 19227
rect 9582 19224 9588 19236
rect 9171 19196 9588 19224
rect 9171 19193 9183 19196
rect 9125 19187 9183 19193
rect 9582 19184 9588 19196
rect 9640 19184 9646 19236
rect 9950 19184 9956 19236
rect 10008 19224 10014 19236
rect 10428 19224 10456 19255
rect 11054 19252 11060 19304
rect 11112 19292 11118 19304
rect 12897 19295 12955 19301
rect 12897 19292 12909 19295
rect 11112 19264 12909 19292
rect 11112 19252 11118 19264
rect 12897 19261 12909 19264
rect 12943 19292 12955 19295
rect 13357 19295 13415 19301
rect 13357 19292 13369 19295
rect 12943 19264 13369 19292
rect 12943 19261 12955 19264
rect 12897 19255 12955 19261
rect 13357 19261 13369 19264
rect 13403 19261 13415 19295
rect 14182 19292 14188 19304
rect 13357 19255 13415 19261
rect 13786 19264 14188 19292
rect 13786 19236 13814 19264
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 14461 19295 14519 19301
rect 14461 19261 14473 19295
rect 14507 19261 14519 19295
rect 14461 19255 14519 19261
rect 13786 19224 13820 19236
rect 10008 19196 10456 19224
rect 13233 19196 13820 19224
rect 10008 19184 10014 19196
rect 8343 19128 8616 19156
rect 8343 19125 8355 19128
rect 8297 19119 8355 19125
rect 9398 19116 9404 19168
rect 9456 19156 9462 19168
rect 9769 19159 9827 19165
rect 9769 19156 9781 19159
rect 9456 19128 9781 19156
rect 9456 19116 9462 19128
rect 9769 19125 9781 19128
rect 9815 19125 9827 19159
rect 10042 19156 10048 19168
rect 10003 19128 10048 19156
rect 9769 19119 9827 19125
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 12802 19156 12808 19168
rect 12763 19128 12808 19156
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 13081 19159 13139 19165
rect 13081 19125 13093 19159
rect 13127 19156 13139 19159
rect 13233 19156 13261 19196
rect 13814 19184 13820 19196
rect 13872 19184 13878 19236
rect 13127 19128 13261 19156
rect 13541 19159 13599 19165
rect 13127 19125 13139 19128
rect 13081 19119 13139 19125
rect 13541 19125 13553 19159
rect 13587 19156 13599 19159
rect 13725 19159 13783 19165
rect 13725 19156 13737 19159
rect 13587 19128 13737 19156
rect 13587 19125 13599 19128
rect 13541 19119 13599 19125
rect 13725 19125 13737 19128
rect 13771 19156 13783 19159
rect 14366 19156 14372 19168
rect 13771 19128 14372 19156
rect 13771 19125 13783 19128
rect 13725 19119 13783 19125
rect 14366 19116 14372 19128
rect 14424 19156 14430 19168
rect 14476 19156 14504 19255
rect 14642 19224 14648 19236
rect 14603 19196 14648 19224
rect 14642 19184 14648 19196
rect 14700 19184 14706 19236
rect 15396 19224 15424 19320
rect 19536 19306 19610 19334
rect 19674 19360 19702 19468
rect 19889 19363 19947 19369
rect 19889 19360 19901 19363
rect 19674 19332 19901 19360
rect 19889 19329 19901 19332
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 20070 19320 20076 19372
rect 20128 19360 20134 19372
rect 20165 19363 20223 19369
rect 20165 19360 20177 19363
rect 20128 19332 20177 19360
rect 20128 19320 20134 19332
rect 20165 19329 20177 19332
rect 20211 19329 20223 19363
rect 20165 19323 20223 19329
rect 15562 19292 15568 19304
rect 15523 19264 15568 19292
rect 15562 19252 15568 19264
rect 15620 19252 15626 19304
rect 15886 19227 15944 19233
rect 15886 19224 15898 19227
rect 15396 19196 15898 19224
rect 15886 19193 15898 19196
rect 15932 19224 15944 19227
rect 15932 19196 16252 19224
rect 15932 19193 15944 19196
rect 15886 19187 15944 19193
rect 14424 19128 14504 19156
rect 16224 19156 16252 19196
rect 16298 19184 16304 19236
rect 16356 19224 16362 19236
rect 17405 19227 17463 19233
rect 17405 19224 17417 19227
rect 16356 19196 17417 19224
rect 16356 19184 16362 19196
rect 17405 19193 17417 19196
rect 17451 19193 17463 19227
rect 18322 19224 18328 19236
rect 18283 19196 18328 19224
rect 17405 19187 17463 19193
rect 16574 19156 16580 19168
rect 16224 19128 16580 19156
rect 14424 19116 14430 19128
rect 16574 19116 16580 19128
rect 16632 19156 16638 19168
rect 16761 19159 16819 19165
rect 16761 19156 16773 19159
rect 16632 19128 16773 19156
rect 16632 19116 16638 19128
rect 16761 19125 16773 19128
rect 16807 19125 16819 19159
rect 17420 19156 17448 19187
rect 18322 19184 18328 19196
rect 18380 19184 18386 19236
rect 18417 19227 18475 19233
rect 18417 19193 18429 19227
rect 18463 19193 18475 19227
rect 19536 19224 19564 19306
rect 19702 19292 19708 19304
rect 19663 19264 19708 19292
rect 19702 19252 19708 19264
rect 19760 19252 19766 19304
rect 19981 19227 20039 19233
rect 19981 19224 19993 19227
rect 19536 19196 19993 19224
rect 18417 19187 18475 19193
rect 19981 19193 19993 19196
rect 20027 19224 20039 19227
rect 20070 19224 20076 19236
rect 20027 19196 20076 19224
rect 20027 19193 20039 19196
rect 19981 19187 20039 19193
rect 18432 19156 18460 19187
rect 20070 19184 20076 19196
rect 20128 19184 20134 19236
rect 19518 19156 19524 19168
rect 17420 19128 19524 19156
rect 16761 19119 16819 19125
rect 19518 19116 19524 19128
rect 19576 19116 19582 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 3878 18952 3884 18964
rect 3839 18924 3884 18952
rect 3878 18912 3884 18924
rect 3936 18912 3942 18964
rect 7374 18912 7380 18964
rect 7432 18952 7438 18964
rect 8389 18955 8447 18961
rect 8389 18952 8401 18955
rect 7432 18924 8401 18952
rect 7432 18912 7438 18924
rect 8389 18921 8401 18924
rect 8435 18921 8447 18955
rect 8389 18915 8447 18921
rect 8662 18912 8668 18964
rect 8720 18952 8726 18964
rect 8757 18955 8815 18961
rect 8757 18952 8769 18955
rect 8720 18924 8769 18952
rect 8720 18912 8726 18924
rect 8757 18921 8769 18924
rect 8803 18921 8815 18955
rect 12710 18952 12716 18964
rect 12671 18924 12716 18952
rect 8757 18915 8815 18921
rect 12710 18912 12716 18924
rect 12768 18912 12774 18964
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 13906 18952 13912 18964
rect 12860 18924 13912 18952
rect 12860 18912 12866 18924
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 14642 18912 14648 18964
rect 14700 18952 14706 18964
rect 14737 18955 14795 18961
rect 14737 18952 14749 18955
rect 14700 18924 14749 18952
rect 14700 18912 14706 18924
rect 14737 18921 14749 18924
rect 14783 18921 14795 18955
rect 16114 18952 16120 18964
rect 16075 18924 16120 18952
rect 14737 18915 14795 18921
rect 16114 18912 16120 18924
rect 16172 18912 16178 18964
rect 16574 18952 16580 18964
rect 16535 18924 16580 18952
rect 16574 18912 16580 18924
rect 16632 18912 16638 18964
rect 17129 18955 17187 18961
rect 17129 18921 17141 18955
rect 17175 18952 17187 18955
rect 18230 18952 18236 18964
rect 17175 18924 18236 18952
rect 17175 18921 17187 18924
rect 17129 18915 17187 18921
rect 18230 18912 18236 18924
rect 18288 18912 18294 18964
rect 18322 18912 18328 18964
rect 18380 18952 18386 18964
rect 18969 18955 19027 18961
rect 18969 18952 18981 18955
rect 18380 18924 18981 18952
rect 18380 18912 18386 18924
rect 18969 18921 18981 18924
rect 19015 18952 19027 18955
rect 19659 18955 19717 18961
rect 19659 18952 19671 18955
rect 19015 18924 19671 18952
rect 19015 18921 19027 18924
rect 18969 18915 19027 18921
rect 19659 18921 19671 18924
rect 19705 18921 19717 18955
rect 20070 18952 20076 18964
rect 20031 18924 20076 18952
rect 19659 18915 19717 18921
rect 20070 18912 20076 18924
rect 20128 18912 20134 18964
rect 3234 18884 3240 18896
rect 3195 18856 3240 18884
rect 3234 18844 3240 18856
rect 3292 18844 3298 18896
rect 4062 18884 4068 18896
rect 3975 18856 4068 18884
rect 4062 18844 4068 18856
rect 4120 18884 4126 18896
rect 4522 18884 4528 18896
rect 4120 18856 4528 18884
rect 4120 18844 4126 18856
rect 4522 18844 4528 18856
rect 4580 18844 4586 18896
rect 5997 18887 6055 18893
rect 5997 18853 6009 18887
rect 6043 18884 6055 18887
rect 6917 18887 6975 18893
rect 6917 18884 6929 18887
rect 6043 18856 6929 18884
rect 6043 18853 6055 18856
rect 5997 18847 6055 18853
rect 6917 18853 6929 18856
rect 6963 18884 6975 18887
rect 7006 18884 7012 18896
rect 6963 18856 7012 18884
rect 6963 18853 6975 18856
rect 6917 18847 6975 18853
rect 7006 18844 7012 18856
rect 7064 18884 7070 18896
rect 7558 18884 7564 18896
rect 7064 18856 7564 18884
rect 7064 18844 7070 18856
rect 7558 18844 7564 18856
rect 7616 18844 7622 18896
rect 9861 18887 9919 18893
rect 9861 18853 9873 18887
rect 9907 18884 9919 18887
rect 10134 18884 10140 18896
rect 9907 18856 10140 18884
rect 9907 18853 9919 18856
rect 9861 18847 9919 18853
rect 10134 18844 10140 18856
rect 10192 18844 10198 18896
rect 11701 18887 11759 18893
rect 11701 18853 11713 18887
rect 11747 18884 11759 18887
rect 11790 18884 11796 18896
rect 11747 18856 11796 18884
rect 11747 18853 11759 18856
rect 11701 18847 11759 18853
rect 11790 18844 11796 18856
rect 11848 18844 11854 18896
rect 13078 18844 13084 18896
rect 13136 18884 13142 18896
rect 14369 18887 14427 18893
rect 13136 18856 14136 18884
rect 13136 18844 13142 18856
rect 14108 18828 14136 18856
rect 14369 18853 14381 18887
rect 14415 18884 14427 18887
rect 15562 18884 15568 18896
rect 14415 18856 15568 18884
rect 14415 18853 14427 18856
rect 14369 18847 14427 18853
rect 15562 18844 15568 18856
rect 15620 18844 15626 18896
rect 17862 18844 17868 18896
rect 17920 18884 17926 18896
rect 18141 18887 18199 18893
rect 18141 18884 18153 18887
rect 17920 18856 18153 18884
rect 17920 18844 17926 18856
rect 18141 18853 18153 18856
rect 18187 18853 18199 18887
rect 18141 18847 18199 18853
rect 1302 18776 1308 18828
rect 1360 18816 1366 18828
rect 1432 18819 1490 18825
rect 1432 18816 1444 18819
rect 1360 18788 1444 18816
rect 1360 18776 1366 18788
rect 1432 18785 1444 18788
rect 1478 18785 1490 18819
rect 1432 18779 1490 18785
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18816 2927 18819
rect 3050 18816 3056 18828
rect 2915 18788 3056 18816
rect 2915 18785 2927 18788
rect 2869 18779 2927 18785
rect 3050 18776 3056 18788
rect 3108 18776 3114 18828
rect 3970 18776 3976 18828
rect 4028 18816 4034 18828
rect 4709 18819 4767 18825
rect 4709 18816 4721 18819
rect 4028 18788 4721 18816
rect 4028 18776 4034 18788
rect 4709 18785 4721 18788
rect 4755 18816 4767 18819
rect 4798 18816 4804 18828
rect 4755 18788 4804 18816
rect 4755 18785 4767 18788
rect 4709 18779 4767 18785
rect 4798 18776 4804 18788
rect 4856 18776 4862 18828
rect 6549 18819 6607 18825
rect 6549 18785 6561 18819
rect 6595 18816 6607 18819
rect 7282 18816 7288 18828
rect 6595 18788 7288 18816
rect 6595 18785 6607 18788
rect 6549 18779 6607 18785
rect 7282 18776 7288 18788
rect 7340 18776 7346 18828
rect 13814 18776 13820 18828
rect 13872 18816 13878 18828
rect 14090 18816 14096 18828
rect 13872 18788 13917 18816
rect 14051 18788 14096 18816
rect 13872 18776 13878 18788
rect 14090 18776 14096 18788
rect 14148 18776 14154 18828
rect 19242 18776 19248 18828
rect 19300 18816 19306 18828
rect 19556 18819 19614 18825
rect 19556 18816 19568 18819
rect 19300 18788 19568 18816
rect 19300 18776 19306 18788
rect 19556 18785 19568 18788
rect 19602 18785 19614 18819
rect 19556 18779 19614 18785
rect 5905 18751 5963 18757
rect 5905 18717 5917 18751
rect 5951 18717 5963 18751
rect 5905 18711 5963 18717
rect 4430 18640 4436 18692
rect 4488 18680 4494 18692
rect 5629 18683 5687 18689
rect 5629 18680 5641 18683
rect 4488 18652 5641 18680
rect 4488 18640 4494 18652
rect 5629 18649 5641 18652
rect 5675 18680 5687 18683
rect 5920 18680 5948 18711
rect 6638 18708 6644 18760
rect 6696 18748 6702 18760
rect 7469 18751 7527 18757
rect 7469 18748 7481 18751
rect 6696 18720 7481 18748
rect 6696 18708 6702 18720
rect 7469 18717 7481 18720
rect 7515 18717 7527 18751
rect 7469 18711 7527 18717
rect 7745 18751 7803 18757
rect 7745 18717 7757 18751
rect 7791 18748 7803 18751
rect 9401 18751 9459 18757
rect 9401 18748 9413 18751
rect 7791 18720 9413 18748
rect 7791 18717 7803 18720
rect 7745 18711 7803 18717
rect 9401 18717 9413 18720
rect 9447 18748 9459 18751
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 9447 18720 9781 18748
rect 9447 18717 9459 18720
rect 9401 18711 9459 18717
rect 9769 18717 9781 18720
rect 9815 18717 9827 18751
rect 9769 18711 9827 18717
rect 10045 18751 10103 18757
rect 10045 18717 10057 18751
rect 10091 18717 10103 18751
rect 11609 18751 11667 18757
rect 11609 18748 11621 18751
rect 10045 18711 10103 18717
rect 11348 18720 11621 18748
rect 5675 18652 5948 18680
rect 5675 18649 5687 18652
rect 5629 18643 5687 18649
rect 7190 18640 7196 18692
rect 7248 18680 7254 18692
rect 7760 18680 7788 18711
rect 7248 18652 7788 18680
rect 7248 18640 7254 18652
rect 9582 18640 9588 18692
rect 9640 18680 9646 18692
rect 10060 18680 10088 18711
rect 9640 18652 10088 18680
rect 9640 18640 9646 18652
rect 1535 18615 1593 18621
rect 1535 18581 1547 18615
rect 1581 18612 1593 18615
rect 1670 18612 1676 18624
rect 1581 18584 1676 18612
rect 1581 18581 1593 18584
rect 1535 18575 1593 18581
rect 1670 18572 1676 18584
rect 1728 18572 1734 18624
rect 3510 18612 3516 18624
rect 3471 18584 3516 18612
rect 3510 18572 3516 18584
rect 3568 18572 3574 18624
rect 5258 18612 5264 18624
rect 5219 18584 5264 18612
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 7285 18615 7343 18621
rect 7285 18581 7297 18615
rect 7331 18612 7343 18615
rect 7466 18612 7472 18624
rect 7331 18584 7472 18612
rect 7331 18581 7343 18584
rect 7285 18575 7343 18581
rect 7466 18572 7472 18584
rect 7524 18572 7530 18624
rect 11238 18572 11244 18624
rect 11296 18612 11302 18624
rect 11348 18621 11376 18720
rect 11609 18717 11621 18720
rect 11655 18717 11667 18751
rect 11609 18711 11667 18717
rect 12253 18751 12311 18757
rect 12253 18717 12265 18751
rect 12299 18748 12311 18751
rect 12802 18748 12808 18760
rect 12299 18720 12808 18748
rect 12299 18717 12311 18720
rect 12253 18711 12311 18717
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 16206 18748 16212 18760
rect 16167 18720 16212 18748
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 17865 18751 17923 18757
rect 17865 18717 17877 18751
rect 17911 18748 17923 18751
rect 18046 18748 18052 18760
rect 17911 18720 18052 18748
rect 17911 18717 17923 18720
rect 17865 18711 17923 18717
rect 18046 18708 18052 18720
rect 18104 18708 18110 18760
rect 18414 18748 18420 18760
rect 18375 18720 18420 18748
rect 18414 18708 18420 18720
rect 18472 18748 18478 18760
rect 19426 18748 19432 18760
rect 18472 18720 19432 18748
rect 18472 18708 18478 18720
rect 19426 18708 19432 18720
rect 19484 18708 19490 18760
rect 14458 18640 14464 18692
rect 14516 18680 14522 18692
rect 18506 18680 18512 18692
rect 14516 18652 18512 18680
rect 14516 18640 14522 18652
rect 18506 18640 18512 18652
rect 18564 18680 18570 18692
rect 19334 18680 19340 18692
rect 18564 18652 19340 18680
rect 18564 18640 18570 18652
rect 19334 18640 19340 18652
rect 19392 18640 19398 18692
rect 11333 18615 11391 18621
rect 11333 18612 11345 18615
rect 11296 18584 11345 18612
rect 11296 18572 11302 18584
rect 11333 18581 11345 18584
rect 11379 18581 11391 18615
rect 11333 18575 11391 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 4338 18408 4344 18420
rect 4299 18380 4344 18408
rect 4338 18368 4344 18380
rect 4396 18368 4402 18420
rect 6638 18408 6644 18420
rect 6599 18380 6644 18408
rect 6638 18368 6644 18380
rect 6696 18368 6702 18420
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 8665 18411 8723 18417
rect 8665 18408 8677 18411
rect 7616 18380 8677 18408
rect 7616 18368 7622 18380
rect 8665 18377 8677 18380
rect 8711 18377 8723 18411
rect 8665 18371 8723 18377
rect 14734 18368 14740 18420
rect 14792 18408 14798 18420
rect 17862 18408 17868 18420
rect 14792 18380 16573 18408
rect 17823 18380 17868 18408
rect 14792 18368 14798 18380
rect 2593 18343 2651 18349
rect 2593 18309 2605 18343
rect 2639 18340 2651 18343
rect 5258 18340 5264 18352
rect 2639 18312 5264 18340
rect 2639 18309 2651 18312
rect 2593 18303 2651 18309
rect 5258 18300 5264 18312
rect 5316 18300 5322 18352
rect 6273 18343 6331 18349
rect 6273 18309 6285 18343
rect 6319 18340 6331 18343
rect 6454 18340 6460 18352
rect 6319 18312 6460 18340
rect 6319 18309 6331 18312
rect 6273 18303 6331 18309
rect 6454 18300 6460 18312
rect 6512 18340 6518 18352
rect 7576 18340 7604 18368
rect 6512 18312 7604 18340
rect 6512 18300 6518 18312
rect 9214 18300 9220 18352
rect 9272 18340 9278 18352
rect 11882 18340 11888 18352
rect 9272 18312 11888 18340
rect 9272 18300 9278 18312
rect 11882 18300 11888 18312
rect 11940 18340 11946 18352
rect 13538 18340 13544 18352
rect 11940 18312 13544 18340
rect 11940 18300 11946 18312
rect 13538 18300 13544 18312
rect 13596 18300 13602 18352
rect 13722 18300 13728 18352
rect 13780 18340 13786 18352
rect 14458 18340 14464 18352
rect 13780 18312 14464 18340
rect 13780 18300 13786 18312
rect 14458 18300 14464 18312
rect 14516 18300 14522 18352
rect 15378 18300 15384 18352
rect 15436 18340 15442 18352
rect 16209 18343 16267 18349
rect 16209 18340 16221 18343
rect 15436 18312 16221 18340
rect 15436 18300 15442 18312
rect 16209 18309 16221 18312
rect 16255 18309 16267 18343
rect 16545 18340 16573 18380
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 19242 18340 19248 18352
rect 16545 18312 19248 18340
rect 16209 18303 16267 18309
rect 19242 18300 19248 18312
rect 19300 18340 19306 18352
rect 19429 18343 19487 18349
rect 19429 18340 19441 18343
rect 19300 18312 19441 18340
rect 19300 18300 19306 18312
rect 19429 18309 19441 18312
rect 19475 18309 19487 18343
rect 19429 18303 19487 18309
rect 1302 18232 1308 18284
rect 1360 18272 1366 18284
rect 2225 18275 2283 18281
rect 2225 18272 2237 18275
rect 1360 18244 2237 18272
rect 1360 18232 1366 18244
rect 2225 18241 2237 18244
rect 2271 18241 2283 18275
rect 2225 18235 2283 18241
rect 7282 18232 7288 18284
rect 7340 18272 7346 18284
rect 9306 18272 9312 18284
rect 7340 18244 9312 18272
rect 7340 18232 7346 18244
rect 9306 18232 9312 18244
rect 9364 18232 9370 18284
rect 9582 18272 9588 18284
rect 9543 18244 9588 18272
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18272 12587 18275
rect 12618 18272 12624 18284
rect 12575 18244 12624 18272
rect 12575 18241 12587 18244
rect 12529 18235 12587 18241
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 12802 18272 12808 18284
rect 12763 18244 12808 18272
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 14642 18232 14648 18284
rect 14700 18272 14706 18284
rect 14737 18275 14795 18281
rect 14737 18272 14749 18275
rect 14700 18244 14749 18272
rect 14700 18232 14706 18244
rect 14737 18241 14749 18244
rect 14783 18241 14795 18275
rect 18414 18272 18420 18284
rect 18375 18244 18420 18272
rect 14737 18235 14795 18241
rect 18414 18232 18420 18244
rect 18472 18232 18478 18284
rect 20346 18272 20352 18284
rect 20307 18244 20352 18272
rect 20346 18232 20352 18244
rect 20404 18232 20410 18284
rect 1464 18207 1522 18213
rect 1464 18173 1476 18207
rect 1510 18204 1522 18207
rect 2409 18207 2467 18213
rect 1510 18176 1992 18204
rect 1510 18173 1522 18176
rect 1464 18167 1522 18173
rect 1535 18071 1593 18077
rect 1535 18037 1547 18071
rect 1581 18068 1593 18071
rect 1854 18068 1860 18080
rect 1581 18040 1860 18068
rect 1581 18037 1593 18040
rect 1535 18031 1593 18037
rect 1854 18028 1860 18040
rect 1912 18028 1918 18080
rect 1964 18077 1992 18176
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 2498 18204 2504 18216
rect 2455 18176 2504 18204
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 2498 18164 2504 18176
rect 2556 18164 2562 18216
rect 3421 18207 3479 18213
rect 3421 18173 3433 18207
rect 3467 18204 3479 18207
rect 3510 18204 3516 18216
rect 3467 18176 3516 18204
rect 3467 18173 3479 18176
rect 3421 18167 3479 18173
rect 3510 18164 3516 18176
rect 3568 18204 3574 18216
rect 3878 18204 3884 18216
rect 3568 18176 3884 18204
rect 3568 18164 3574 18176
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 5169 18207 5227 18213
rect 5169 18173 5181 18207
rect 5215 18204 5227 18207
rect 5534 18204 5540 18216
rect 5215 18176 5540 18204
rect 5215 18173 5227 18176
rect 5169 18167 5227 18173
rect 1949 18071 2007 18077
rect 1949 18037 1961 18071
rect 1995 18068 2007 18071
rect 2130 18068 2136 18080
rect 1995 18040 2136 18068
rect 1995 18037 2007 18040
rect 1949 18031 2007 18037
rect 2130 18028 2136 18040
rect 2188 18028 2194 18080
rect 3050 18068 3056 18080
rect 3011 18040 3056 18068
rect 3050 18028 3056 18040
rect 3108 18028 3114 18080
rect 3418 18028 3424 18080
rect 3476 18068 3482 18080
rect 3789 18071 3847 18077
rect 3789 18068 3801 18071
rect 3476 18040 3801 18068
rect 3476 18028 3482 18040
rect 3789 18037 3801 18040
rect 3835 18037 3847 18071
rect 3789 18031 3847 18037
rect 4709 18071 4767 18077
rect 4709 18037 4721 18071
rect 4755 18068 4767 18071
rect 4798 18068 4804 18080
rect 4755 18040 4804 18068
rect 4755 18037 4767 18040
rect 4709 18031 4767 18037
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 5074 18068 5080 18080
rect 5035 18040 5080 18068
rect 5074 18028 5080 18040
rect 5132 18068 5138 18080
rect 5184 18068 5212 18167
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 5721 18207 5779 18213
rect 5721 18173 5733 18207
rect 5767 18173 5779 18207
rect 7466 18204 7472 18216
rect 7427 18176 7472 18204
rect 5721 18167 5779 18173
rect 5258 18096 5264 18148
rect 5316 18136 5322 18148
rect 5736 18136 5764 18167
rect 7466 18164 7472 18176
rect 7524 18164 7530 18216
rect 8389 18207 8447 18213
rect 8389 18173 8401 18207
rect 8435 18204 8447 18207
rect 9033 18207 9091 18213
rect 9033 18204 9045 18207
rect 8435 18176 9045 18204
rect 8435 18173 8447 18176
rect 8389 18167 8447 18173
rect 9033 18173 9045 18176
rect 9079 18173 9091 18207
rect 9033 18167 9091 18173
rect 10689 18207 10747 18213
rect 10689 18173 10701 18207
rect 10735 18204 10747 18207
rect 11422 18204 11428 18216
rect 10735 18176 11428 18204
rect 10735 18173 10747 18176
rect 10689 18167 10747 18173
rect 6730 18136 6736 18148
rect 5316 18108 6736 18136
rect 5316 18096 5322 18108
rect 6730 18096 6736 18108
rect 6788 18136 6794 18148
rect 7374 18136 7380 18148
rect 6788 18108 7380 18136
rect 6788 18096 6794 18108
rect 7374 18096 7380 18108
rect 7432 18096 7438 18148
rect 5132 18040 5212 18068
rect 5445 18071 5503 18077
rect 5132 18028 5138 18040
rect 5445 18037 5457 18071
rect 5491 18068 5503 18071
rect 5534 18068 5540 18080
rect 5491 18040 5540 18068
rect 5491 18037 5503 18040
rect 5445 18031 5503 18037
rect 5534 18028 5540 18040
rect 5592 18028 5598 18080
rect 7285 18071 7343 18077
rect 7285 18037 7297 18071
rect 7331 18068 7343 18071
rect 7742 18068 7748 18080
rect 7331 18040 7748 18068
rect 7331 18037 7343 18040
rect 7285 18031 7343 18037
rect 7742 18028 7748 18040
rect 7800 18068 7806 18080
rect 7837 18071 7895 18077
rect 7837 18068 7849 18071
rect 7800 18040 7849 18068
rect 7800 18028 7806 18040
rect 7837 18037 7849 18040
rect 7883 18037 7895 18071
rect 9048 18068 9076 18167
rect 11422 18164 11428 18176
rect 11480 18164 11486 18216
rect 13725 18207 13783 18213
rect 13725 18173 13737 18207
rect 13771 18204 13783 18207
rect 13814 18204 13820 18216
rect 13771 18176 13820 18204
rect 13771 18173 13783 18176
rect 13725 18167 13783 18173
rect 13814 18164 13820 18176
rect 13872 18164 13878 18216
rect 16206 18164 16212 18216
rect 16264 18204 16270 18216
rect 16945 18207 17003 18213
rect 16945 18204 16957 18207
rect 16264 18176 16957 18204
rect 16264 18164 16270 18176
rect 16945 18173 16957 18176
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 9401 18139 9459 18145
rect 9401 18105 9413 18139
rect 9447 18105 9459 18139
rect 11514 18136 11520 18148
rect 11475 18108 11520 18136
rect 9401 18099 9459 18105
rect 9416 18068 9444 18099
rect 11514 18096 11520 18108
rect 11572 18096 11578 18148
rect 12621 18139 12679 18145
rect 12621 18105 12633 18139
rect 12667 18105 12679 18139
rect 12621 18099 12679 18105
rect 9048 18040 9444 18068
rect 7837 18031 7895 18037
rect 10134 18028 10140 18080
rect 10192 18068 10198 18080
rect 10229 18071 10287 18077
rect 10229 18068 10241 18071
rect 10192 18040 10241 18068
rect 10192 18028 10198 18040
rect 10229 18037 10241 18040
rect 10275 18037 10287 18071
rect 11790 18068 11796 18080
rect 11751 18040 11796 18068
rect 10229 18031 10287 18037
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 12250 18068 12256 18080
rect 12211 18040 12256 18068
rect 12250 18028 12256 18040
rect 12308 18068 12314 18080
rect 12636 18068 12664 18099
rect 15194 18096 15200 18148
rect 15252 18136 15258 18148
rect 16485 18139 16543 18145
rect 16485 18136 16497 18139
rect 15252 18108 16497 18136
rect 15252 18096 15258 18108
rect 16485 18105 16497 18108
rect 16531 18105 16543 18139
rect 16485 18099 16543 18105
rect 17126 18096 17132 18148
rect 17184 18136 17190 18148
rect 18141 18139 18199 18145
rect 18141 18136 18153 18139
rect 17184 18108 18153 18136
rect 17184 18096 17190 18108
rect 18141 18105 18153 18108
rect 18187 18105 18199 18139
rect 18141 18099 18199 18105
rect 18230 18096 18236 18148
rect 18288 18136 18294 18148
rect 19153 18139 19211 18145
rect 18288 18108 18333 18136
rect 18288 18096 18294 18108
rect 19153 18105 19165 18139
rect 19199 18136 19211 18139
rect 19334 18136 19340 18148
rect 19199 18108 19340 18136
rect 19199 18105 19211 18108
rect 19153 18099 19211 18105
rect 19334 18096 19340 18108
rect 19392 18136 19398 18148
rect 19705 18139 19763 18145
rect 19705 18136 19717 18139
rect 19392 18108 19717 18136
rect 19392 18096 19398 18108
rect 19705 18105 19717 18108
rect 19751 18105 19763 18139
rect 19705 18099 19763 18105
rect 19797 18139 19855 18145
rect 19797 18105 19809 18139
rect 19843 18105 19855 18139
rect 19797 18099 19855 18105
rect 14090 18068 14096 18080
rect 12308 18040 12664 18068
rect 14051 18040 14096 18068
rect 12308 18028 12314 18040
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 14645 18071 14703 18077
rect 14645 18037 14657 18071
rect 14691 18068 14703 18071
rect 15105 18071 15163 18077
rect 15105 18068 15117 18071
rect 14691 18040 15117 18068
rect 14691 18037 14703 18040
rect 14645 18031 14703 18037
rect 15105 18037 15117 18040
rect 15151 18068 15163 18071
rect 15378 18068 15384 18080
rect 15151 18040 15384 18068
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 15654 18068 15660 18080
rect 15615 18040 15660 18068
rect 15654 18028 15660 18040
rect 15712 18028 15718 18080
rect 17497 18071 17555 18077
rect 17497 18037 17509 18071
rect 17543 18068 17555 18071
rect 18248 18068 18276 18096
rect 17543 18040 18276 18068
rect 17543 18037 17555 18040
rect 17497 18031 17555 18037
rect 19518 18028 19524 18080
rect 19576 18068 19582 18080
rect 19812 18068 19840 18099
rect 19576 18040 19840 18068
rect 19576 18028 19582 18040
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1670 17864 1676 17876
rect 1631 17836 1676 17864
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 5258 17864 5264 17876
rect 5219 17836 5264 17864
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 6454 17864 6460 17876
rect 6415 17836 6460 17864
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 6914 17864 6920 17876
rect 6875 17836 6920 17864
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 7742 17864 7748 17876
rect 7703 17836 7748 17864
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 8297 17867 8355 17873
rect 8297 17833 8309 17867
rect 8343 17864 8355 17867
rect 10134 17864 10140 17876
rect 8343 17836 10140 17864
rect 8343 17833 8355 17836
rect 8297 17827 8355 17833
rect 10134 17824 10140 17836
rect 10192 17824 10198 17876
rect 13906 17864 13912 17876
rect 10244 17836 13912 17864
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 5899 17799 5957 17805
rect 1820 17768 4154 17796
rect 1820 17756 1826 17768
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 2406 17728 2412 17740
rect 1995 17700 2412 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 2406 17688 2412 17700
rect 2464 17688 2470 17740
rect 2961 17731 3019 17737
rect 2961 17697 2973 17731
rect 3007 17728 3019 17731
rect 3326 17728 3332 17740
rect 3007 17700 3332 17728
rect 3007 17697 3019 17700
rect 2961 17691 3019 17697
rect 3326 17688 3332 17700
rect 3384 17688 3390 17740
rect 4126 17728 4154 17768
rect 5899 17765 5911 17799
rect 5945 17796 5957 17799
rect 5994 17796 6000 17808
rect 5945 17768 6000 17796
rect 5945 17765 5957 17768
rect 5899 17759 5957 17765
rect 5994 17756 6000 17768
rect 6052 17796 6058 17808
rect 7760 17796 7788 17824
rect 9306 17796 9312 17808
rect 6052 17768 7788 17796
rect 9267 17768 9312 17796
rect 6052 17756 6058 17768
rect 9306 17756 9312 17768
rect 9364 17756 9370 17808
rect 10244 17796 10272 17836
rect 13906 17824 13912 17836
rect 13964 17824 13970 17876
rect 15470 17824 15476 17876
rect 15528 17864 15534 17876
rect 15841 17867 15899 17873
rect 15841 17864 15853 17867
rect 15528 17836 15853 17864
rect 15528 17824 15534 17836
rect 15841 17833 15853 17836
rect 15887 17864 15899 17867
rect 15887 17836 16160 17864
rect 15887 17833 15899 17836
rect 15841 17827 15899 17833
rect 9968 17768 10272 17796
rect 4592 17731 4650 17737
rect 4592 17728 4604 17731
rect 4126 17700 4604 17728
rect 4592 17697 4604 17700
rect 4638 17728 4650 17731
rect 5166 17728 5172 17740
rect 4638 17700 5172 17728
rect 4638 17697 4650 17700
rect 4592 17691 4650 17697
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 9490 17688 9496 17740
rect 9548 17728 9554 17740
rect 9968 17737 9996 17768
rect 11514 17756 11520 17808
rect 11572 17796 11578 17808
rect 11609 17799 11667 17805
rect 11609 17796 11621 17799
rect 11572 17768 11621 17796
rect 11572 17756 11578 17768
rect 11609 17765 11621 17768
rect 11655 17765 11667 17799
rect 11609 17759 11667 17765
rect 12802 17756 12808 17808
rect 12860 17796 12866 17808
rect 13081 17799 13139 17805
rect 13081 17796 13093 17799
rect 12860 17768 13093 17796
rect 12860 17756 12866 17768
rect 13081 17765 13093 17768
rect 13127 17765 13139 17799
rect 13081 17759 13139 17765
rect 13173 17799 13231 17805
rect 13173 17765 13185 17799
rect 13219 17796 13231 17799
rect 13446 17796 13452 17808
rect 13219 17768 13452 17796
rect 13219 17765 13231 17768
rect 13173 17759 13231 17765
rect 13446 17756 13452 17768
rect 13504 17756 13510 17808
rect 13538 17756 13544 17808
rect 13596 17796 13602 17808
rect 13725 17799 13783 17805
rect 13725 17796 13737 17799
rect 13596 17768 13737 17796
rect 13596 17756 13602 17768
rect 13725 17765 13737 17768
rect 13771 17765 13783 17799
rect 13725 17759 13783 17765
rect 13814 17756 13820 17808
rect 13872 17796 13878 17808
rect 14550 17796 14556 17808
rect 13872 17768 14556 17796
rect 13872 17756 13878 17768
rect 14550 17756 14556 17768
rect 14608 17756 14614 17808
rect 16132 17805 16160 17836
rect 17494 17824 17500 17876
rect 17552 17864 17558 17876
rect 17681 17867 17739 17873
rect 17681 17864 17693 17867
rect 17552 17836 17693 17864
rect 17552 17824 17558 17836
rect 17681 17833 17693 17836
rect 17727 17833 17739 17867
rect 17681 17827 17739 17833
rect 18046 17824 18052 17876
rect 18104 17864 18110 17876
rect 19291 17867 19349 17873
rect 19291 17864 19303 17867
rect 18104 17836 19303 17864
rect 18104 17824 18110 17836
rect 19291 17833 19303 17836
rect 19337 17833 19349 17867
rect 19291 17827 19349 17833
rect 19518 17824 19524 17876
rect 19576 17864 19582 17876
rect 19613 17867 19671 17873
rect 19613 17864 19625 17867
rect 19576 17836 19625 17864
rect 19576 17824 19582 17836
rect 19613 17833 19625 17836
rect 19659 17833 19671 17867
rect 19613 17827 19671 17833
rect 16117 17799 16175 17805
rect 16117 17765 16129 17799
rect 16163 17765 16175 17799
rect 16117 17759 16175 17765
rect 16209 17799 16267 17805
rect 16209 17765 16221 17799
rect 16255 17796 16267 17799
rect 16298 17796 16304 17808
rect 16255 17768 16304 17796
rect 16255 17765 16267 17768
rect 16209 17759 16267 17765
rect 16298 17756 16304 17768
rect 16356 17756 16362 17808
rect 16761 17799 16819 17805
rect 16761 17765 16773 17799
rect 16807 17796 16819 17799
rect 18414 17796 18420 17808
rect 16807 17768 18420 17796
rect 16807 17765 16819 17768
rect 16761 17759 16819 17765
rect 18414 17756 18420 17768
rect 18472 17756 18478 17808
rect 9953 17731 10011 17737
rect 9953 17728 9965 17731
rect 9548 17700 9965 17728
rect 9548 17688 9554 17700
rect 9953 17697 9965 17700
rect 9999 17697 10011 17731
rect 10134 17728 10140 17740
rect 10095 17700 10140 17728
rect 9953 17691 10011 17697
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 17586 17728 17592 17740
rect 17547 17700 17592 17728
rect 17586 17688 17592 17700
rect 17644 17688 17650 17740
rect 17770 17688 17776 17740
rect 17828 17728 17834 17740
rect 18049 17731 18107 17737
rect 18049 17728 18061 17731
rect 17828 17700 18061 17728
rect 17828 17688 17834 17700
rect 18049 17697 18061 17700
rect 18095 17697 18107 17731
rect 19150 17728 19156 17740
rect 19111 17700 19156 17728
rect 18049 17691 18107 17697
rect 19150 17688 19156 17700
rect 19208 17688 19214 17740
rect 5534 17660 5540 17672
rect 5495 17632 5540 17660
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 6638 17620 6644 17672
rect 6696 17660 6702 17672
rect 7377 17663 7435 17669
rect 7377 17660 7389 17663
rect 6696 17632 7389 17660
rect 6696 17620 6702 17632
rect 7377 17629 7389 17632
rect 7423 17660 7435 17663
rect 10229 17663 10287 17669
rect 10229 17660 10241 17663
rect 7423 17632 10241 17660
rect 7423 17629 7435 17632
rect 7377 17623 7435 17629
rect 10229 17629 10241 17632
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 11330 17620 11336 17672
rect 11388 17660 11394 17672
rect 11517 17663 11575 17669
rect 11517 17660 11529 17663
rect 11388 17632 11529 17660
rect 11388 17620 11394 17632
rect 11517 17629 11529 17632
rect 11563 17629 11575 17663
rect 11882 17660 11888 17672
rect 11843 17632 11888 17660
rect 11517 17623 11575 17629
rect 11882 17620 11888 17632
rect 11940 17620 11946 17672
rect 15194 17660 15200 17672
rect 13188 17632 15200 17660
rect 2498 17592 2504 17604
rect 2411 17564 2504 17592
rect 2498 17552 2504 17564
rect 2556 17592 2562 17604
rect 3510 17592 3516 17604
rect 2556 17564 3516 17592
rect 2556 17552 2562 17564
rect 3510 17552 3516 17564
rect 3568 17552 3574 17604
rect 4663 17595 4721 17601
rect 4663 17561 4675 17595
rect 4709 17592 4721 17595
rect 11606 17592 11612 17604
rect 4709 17564 11612 17592
rect 4709 17561 4721 17564
rect 4663 17555 4721 17561
rect 11606 17552 11612 17564
rect 11664 17552 11670 17604
rect 12526 17592 12532 17604
rect 12439 17564 12532 17592
rect 12526 17552 12532 17564
rect 12584 17592 12590 17604
rect 13188 17592 13216 17632
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 12584 17564 13216 17592
rect 12584 17552 12590 17564
rect 2133 17527 2191 17533
rect 2133 17493 2145 17527
rect 2179 17524 2191 17527
rect 2866 17524 2872 17536
rect 2179 17496 2872 17524
rect 2179 17493 2191 17496
rect 2133 17487 2191 17493
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 3142 17524 3148 17536
rect 3103 17496 3148 17524
rect 3142 17484 3148 17496
rect 3200 17484 3206 17536
rect 3418 17524 3424 17536
rect 3379 17496 3424 17524
rect 3418 17484 3424 17496
rect 3476 17484 3482 17536
rect 4062 17484 4068 17536
rect 4120 17524 4126 17536
rect 4249 17527 4307 17533
rect 4249 17524 4261 17527
rect 4120 17496 4261 17524
rect 4120 17484 4126 17496
rect 4249 17493 4261 17496
rect 4295 17493 4307 17527
rect 4249 17487 4307 17493
rect 6730 17484 6736 17536
rect 6788 17524 6794 17536
rect 7193 17527 7251 17533
rect 7193 17524 7205 17527
rect 6788 17496 7205 17524
rect 6788 17484 6794 17496
rect 7193 17493 7205 17496
rect 7239 17493 7251 17527
rect 7193 17487 7251 17493
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 8573 17527 8631 17533
rect 8573 17524 8585 17527
rect 7984 17496 8585 17524
rect 7984 17484 7990 17496
rect 8573 17493 8585 17496
rect 8619 17524 8631 17527
rect 9030 17524 9036 17536
rect 8619 17496 9036 17524
rect 8619 17493 8631 17496
rect 8573 17487 8631 17493
rect 9030 17484 9036 17496
rect 9088 17484 9094 17536
rect 10686 17524 10692 17536
rect 10647 17496 10692 17524
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 12618 17484 12624 17536
rect 12676 17524 12682 17536
rect 12897 17527 12955 17533
rect 12897 17524 12909 17527
rect 12676 17496 12909 17524
rect 12676 17484 12682 17496
rect 12897 17493 12909 17496
rect 12943 17524 12955 17527
rect 13354 17524 13360 17536
rect 12943 17496 13360 17524
rect 12943 17493 12955 17496
rect 12897 17487 12955 17493
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 17126 17484 17132 17536
rect 17184 17524 17190 17536
rect 17405 17527 17463 17533
rect 17405 17524 17417 17527
rect 17184 17496 17417 17524
rect 17184 17484 17190 17496
rect 17405 17493 17417 17496
rect 17451 17493 17463 17527
rect 18598 17524 18604 17536
rect 18559 17496 18604 17524
rect 17405 17487 17463 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 18966 17524 18972 17536
rect 18927 17496 18972 17524
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2041 17323 2099 17329
rect 2041 17289 2053 17323
rect 2087 17320 2099 17323
rect 3050 17320 3056 17332
rect 2087 17292 3056 17320
rect 2087 17289 2099 17292
rect 2041 17283 2099 17289
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2056 17116 2084 17283
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 3326 17320 3332 17332
rect 3287 17292 3332 17320
rect 3326 17280 3332 17292
rect 3384 17320 3390 17332
rect 4614 17320 4620 17332
rect 3384 17292 4620 17320
rect 3384 17280 3390 17292
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 4798 17320 4804 17332
rect 4759 17292 4804 17320
rect 4798 17280 4804 17292
rect 4856 17280 4862 17332
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 6181 17323 6239 17329
rect 6181 17320 6193 17323
rect 5592 17292 6193 17320
rect 5592 17280 5598 17292
rect 6181 17289 6193 17292
rect 6227 17289 6239 17323
rect 6638 17320 6644 17332
rect 6599 17292 6644 17320
rect 6181 17283 6239 17289
rect 6638 17280 6644 17292
rect 6696 17280 6702 17332
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 7101 17323 7159 17329
rect 7101 17320 7113 17323
rect 6972 17292 7113 17320
rect 6972 17280 6978 17292
rect 7101 17289 7113 17292
rect 7147 17289 7159 17323
rect 7101 17283 7159 17289
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 9861 17323 9919 17329
rect 9861 17320 9873 17323
rect 7432 17292 9873 17320
rect 7432 17280 7438 17292
rect 9861 17289 9873 17292
rect 9907 17320 9919 17323
rect 10134 17320 10140 17332
rect 9907 17292 10140 17320
rect 9907 17289 9919 17292
rect 9861 17283 9919 17289
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 11514 17320 11520 17332
rect 11475 17292 11520 17320
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 12802 17280 12808 17332
rect 12860 17320 12866 17332
rect 13817 17323 13875 17329
rect 13817 17320 13829 17323
rect 12860 17292 13829 17320
rect 12860 17280 12866 17292
rect 13817 17289 13829 17292
rect 13863 17289 13875 17323
rect 15654 17320 15660 17332
rect 15615 17292 15660 17320
rect 13817 17283 13875 17289
rect 15654 17280 15660 17292
rect 15712 17320 15718 17332
rect 16298 17320 16304 17332
rect 15712 17292 16304 17320
rect 15712 17280 15718 17292
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 19978 17280 19984 17332
rect 20036 17320 20042 17332
rect 20073 17323 20131 17329
rect 20073 17320 20085 17323
rect 20036 17292 20085 17320
rect 20036 17280 20042 17292
rect 20073 17289 20085 17292
rect 20119 17289 20131 17323
rect 20073 17283 20131 17289
rect 4893 17255 4951 17261
rect 4893 17221 4905 17255
rect 4939 17252 4951 17255
rect 5629 17255 5687 17261
rect 5629 17252 5641 17255
rect 4939 17224 5641 17252
rect 4939 17221 4951 17224
rect 4893 17215 4951 17221
rect 5629 17221 5641 17224
rect 5675 17252 5687 17255
rect 5994 17252 6000 17264
rect 5675 17224 6000 17252
rect 5675 17221 5687 17224
rect 5629 17215 5687 17221
rect 5994 17212 6000 17224
rect 6052 17212 6058 17264
rect 11241 17255 11299 17261
rect 11241 17221 11253 17255
rect 11287 17252 11299 17255
rect 11422 17252 11428 17264
rect 11287 17224 11428 17252
rect 11287 17221 11299 17224
rect 11241 17215 11299 17221
rect 11422 17212 11428 17224
rect 11480 17252 11486 17264
rect 13446 17252 13452 17264
rect 11480 17224 13452 17252
rect 11480 17212 11486 17224
rect 13446 17212 13452 17224
rect 13504 17212 13510 17264
rect 24765 17255 24823 17261
rect 24765 17221 24777 17255
rect 24811 17252 24823 17255
rect 27614 17252 27620 17264
rect 24811 17224 27620 17252
rect 24811 17221 24823 17224
rect 24765 17215 24823 17221
rect 27614 17212 27620 17224
rect 27672 17212 27678 17264
rect 5721 17187 5779 17193
rect 2884 17156 5672 17184
rect 2884 17125 2912 17156
rect 1443 17088 2084 17116
rect 2777 17119 2835 17125
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 2777 17085 2789 17119
rect 2823 17116 2835 17119
rect 2869 17119 2927 17125
rect 2869 17116 2881 17119
rect 2823 17088 2881 17116
rect 2823 17085 2835 17088
rect 2777 17079 2835 17085
rect 2869 17085 2881 17088
rect 2915 17085 2927 17119
rect 2869 17079 2927 17085
rect 3881 17119 3939 17125
rect 3881 17085 3893 17119
rect 3927 17116 3939 17119
rect 4062 17116 4068 17128
rect 3927 17088 4068 17116
rect 3927 17085 3939 17088
rect 3881 17079 3939 17085
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 5644 17116 5672 17156
rect 5721 17153 5733 17187
rect 5767 17184 5779 17187
rect 6546 17184 6552 17196
rect 5767 17156 6552 17184
rect 5767 17153 5779 17156
rect 5721 17147 5779 17153
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 9398 17184 9404 17196
rect 6748 17156 6960 17184
rect 6270 17116 6276 17128
rect 5644 17088 6276 17116
rect 6270 17076 6276 17088
rect 6328 17076 6334 17128
rect 6748 17125 6776 17156
rect 6932 17128 6960 17156
rect 7300 17156 9404 17184
rect 6733 17119 6791 17125
rect 6733 17085 6745 17119
rect 6779 17085 6791 17119
rect 6733 17079 6791 17085
rect 6914 17076 6920 17128
rect 6972 17116 6978 17128
rect 7300 17125 7328 17156
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17184 9551 17187
rect 10321 17187 10379 17193
rect 10321 17184 10333 17187
rect 9539 17156 10333 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 10321 17153 10333 17156
rect 10367 17184 10379 17187
rect 10686 17184 10692 17196
rect 10367 17156 10692 17184
rect 10367 17153 10379 17156
rect 10321 17147 10379 17153
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 12526 17184 12532 17196
rect 12487 17156 12532 17184
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 12802 17184 12808 17196
rect 12763 17156 12808 17184
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17184 15347 17187
rect 16206 17184 16212 17196
rect 15335 17156 16212 17184
rect 15335 17153 15347 17156
rect 15289 17147 15347 17153
rect 16206 17144 16212 17156
rect 16264 17144 16270 17196
rect 18233 17187 18291 17193
rect 18233 17153 18245 17187
rect 18279 17184 18291 17187
rect 18966 17184 18972 17196
rect 18279 17156 18972 17184
rect 18279 17153 18291 17156
rect 18233 17147 18291 17153
rect 18966 17144 18972 17156
rect 19024 17144 19030 17196
rect 7285 17119 7343 17125
rect 7285 17116 7297 17119
rect 6972 17088 7297 17116
rect 6972 17076 6978 17088
rect 7285 17085 7297 17088
rect 7331 17085 7343 17119
rect 7285 17079 7343 17085
rect 7926 17076 7932 17128
rect 7984 17116 7990 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7984 17088 8033 17116
rect 7984 17076 7990 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 8110 17076 8116 17128
rect 8168 17116 8174 17128
rect 8481 17119 8539 17125
rect 8481 17116 8493 17119
rect 8168 17088 8493 17116
rect 8168 17076 8174 17088
rect 8481 17085 8493 17088
rect 8527 17085 8539 17119
rect 8938 17116 8944 17128
rect 8899 17088 8944 17116
rect 8481 17079 8539 17085
rect 8938 17076 8944 17088
rect 8996 17076 9002 17128
rect 9214 17116 9220 17128
rect 9175 17088 9220 17116
rect 9214 17076 9220 17088
rect 9272 17076 9278 17128
rect 10134 17076 10140 17128
rect 10192 17116 10198 17128
rect 14550 17116 14556 17128
rect 10192 17088 10726 17116
rect 14511 17088 14556 17116
rect 10192 17076 10198 17088
rect 3418 17008 3424 17060
rect 3476 17048 3482 17060
rect 3697 17051 3755 17057
rect 3697 17048 3709 17051
rect 3476 17020 3709 17048
rect 3476 17008 3482 17020
rect 3697 17017 3709 17020
rect 3743 17048 3755 17051
rect 4243 17051 4301 17057
rect 4243 17048 4255 17051
rect 3743 17020 4255 17048
rect 3743 17017 3755 17020
rect 3697 17011 3755 17017
rect 4243 17017 4255 17020
rect 4289 17048 4301 17051
rect 4893 17051 4951 17057
rect 4893 17048 4905 17051
rect 4289 17020 4905 17048
rect 4289 17017 4301 17020
rect 4243 17011 4301 17017
rect 4893 17017 4905 17020
rect 4939 17017 4951 17051
rect 5166 17048 5172 17060
rect 5079 17020 5172 17048
rect 4893 17011 4951 17017
rect 5166 17008 5172 17020
rect 5224 17048 5230 17060
rect 10698 17057 10726 17088
rect 14550 17076 14556 17088
rect 14608 17076 14614 17128
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17085 15071 17119
rect 15013 17079 15071 17085
rect 10683 17051 10741 17057
rect 5224 17020 10594 17048
rect 5224 17008 5230 17020
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 2406 16980 2412 16992
rect 2367 16952 2412 16980
rect 2406 16940 2412 16952
rect 2464 16940 2470 16992
rect 3053 16983 3111 16989
rect 3053 16949 3065 16983
rect 3099 16980 3111 16983
rect 3602 16980 3608 16992
rect 3099 16952 3608 16980
rect 3099 16949 3111 16952
rect 3053 16943 3111 16949
rect 3602 16940 3608 16952
rect 3660 16940 3666 16992
rect 7742 16980 7748 16992
rect 7655 16952 7748 16980
rect 7742 16940 7748 16952
rect 7800 16980 7806 16992
rect 10134 16980 10140 16992
rect 7800 16952 10140 16980
rect 7800 16940 7806 16952
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 10566 16980 10594 17020
rect 10683 17017 10695 17051
rect 10729 17017 10741 17051
rect 12250 17048 12256 17060
rect 12163 17020 12256 17048
rect 10683 17011 10741 17017
rect 12250 17008 12256 17020
rect 12308 17048 12314 17060
rect 12618 17048 12624 17060
rect 12308 17020 12624 17048
rect 12308 17008 12314 17020
rect 12618 17008 12624 17020
rect 12676 17008 12682 17060
rect 15028 17048 15056 17079
rect 16022 17076 16028 17128
rect 16080 17116 16086 17128
rect 16117 17119 16175 17125
rect 16117 17116 16129 17119
rect 16080 17088 16129 17116
rect 16080 17076 16086 17088
rect 16117 17085 16129 17088
rect 16163 17085 16175 17119
rect 16117 17079 16175 17085
rect 18874 17076 18880 17128
rect 18932 17116 18938 17128
rect 19864 17119 19922 17125
rect 19864 17116 19876 17119
rect 18932 17088 19876 17116
rect 18932 17076 18938 17088
rect 19864 17085 19876 17088
rect 19910 17116 19922 17119
rect 20257 17119 20315 17125
rect 20257 17116 20269 17119
rect 19910 17088 20269 17116
rect 19910 17085 19922 17088
rect 19864 17079 19922 17085
rect 20257 17085 20269 17088
rect 20303 17085 20315 17119
rect 20257 17079 20315 17085
rect 24210 17076 24216 17128
rect 24268 17116 24274 17128
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 24268 17088 24593 17116
rect 24268 17076 24274 17088
rect 24581 17085 24593 17088
rect 24627 17116 24639 17119
rect 25133 17119 25191 17125
rect 25133 17116 25145 17119
rect 24627 17088 25145 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 25133 17085 25145 17088
rect 25179 17085 25191 17119
rect 25133 17079 25191 17085
rect 16438 17051 16496 17057
rect 16438 17048 16450 17051
rect 14568 17020 15056 17048
rect 15948 17020 16450 17048
rect 14568 16992 14596 17020
rect 12526 16980 12532 16992
rect 10566 16952 12532 16980
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 14461 16983 14519 16989
rect 14461 16949 14473 16983
rect 14507 16980 14519 16983
rect 14550 16980 14556 16992
rect 14507 16952 14556 16980
rect 14507 16949 14519 16952
rect 14461 16943 14519 16949
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 15948 16989 15976 17020
rect 16438 17017 16450 17020
rect 16484 17048 16496 17051
rect 16758 17048 16764 17060
rect 16484 17020 16764 17048
rect 16484 17017 16496 17020
rect 16438 17011 16496 17017
rect 16758 17008 16764 17020
rect 16816 17008 16822 17060
rect 18325 17051 18383 17057
rect 18325 17017 18337 17051
rect 18371 17048 18383 17051
rect 18598 17048 18604 17060
rect 18371 17020 18604 17048
rect 18371 17017 18383 17020
rect 18325 17011 18383 17017
rect 18598 17008 18604 17020
rect 18656 17008 18662 17060
rect 15933 16983 15991 16989
rect 15933 16980 15945 16983
rect 15528 16952 15945 16980
rect 15528 16940 15534 16952
rect 15933 16949 15945 16952
rect 15979 16949 15991 16983
rect 17034 16980 17040 16992
rect 16995 16952 17040 16980
rect 15933 16943 15991 16949
rect 17034 16940 17040 16952
rect 17092 16940 17098 16992
rect 17586 16980 17592 16992
rect 17547 16952 17592 16980
rect 17586 16940 17592 16952
rect 17644 16940 17650 16992
rect 17678 16940 17684 16992
rect 17736 16980 17742 16992
rect 19150 16980 19156 16992
rect 17736 16952 19156 16980
rect 17736 16940 17742 16952
rect 19150 16940 19156 16952
rect 19208 16940 19214 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 3142 16736 3148 16788
rect 3200 16776 3206 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 3200 16748 3801 16776
rect 3200 16736 3206 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 3789 16739 3847 16745
rect 2866 16668 2872 16720
rect 2924 16708 2930 16720
rect 3804 16708 3832 16739
rect 4062 16736 4068 16788
rect 4120 16776 4126 16788
rect 4157 16779 4215 16785
rect 4157 16776 4169 16779
rect 4120 16748 4169 16776
rect 4120 16736 4126 16748
rect 4157 16745 4169 16748
rect 4203 16745 4215 16779
rect 8018 16776 8024 16788
rect 4157 16739 4215 16745
rect 4724 16748 8024 16776
rect 4724 16708 4752 16748
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 8481 16779 8539 16785
rect 8481 16745 8493 16779
rect 8527 16776 8539 16779
rect 9214 16776 9220 16788
rect 8527 16748 9220 16776
rect 8527 16745 8539 16748
rect 8481 16739 8539 16745
rect 8496 16708 8524 16739
rect 9214 16736 9220 16748
rect 9272 16736 9278 16788
rect 9490 16776 9496 16788
rect 9451 16748 9496 16776
rect 9490 16736 9496 16748
rect 9548 16736 9554 16788
rect 10134 16776 10140 16788
rect 10095 16748 10140 16776
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 10689 16779 10747 16785
rect 10689 16745 10701 16779
rect 10735 16745 10747 16779
rect 11330 16776 11336 16788
rect 11291 16748 11336 16776
rect 10689 16739 10747 16745
rect 9030 16708 9036 16720
rect 2924 16680 3740 16708
rect 3804 16680 4752 16708
rect 2924 16668 2930 16680
rect 1946 16640 1952 16652
rect 1907 16612 1952 16640
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 2774 16600 2780 16652
rect 2832 16640 2838 16652
rect 2996 16643 3054 16649
rect 2996 16640 3008 16643
rect 2832 16612 3008 16640
rect 2832 16600 2838 16612
rect 2996 16609 3008 16612
rect 3042 16609 3054 16643
rect 3712 16640 3740 16680
rect 4724 16652 4752 16680
rect 5460 16680 8524 16708
rect 8991 16680 9036 16708
rect 4062 16640 4068 16652
rect 3712 16612 4068 16640
rect 2996 16603 3054 16609
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 4706 16640 4712 16652
rect 4619 16612 4712 16640
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 4890 16640 4896 16652
rect 4851 16612 4896 16640
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 5460 16649 5488 16680
rect 9030 16668 9036 16680
rect 9088 16668 9094 16720
rect 10704 16708 10732 16739
rect 11330 16736 11336 16748
rect 11388 16776 11394 16788
rect 12802 16776 12808 16788
rect 11388 16748 12808 16776
rect 11388 16736 11394 16748
rect 11701 16711 11759 16717
rect 11701 16708 11713 16711
rect 10704 16680 11713 16708
rect 11701 16677 11713 16680
rect 11747 16708 11759 16711
rect 11790 16708 11796 16720
rect 11747 16680 11796 16708
rect 11747 16677 11759 16680
rect 11701 16671 11759 16677
rect 11790 16668 11796 16680
rect 11848 16668 11854 16720
rect 12268 16717 12296 16748
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 16758 16776 16764 16788
rect 16719 16748 16764 16776
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 17313 16779 17371 16785
rect 17313 16745 17325 16779
rect 17359 16776 17371 16779
rect 18598 16776 18604 16788
rect 17359 16748 18604 16776
rect 17359 16745 17371 16748
rect 17313 16739 17371 16745
rect 18598 16736 18604 16748
rect 18656 16736 18662 16788
rect 19518 16736 19524 16788
rect 19576 16776 19582 16788
rect 19705 16779 19763 16785
rect 19705 16776 19717 16779
rect 19576 16748 19717 16776
rect 19576 16736 19582 16748
rect 19705 16745 19717 16748
rect 19751 16745 19763 16779
rect 19705 16739 19763 16745
rect 12253 16711 12311 16717
rect 12253 16677 12265 16711
rect 12299 16677 12311 16711
rect 12253 16671 12311 16677
rect 12618 16668 12624 16720
rect 12676 16708 12682 16720
rect 13081 16711 13139 16717
rect 13081 16708 13093 16711
rect 12676 16680 13093 16708
rect 12676 16668 12682 16680
rect 13081 16677 13093 16680
rect 13127 16677 13139 16711
rect 13081 16671 13139 16677
rect 16942 16668 16948 16720
rect 17000 16708 17006 16720
rect 18325 16711 18383 16717
rect 18325 16708 18337 16711
rect 17000 16680 18337 16708
rect 17000 16668 17006 16680
rect 18325 16677 18337 16680
rect 18371 16708 18383 16711
rect 18690 16708 18696 16720
rect 18371 16680 18696 16708
rect 18371 16677 18383 16680
rect 18325 16671 18383 16677
rect 18690 16668 18696 16680
rect 18748 16668 18754 16720
rect 18874 16708 18880 16720
rect 18835 16680 18880 16708
rect 18874 16668 18880 16680
rect 18932 16668 18938 16720
rect 5445 16643 5503 16649
rect 5445 16609 5457 16643
rect 5491 16609 5503 16643
rect 5445 16603 5503 16609
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16609 7251 16643
rect 7374 16640 7380 16652
rect 7335 16612 7380 16640
rect 7193 16603 7251 16609
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16572 2191 16575
rect 2222 16572 2228 16584
rect 2179 16544 2228 16572
rect 2179 16541 2191 16544
rect 2133 16535 2191 16541
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 2406 16532 2412 16584
rect 2464 16572 2470 16584
rect 5350 16572 5356 16584
rect 2464 16544 5356 16572
rect 2464 16532 2470 16544
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 1762 16464 1768 16516
rect 1820 16504 1826 16516
rect 2777 16507 2835 16513
rect 2777 16504 2789 16507
rect 1820 16476 2789 16504
rect 1820 16464 1826 16476
rect 2777 16473 2789 16476
rect 2823 16504 2835 16507
rect 3099 16507 3157 16513
rect 3099 16504 3111 16507
rect 2823 16476 3111 16504
rect 2823 16473 2835 16476
rect 2777 16467 2835 16473
rect 3099 16473 3111 16476
rect 3145 16473 3157 16507
rect 5460 16504 5488 16603
rect 3099 16467 3157 16473
rect 3436 16476 5488 16504
rect 7208 16504 7236 16603
rect 7374 16600 7380 16612
rect 7432 16600 7438 16652
rect 8570 16640 8576 16652
rect 8531 16612 8576 16640
rect 8570 16600 8576 16612
rect 8628 16600 8634 16652
rect 13446 16640 13452 16652
rect 13407 16612 13452 16640
rect 13446 16600 13452 16612
rect 13504 16600 13510 16652
rect 15197 16643 15255 16649
rect 15197 16609 15209 16643
rect 15243 16640 15255 16643
rect 15286 16640 15292 16652
rect 15243 16612 15292 16640
rect 15243 16609 15255 16612
rect 15197 16603 15255 16609
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 16393 16643 16451 16649
rect 16393 16609 16405 16643
rect 16439 16640 16451 16643
rect 17494 16640 17500 16652
rect 16439 16612 17500 16640
rect 16439 16609 16451 16612
rect 16393 16603 16451 16609
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 24489 16643 24547 16649
rect 24489 16609 24501 16643
rect 24535 16640 24547 16643
rect 24670 16640 24676 16652
rect 24535 16612 24676 16640
rect 24535 16609 24547 16612
rect 24489 16603 24547 16609
rect 24670 16600 24676 16612
rect 24728 16600 24734 16652
rect 7466 16572 7472 16584
rect 7427 16544 7472 16572
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 9490 16532 9496 16584
rect 9548 16572 9554 16584
rect 9769 16575 9827 16581
rect 9769 16572 9781 16575
rect 9548 16544 9781 16572
rect 9548 16532 9554 16544
rect 9769 16541 9781 16544
rect 9815 16572 9827 16575
rect 10965 16575 11023 16581
rect 10965 16572 10977 16575
rect 9815 16544 10977 16572
rect 9815 16541 9827 16544
rect 9769 16535 9827 16541
rect 10965 16541 10977 16544
rect 11011 16541 11023 16575
rect 11606 16572 11612 16584
rect 11567 16544 11612 16572
rect 10965 16535 11023 16541
rect 11606 16532 11612 16544
rect 11664 16532 11670 16584
rect 18233 16575 18291 16581
rect 18233 16541 18245 16575
rect 18279 16572 18291 16575
rect 18414 16572 18420 16584
rect 18279 16544 18420 16572
rect 18279 16541 18291 16544
rect 18233 16535 18291 16541
rect 18414 16532 18420 16544
rect 18472 16532 18478 16584
rect 7742 16504 7748 16516
rect 7208 16476 7748 16504
rect 1946 16396 1952 16448
rect 2004 16436 2010 16448
rect 2409 16439 2467 16445
rect 2409 16436 2421 16439
rect 2004 16408 2421 16436
rect 2004 16396 2010 16408
rect 2409 16405 2421 16408
rect 2455 16405 2467 16439
rect 2409 16399 2467 16405
rect 3326 16396 3332 16448
rect 3384 16436 3390 16448
rect 3436 16445 3464 16476
rect 7742 16464 7748 16476
rect 7800 16464 7806 16516
rect 8757 16507 8815 16513
rect 8757 16473 8769 16507
rect 8803 16504 8815 16507
rect 9950 16504 9956 16516
rect 8803 16476 9956 16504
rect 8803 16473 8815 16476
rect 8757 16467 8815 16473
rect 9950 16464 9956 16476
rect 10008 16464 10014 16516
rect 15427 16507 15485 16513
rect 15427 16473 15439 16507
rect 15473 16504 15485 16507
rect 17218 16504 17224 16516
rect 15473 16476 17224 16504
rect 15473 16473 15485 16476
rect 15427 16467 15485 16473
rect 17218 16464 17224 16476
rect 17276 16464 17282 16516
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 3384 16408 3433 16436
rect 3384 16396 3390 16408
rect 3421 16405 3433 16408
rect 3467 16405 3479 16439
rect 8018 16436 8024 16448
rect 7979 16408 8024 16436
rect 3421 16399 3479 16405
rect 8018 16396 8024 16408
rect 8076 16396 8082 16448
rect 14369 16439 14427 16445
rect 14369 16405 14381 16439
rect 14415 16436 14427 16439
rect 14826 16436 14832 16448
rect 14415 16408 14832 16436
rect 14415 16405 14427 16408
rect 14369 16399 14427 16405
rect 14826 16396 14832 16408
rect 14884 16396 14890 16448
rect 15838 16436 15844 16448
rect 15799 16408 15844 16436
rect 15838 16396 15844 16408
rect 15896 16396 15902 16448
rect 16022 16396 16028 16448
rect 16080 16436 16086 16448
rect 16117 16439 16175 16445
rect 16117 16436 16129 16439
rect 16080 16408 16129 16436
rect 16080 16396 16086 16408
rect 16117 16405 16129 16408
rect 16163 16405 16175 16439
rect 16117 16399 16175 16405
rect 17681 16439 17739 16445
rect 17681 16405 17693 16439
rect 17727 16436 17739 16439
rect 17770 16436 17776 16448
rect 17727 16408 17776 16436
rect 17727 16405 17739 16408
rect 17681 16399 17739 16405
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 18046 16436 18052 16448
rect 18007 16408 18052 16436
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 21358 16436 21364 16448
rect 21271 16408 21364 16436
rect 21358 16396 21364 16408
rect 21416 16436 21422 16448
rect 24719 16439 24777 16445
rect 24719 16436 24731 16439
rect 21416 16408 24731 16436
rect 21416 16396 21422 16408
rect 24719 16405 24731 16408
rect 24765 16405 24777 16439
rect 24719 16399 24777 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2774 16192 2780 16244
rect 2832 16232 2838 16244
rect 2961 16235 3019 16241
rect 2961 16232 2973 16235
rect 2832 16204 2973 16232
rect 2832 16192 2838 16204
rect 2961 16201 2973 16204
rect 3007 16232 3019 16235
rect 6546 16232 6552 16244
rect 3007 16204 6552 16232
rect 3007 16201 3019 16204
rect 2961 16195 3019 16201
rect 6546 16192 6552 16204
rect 6604 16192 6610 16244
rect 7147 16235 7205 16241
rect 7147 16201 7159 16235
rect 7193 16232 7205 16235
rect 11238 16232 11244 16244
rect 7193 16204 11244 16232
rect 7193 16201 7205 16204
rect 7147 16195 7205 16201
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 11790 16232 11796 16244
rect 11703 16204 11796 16232
rect 11790 16192 11796 16204
rect 11848 16232 11854 16244
rect 13446 16232 13452 16244
rect 11848 16204 13452 16232
rect 11848 16192 11854 16204
rect 13446 16192 13452 16204
rect 13504 16192 13510 16244
rect 15286 16232 15292 16244
rect 15247 16204 15292 16232
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 16761 16235 16819 16241
rect 16761 16201 16773 16235
rect 16807 16232 16819 16235
rect 16942 16232 16948 16244
rect 16807 16204 16948 16232
rect 16807 16201 16819 16204
rect 16761 16195 16819 16201
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 17034 16192 17040 16244
rect 17092 16232 17098 16244
rect 17773 16235 17831 16241
rect 17773 16232 17785 16235
rect 17092 16204 17785 16232
rect 17092 16192 17098 16204
rect 17773 16201 17785 16204
rect 17819 16232 17831 16235
rect 18322 16232 18328 16244
rect 17819 16204 18328 16232
rect 17819 16201 17831 16204
rect 17773 16195 17831 16201
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 18690 16192 18696 16244
rect 18748 16232 18754 16244
rect 19153 16235 19211 16241
rect 19153 16232 19165 16235
rect 18748 16204 19165 16232
rect 18748 16192 18754 16204
rect 19153 16201 19165 16204
rect 19199 16201 19211 16235
rect 24670 16232 24676 16244
rect 24631 16204 24676 16232
rect 19153 16195 19211 16201
rect 24670 16192 24676 16204
rect 24728 16192 24734 16244
rect 4062 16124 4068 16176
rect 4120 16164 4126 16176
rect 5721 16167 5779 16173
rect 5721 16164 5733 16167
rect 4120 16136 5733 16164
rect 4120 16124 4126 16136
rect 5721 16133 5733 16136
rect 5767 16133 5779 16167
rect 5721 16127 5779 16133
rect 6641 16167 6699 16173
rect 6641 16133 6653 16167
rect 6687 16164 6699 16167
rect 7374 16164 7380 16176
rect 6687 16136 7380 16164
rect 6687 16133 6699 16136
rect 6641 16127 6699 16133
rect 7374 16124 7380 16136
rect 7432 16124 7438 16176
rect 9861 16167 9919 16173
rect 9861 16133 9873 16167
rect 9907 16164 9919 16167
rect 10134 16164 10140 16176
rect 9907 16136 10140 16164
rect 9907 16133 9919 16136
rect 9861 16127 9919 16133
rect 10134 16124 10140 16136
rect 10192 16124 10198 16176
rect 11333 16167 11391 16173
rect 11333 16164 11345 16167
rect 10336 16136 11345 16164
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 6917 16099 6975 16105
rect 2731 16068 5396 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 4062 16028 4068 16040
rect 4023 16000 4068 16028
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 4706 16028 4712 16040
rect 4667 16000 4712 16028
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 4890 16028 4896 16040
rect 4851 16000 4896 16028
rect 4890 15988 4896 16000
rect 4948 15988 4954 16040
rect 5368 16037 5396 16068
rect 6917 16065 6929 16099
rect 6963 16096 6975 16099
rect 9490 16096 9496 16108
rect 6963 16068 7328 16096
rect 9451 16068 9496 16096
rect 6963 16065 6975 16068
rect 6917 16059 6975 16065
rect 7300 16040 7328 16068
rect 9490 16056 9496 16068
rect 9548 16056 9554 16108
rect 5353 16031 5411 16037
rect 5353 15997 5365 16031
rect 5399 16028 5411 16031
rect 5994 16028 6000 16040
rect 5399 16000 6000 16028
rect 5399 15997 5411 16000
rect 5353 15991 5411 15997
rect 5994 15988 6000 16000
rect 6052 15988 6058 16040
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 7340 16000 7481 16028
rect 7340 15988 7346 16000
rect 7469 15997 7481 16000
rect 7515 15997 7527 16031
rect 7469 15991 7527 15997
rect 7926 15988 7932 16040
rect 7984 16028 7990 16040
rect 8021 16031 8079 16037
rect 8021 16028 8033 16031
rect 7984 16000 8033 16028
rect 7984 15988 7990 16000
rect 8021 15997 8033 16000
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 8481 16031 8539 16037
rect 8481 15997 8493 16031
rect 8527 15997 8539 16031
rect 8938 16028 8944 16040
rect 8899 16000 8944 16028
rect 8481 15991 8539 15997
rect 1765 15963 1823 15969
rect 1765 15929 1777 15963
rect 1811 15960 1823 15963
rect 1946 15960 1952 15972
rect 1811 15932 1952 15960
rect 1811 15929 1823 15932
rect 1765 15923 1823 15929
rect 1946 15920 1952 15932
rect 2004 15920 2010 15972
rect 2317 15963 2375 15969
rect 2317 15929 2329 15963
rect 2363 15960 2375 15963
rect 2406 15960 2412 15972
rect 2363 15932 2412 15960
rect 2363 15929 2375 15932
rect 2317 15923 2375 15929
rect 2406 15920 2412 15932
rect 2464 15920 2470 15972
rect 3513 15963 3571 15969
rect 3513 15929 3525 15963
rect 3559 15960 3571 15963
rect 3786 15960 3792 15972
rect 3559 15932 3792 15960
rect 3559 15929 3571 15932
rect 3513 15923 3571 15929
rect 3786 15920 3792 15932
rect 3844 15960 3850 15972
rect 4908 15960 4936 15988
rect 3844 15932 4936 15960
rect 6273 15963 6331 15969
rect 3844 15920 3850 15932
rect 6273 15929 6285 15963
rect 6319 15960 6331 15963
rect 7742 15960 7748 15972
rect 6319 15932 7748 15960
rect 6319 15929 6331 15932
rect 6273 15923 6331 15929
rect 7742 15920 7748 15932
rect 7800 15920 7806 15972
rect 8496 15960 8524 15991
rect 8938 15988 8944 16000
rect 8996 15988 9002 16040
rect 9122 15988 9128 16040
rect 9180 16028 9186 16040
rect 9217 16031 9275 16037
rect 9217 16028 9229 16031
rect 9180 16000 9229 16028
rect 9180 15988 9186 16000
rect 9217 15997 9229 16000
rect 9263 15997 9275 16031
rect 9217 15991 9275 15997
rect 9858 15988 9864 16040
rect 9916 16028 9922 16040
rect 10336 16037 10364 16136
rect 11333 16133 11345 16136
rect 11379 16133 11391 16167
rect 17494 16164 17500 16176
rect 17455 16136 17500 16164
rect 11333 16127 11391 16133
rect 17494 16124 17500 16136
rect 17552 16124 17558 16176
rect 20088 16136 21680 16164
rect 11054 16096 11060 16108
rect 11015 16068 11060 16096
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 18046 16056 18052 16108
rect 18104 16096 18110 16108
rect 18230 16096 18236 16108
rect 18104 16068 18236 16096
rect 18104 16056 18110 16068
rect 18230 16056 18236 16068
rect 18288 16056 18294 16108
rect 18874 16096 18880 16108
rect 18835 16068 18880 16096
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 18966 16056 18972 16108
rect 19024 16096 19030 16108
rect 19978 16096 19984 16108
rect 19024 16068 19984 16096
rect 19024 16056 19030 16068
rect 19978 16056 19984 16068
rect 20036 16096 20042 16108
rect 20088 16105 20116 16136
rect 20073 16099 20131 16105
rect 20073 16096 20085 16099
rect 20036 16068 20085 16096
rect 20036 16056 20042 16068
rect 20073 16065 20085 16068
rect 20119 16065 20131 16099
rect 21358 16096 21364 16108
rect 21319 16068 21364 16096
rect 20073 16059 20131 16065
rect 21358 16056 21364 16068
rect 21416 16056 21422 16108
rect 21652 16105 21680 16136
rect 21637 16099 21695 16105
rect 21637 16065 21649 16099
rect 21683 16065 21695 16099
rect 21637 16059 21695 16065
rect 10321 16031 10379 16037
rect 10321 16028 10333 16031
rect 9916 16000 10333 16028
rect 9916 15988 9922 16000
rect 10321 15997 10333 16000
rect 10367 15997 10379 16031
rect 10321 15991 10379 15997
rect 10413 16031 10471 16037
rect 10413 15997 10425 16031
rect 10459 15997 10471 16031
rect 10413 15991 10471 15997
rect 10597 16031 10655 16037
rect 10597 15997 10609 16031
rect 10643 16028 10655 16031
rect 10778 16028 10784 16040
rect 10643 16000 10784 16028
rect 10643 15997 10655 16000
rect 10597 15991 10655 15997
rect 10428 15960 10456 15991
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 12529 16031 12587 16037
rect 12529 15997 12541 16031
rect 12575 15997 12587 16031
rect 12529 15991 12587 15997
rect 14185 16031 14243 16037
rect 14185 15997 14197 16031
rect 14231 16028 14243 16031
rect 14550 16028 14556 16040
rect 14231 16000 14556 16028
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 12434 15960 12440 15972
rect 8036 15932 8524 15960
rect 10152 15932 10456 15960
rect 12395 15932 12440 15960
rect 8036 15904 8064 15932
rect 10152 15904 10180 15932
rect 12434 15920 12440 15932
rect 12492 15920 12498 15972
rect 3878 15852 3884 15904
rect 3936 15892 3942 15904
rect 4065 15895 4123 15901
rect 4065 15892 4077 15895
rect 3936 15864 4077 15892
rect 3936 15852 3942 15864
rect 4065 15861 4077 15864
rect 4111 15861 4123 15895
rect 4065 15855 4123 15861
rect 7558 15852 7564 15904
rect 7616 15892 7622 15904
rect 7837 15895 7895 15901
rect 7837 15892 7849 15895
rect 7616 15864 7849 15892
rect 7616 15852 7622 15864
rect 7837 15861 7849 15864
rect 7883 15892 7895 15895
rect 8018 15892 8024 15904
rect 7883 15864 8024 15892
rect 7883 15861 7895 15864
rect 7837 15855 7895 15861
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 10134 15892 10140 15904
rect 10095 15864 10140 15892
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 12253 15895 12311 15901
rect 12253 15861 12265 15895
rect 12299 15892 12311 15895
rect 12544 15892 12572 15991
rect 14550 15988 14556 16000
rect 14608 15988 14614 16040
rect 14826 16028 14832 16040
rect 14787 16000 14832 16028
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 15838 16028 15844 16040
rect 15799 16000 15844 16028
rect 15838 15988 15844 16000
rect 15896 15988 15902 16040
rect 15010 15960 15016 15972
rect 14971 15932 15016 15960
rect 15010 15920 15016 15932
rect 15068 15920 15074 15972
rect 16206 15969 16212 15972
rect 16162 15963 16212 15969
rect 16162 15960 16174 15963
rect 15672 15932 16174 15960
rect 12894 15892 12900 15904
rect 12299 15864 12900 15892
rect 12299 15861 12311 15864
rect 12253 15855 12311 15861
rect 12894 15852 12900 15864
rect 12952 15852 12958 15904
rect 15470 15852 15476 15904
rect 15528 15892 15534 15904
rect 15672 15901 15700 15932
rect 16162 15929 16174 15932
rect 16208 15929 16212 15963
rect 16162 15923 16212 15929
rect 16206 15920 16212 15923
rect 16264 15960 16270 15972
rect 17037 15963 17095 15969
rect 17037 15960 17049 15963
rect 16264 15932 17049 15960
rect 16264 15920 16270 15932
rect 17037 15929 17049 15932
rect 17083 15929 17095 15963
rect 17037 15923 17095 15929
rect 18322 15920 18328 15972
rect 18380 15960 18386 15972
rect 18380 15932 18425 15960
rect 18380 15920 18386 15932
rect 19610 15920 19616 15972
rect 19668 15960 19674 15972
rect 19797 15963 19855 15969
rect 19797 15960 19809 15963
rect 19668 15932 19809 15960
rect 19668 15920 19674 15932
rect 19797 15929 19809 15932
rect 19843 15929 19855 15963
rect 19797 15923 19855 15929
rect 19889 15963 19947 15969
rect 19889 15929 19901 15963
rect 19935 15929 19947 15963
rect 19889 15923 19947 15929
rect 15657 15895 15715 15901
rect 15657 15892 15669 15895
rect 15528 15864 15669 15892
rect 15528 15852 15534 15864
rect 15657 15861 15669 15864
rect 15703 15861 15715 15895
rect 15657 15855 15715 15861
rect 18874 15852 18880 15904
rect 18932 15892 18938 15904
rect 19521 15895 19579 15901
rect 19521 15892 19533 15895
rect 18932 15864 19533 15892
rect 18932 15852 18938 15864
rect 19521 15861 19533 15864
rect 19567 15892 19579 15895
rect 19904 15892 19932 15923
rect 20070 15920 20076 15972
rect 20128 15960 20134 15972
rect 21177 15963 21235 15969
rect 21177 15960 21189 15963
rect 20128 15932 21189 15960
rect 20128 15920 20134 15932
rect 21177 15929 21189 15932
rect 21223 15960 21235 15963
rect 21453 15963 21511 15969
rect 21453 15960 21465 15963
rect 21223 15932 21465 15960
rect 21223 15929 21235 15932
rect 21177 15923 21235 15929
rect 21453 15929 21465 15932
rect 21499 15929 21511 15963
rect 21453 15923 21511 15929
rect 19567 15864 19932 15892
rect 19567 15861 19579 15864
rect 19521 15855 19579 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 3142 15648 3148 15700
rect 3200 15688 3206 15700
rect 3421 15691 3479 15697
rect 3421 15688 3433 15691
rect 3200 15660 3433 15688
rect 3200 15648 3206 15660
rect 3421 15657 3433 15660
rect 3467 15657 3479 15691
rect 3421 15651 3479 15657
rect 3510 15648 3516 15700
rect 3568 15688 3574 15700
rect 6457 15691 6515 15697
rect 6457 15688 6469 15691
rect 3568 15660 6469 15688
rect 3568 15648 3574 15660
rect 6457 15657 6469 15660
rect 6503 15657 6515 15691
rect 6457 15651 6515 15657
rect 8570 15648 8576 15700
rect 8628 15688 8634 15700
rect 8665 15691 8723 15697
rect 8665 15688 8677 15691
rect 8628 15660 8677 15688
rect 8628 15648 8634 15660
rect 8665 15657 8677 15660
rect 8711 15688 8723 15691
rect 10137 15691 10195 15697
rect 10137 15688 10149 15691
rect 8711 15660 10149 15688
rect 8711 15657 8723 15660
rect 8665 15651 8723 15657
rect 10137 15657 10149 15660
rect 10183 15657 10195 15691
rect 11606 15688 11612 15700
rect 11567 15660 11612 15688
rect 10137 15651 10195 15657
rect 11606 15648 11612 15660
rect 11664 15648 11670 15700
rect 15010 15648 15016 15700
rect 15068 15688 15074 15700
rect 15657 15691 15715 15697
rect 15657 15688 15669 15691
rect 15068 15660 15669 15688
rect 15068 15648 15074 15660
rect 15657 15657 15669 15660
rect 15703 15657 15715 15691
rect 16206 15688 16212 15700
rect 16167 15660 16212 15688
rect 15657 15651 15715 15657
rect 1762 15620 1768 15632
rect 1723 15592 1768 15620
rect 1762 15580 1768 15592
rect 1820 15580 1826 15632
rect 1857 15623 1915 15629
rect 1857 15589 1869 15623
rect 1903 15620 1915 15623
rect 1946 15620 1952 15632
rect 1903 15592 1952 15620
rect 1903 15589 1915 15592
rect 1857 15583 1915 15589
rect 1946 15580 1952 15592
rect 2004 15580 2010 15632
rect 3881 15623 3939 15629
rect 3881 15589 3893 15623
rect 3927 15620 3939 15623
rect 3970 15620 3976 15632
rect 3927 15592 3976 15620
rect 3927 15589 3939 15592
rect 3881 15583 3939 15589
rect 3970 15580 3976 15592
rect 4028 15580 4034 15632
rect 4154 15580 4160 15632
rect 4212 15620 4218 15632
rect 4249 15623 4307 15629
rect 4249 15620 4261 15623
rect 4212 15592 4261 15620
rect 4212 15580 4218 15592
rect 4249 15589 4261 15592
rect 4295 15589 4307 15623
rect 4249 15583 4307 15589
rect 4338 15580 4344 15632
rect 4396 15620 4402 15632
rect 5813 15623 5871 15629
rect 5813 15620 5825 15623
rect 4396 15592 5825 15620
rect 4396 15580 4402 15592
rect 5813 15589 5825 15592
rect 5859 15589 5871 15623
rect 7926 15620 7932 15632
rect 5813 15583 5871 15589
rect 5920 15592 7932 15620
rect 4798 15512 4804 15564
rect 4856 15552 4862 15564
rect 5537 15555 5595 15561
rect 5537 15552 5549 15555
rect 4856 15524 5549 15552
rect 4856 15512 4862 15524
rect 5537 15521 5549 15524
rect 5583 15552 5595 15555
rect 5920 15552 5948 15592
rect 7926 15580 7932 15592
rect 7984 15580 7990 15632
rect 9858 15620 9864 15632
rect 9324 15592 9864 15620
rect 5583 15524 5948 15552
rect 5997 15555 6055 15561
rect 5583 15521 5595 15524
rect 5537 15515 5595 15521
rect 5997 15521 6009 15555
rect 6043 15521 6055 15555
rect 6270 15552 6276 15564
rect 6231 15524 6276 15552
rect 5997 15515 6055 15521
rect 2406 15444 2412 15496
rect 2464 15484 2470 15496
rect 4157 15487 4215 15493
rect 4157 15484 4169 15487
rect 2464 15456 4169 15484
rect 2464 15444 2470 15456
rect 4157 15453 4169 15456
rect 4203 15484 4215 15487
rect 4338 15484 4344 15496
rect 4203 15456 4344 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4338 15444 4344 15456
rect 4396 15444 4402 15496
rect 4433 15487 4491 15493
rect 4433 15453 4445 15487
rect 4479 15453 4491 15487
rect 4433 15447 4491 15453
rect 2314 15416 2320 15428
rect 2275 15388 2320 15416
rect 2314 15376 2320 15388
rect 2372 15376 2378 15428
rect 3142 15416 3148 15428
rect 3055 15388 3148 15416
rect 3142 15376 3148 15388
rect 3200 15416 3206 15428
rect 4246 15416 4252 15428
rect 3200 15388 4252 15416
rect 3200 15376 3206 15388
rect 4246 15376 4252 15388
rect 4304 15376 4310 15428
rect 1946 15308 1952 15360
rect 2004 15348 2010 15360
rect 2685 15351 2743 15357
rect 2685 15348 2697 15351
rect 2004 15320 2697 15348
rect 2004 15308 2010 15320
rect 2685 15317 2697 15320
rect 2731 15317 2743 15351
rect 2685 15311 2743 15317
rect 3878 15308 3884 15360
rect 3936 15348 3942 15360
rect 4448 15348 4476 15447
rect 4614 15444 4620 15496
rect 4672 15484 4678 15496
rect 5077 15487 5135 15493
rect 5077 15484 5089 15487
rect 4672 15456 5089 15484
rect 4672 15444 4678 15456
rect 5077 15453 5089 15456
rect 5123 15453 5135 15487
rect 6012 15484 6040 15515
rect 6270 15512 6276 15524
rect 6328 15552 6334 15564
rect 7377 15555 7435 15561
rect 7377 15552 7389 15555
rect 6328 15524 7389 15552
rect 6328 15512 6334 15524
rect 7377 15521 7389 15524
rect 7423 15521 7435 15555
rect 7650 15552 7656 15564
rect 7611 15524 7656 15552
rect 7377 15515 7435 15521
rect 6638 15484 6644 15496
rect 6012 15456 6644 15484
rect 5077 15447 5135 15453
rect 6638 15444 6644 15456
rect 6696 15444 6702 15496
rect 7392 15484 7420 15515
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 7561 15487 7619 15493
rect 7561 15484 7573 15487
rect 7392 15456 7573 15484
rect 7561 15453 7573 15456
rect 7607 15484 7619 15487
rect 7926 15484 7932 15496
rect 7607 15456 7932 15484
rect 7607 15453 7619 15456
rect 7561 15447 7619 15453
rect 7926 15444 7932 15456
rect 7984 15444 7990 15496
rect 6089 15419 6147 15425
rect 6089 15385 6101 15419
rect 6135 15416 6147 15419
rect 6270 15416 6276 15428
rect 6135 15388 6276 15416
rect 6135 15385 6147 15388
rect 6089 15379 6147 15385
rect 6270 15376 6276 15388
rect 6328 15376 6334 15428
rect 6656 15416 6684 15444
rect 8938 15416 8944 15428
rect 6656 15388 8944 15416
rect 8938 15376 8944 15388
rect 8996 15416 9002 15428
rect 9324 15425 9352 15592
rect 9858 15580 9864 15592
rect 9916 15580 9922 15632
rect 11974 15580 11980 15632
rect 12032 15620 12038 15632
rect 12069 15623 12127 15629
rect 12069 15620 12081 15623
rect 12032 15592 12081 15620
rect 12032 15580 12038 15592
rect 12069 15589 12081 15592
rect 12115 15620 12127 15623
rect 12434 15620 12440 15632
rect 12115 15592 12440 15620
rect 12115 15589 12127 15592
rect 12069 15583 12127 15589
rect 12434 15580 12440 15592
rect 12492 15580 12498 15632
rect 9674 15552 9680 15564
rect 9635 15524 9680 15552
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15552 10011 15555
rect 10778 15552 10784 15564
rect 9999 15524 10784 15552
rect 9999 15521 10011 15524
rect 9953 15515 10011 15521
rect 10778 15512 10784 15524
rect 10836 15512 10842 15564
rect 13538 15552 13544 15564
rect 13499 15524 13544 15552
rect 13538 15512 13544 15524
rect 13596 15512 13602 15564
rect 15672 15552 15700 15651
rect 16206 15648 16212 15660
rect 16264 15648 16270 15700
rect 17402 15580 17408 15632
rect 17460 15620 17466 15632
rect 18049 15623 18107 15629
rect 18049 15620 18061 15623
rect 17460 15592 18061 15620
rect 17460 15580 17466 15592
rect 18049 15589 18061 15592
rect 18095 15620 18107 15623
rect 18874 15620 18880 15632
rect 18095 15592 18880 15620
rect 18095 15589 18107 15592
rect 18049 15583 18107 15589
rect 18874 15580 18880 15592
rect 18932 15580 18938 15632
rect 15841 15555 15899 15561
rect 15841 15552 15853 15555
rect 15672 15524 15853 15552
rect 15841 15521 15853 15524
rect 15887 15521 15899 15555
rect 19426 15552 19432 15564
rect 19387 15524 19432 15552
rect 15841 15515 15899 15521
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 11790 15444 11796 15496
rect 11848 15484 11854 15496
rect 11977 15487 12035 15493
rect 11977 15484 11989 15487
rect 11848 15456 11989 15484
rect 11848 15444 11854 15456
rect 11977 15453 11989 15456
rect 12023 15453 12035 15487
rect 12342 15484 12348 15496
rect 12303 15456 12348 15484
rect 11977 15447 12035 15453
rect 12342 15444 12348 15456
rect 12400 15444 12406 15496
rect 12618 15444 12624 15496
rect 12676 15484 12682 15496
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 12676 15456 13461 15484
rect 12676 15444 12682 15456
rect 13449 15453 13461 15456
rect 13495 15453 13507 15487
rect 17954 15484 17960 15496
rect 17867 15456 17960 15484
rect 13449 15447 13507 15453
rect 17954 15444 17960 15456
rect 18012 15484 18018 15496
rect 20901 15487 20959 15493
rect 20901 15484 20913 15487
rect 18012 15456 20913 15484
rect 18012 15444 18018 15456
rect 20901 15453 20913 15456
rect 20947 15453 20959 15487
rect 20901 15447 20959 15453
rect 9309 15419 9367 15425
rect 9309 15416 9321 15419
rect 8996 15388 9321 15416
rect 8996 15376 9002 15388
rect 9309 15385 9321 15388
rect 9355 15385 9367 15419
rect 9766 15416 9772 15428
rect 9727 15388 9772 15416
rect 9309 15379 9367 15385
rect 9766 15376 9772 15388
rect 9824 15376 9830 15428
rect 18414 15416 18420 15428
rect 17880 15388 18420 15416
rect 17880 15360 17908 15388
rect 18414 15376 18420 15388
rect 18472 15416 18478 15428
rect 18509 15419 18567 15425
rect 18509 15416 18521 15419
rect 18472 15388 18521 15416
rect 18472 15376 18478 15388
rect 18509 15385 18521 15388
rect 18555 15385 18567 15419
rect 18509 15379 18567 15385
rect 3936 15320 4476 15348
rect 3936 15308 3942 15320
rect 5994 15308 6000 15360
rect 6052 15348 6058 15360
rect 7009 15351 7067 15357
rect 7009 15348 7021 15351
rect 6052 15320 7021 15348
rect 6052 15308 6058 15320
rect 7009 15317 7021 15320
rect 7055 15317 7067 15351
rect 7009 15311 7067 15317
rect 9033 15351 9091 15357
rect 9033 15317 9045 15351
rect 9079 15348 9091 15351
rect 9122 15348 9128 15360
rect 9079 15320 9128 15348
rect 9079 15317 9091 15320
rect 9033 15311 9091 15317
rect 9122 15308 9128 15320
rect 9180 15308 9186 15360
rect 10778 15348 10784 15360
rect 10739 15320 10784 15348
rect 10778 15308 10784 15320
rect 10836 15308 10842 15360
rect 11054 15348 11060 15360
rect 11015 15320 11060 15348
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 12894 15348 12900 15360
rect 12855 15320 12900 15348
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 13262 15348 13268 15360
rect 13223 15320 13268 15348
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 16761 15351 16819 15357
rect 16761 15317 16773 15351
rect 16807 15348 16819 15351
rect 17402 15348 17408 15360
rect 16807 15320 17408 15348
rect 16807 15317 16819 15320
rect 16761 15311 16819 15317
rect 17402 15308 17408 15320
rect 17460 15308 17466 15360
rect 17773 15351 17831 15357
rect 17773 15317 17785 15351
rect 17819 15348 17831 15351
rect 17862 15348 17868 15360
rect 17819 15320 17868 15348
rect 17819 15317 17831 15320
rect 17773 15311 17831 15317
rect 17862 15308 17868 15320
rect 17920 15308 17926 15360
rect 18138 15308 18144 15360
rect 18196 15348 18202 15360
rect 18969 15351 19027 15357
rect 18969 15348 18981 15351
rect 18196 15320 18981 15348
rect 18196 15308 18202 15320
rect 18969 15317 18981 15320
rect 19015 15348 19027 15351
rect 19567 15351 19625 15357
rect 19567 15348 19579 15351
rect 19015 15320 19579 15348
rect 19015 15317 19027 15320
rect 18969 15311 19027 15317
rect 19567 15317 19579 15320
rect 19613 15317 19625 15351
rect 19567 15311 19625 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2038 15104 2044 15156
rect 2096 15144 2102 15156
rect 6549 15147 6607 15153
rect 6549 15144 6561 15147
rect 2096 15116 6561 15144
rect 2096 15104 2102 15116
rect 6549 15113 6561 15116
rect 6595 15113 6607 15147
rect 6549 15107 6607 15113
rect 2685 15011 2743 15017
rect 2685 14977 2697 15011
rect 2731 15008 2743 15011
rect 3142 15008 3148 15020
rect 2731 14980 3148 15008
rect 2731 14977 2743 14980
rect 2685 14971 2743 14977
rect 3142 14968 3148 14980
rect 3200 14968 3206 15020
rect 4798 15008 4804 15020
rect 4540 14980 4804 15008
rect 3602 14900 3608 14952
rect 3660 14940 3666 14952
rect 4154 14940 4160 14952
rect 3660 14912 4160 14940
rect 3660 14900 3666 14912
rect 4154 14900 4160 14912
rect 4212 14940 4218 14952
rect 4540 14949 4568 14980
rect 4798 14968 4804 14980
rect 4856 14968 4862 15020
rect 4525 14943 4583 14949
rect 4525 14940 4537 14943
rect 4212 14912 4537 14940
rect 4212 14900 4218 14912
rect 4525 14909 4537 14912
rect 4571 14909 4583 14943
rect 4525 14903 4583 14909
rect 4614 14900 4620 14952
rect 4672 14940 4678 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4672 14912 4905 14940
rect 4672 14900 4678 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 5445 14943 5503 14949
rect 5445 14909 5457 14943
rect 5491 14940 5503 14943
rect 5534 14940 5540 14952
rect 5491 14912 5540 14940
rect 5491 14909 5503 14912
rect 5445 14903 5503 14909
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 5813 14943 5871 14949
rect 5813 14909 5825 14943
rect 5859 14940 5871 14943
rect 5994 14940 6000 14952
rect 5859 14912 6000 14940
rect 5859 14909 5871 14912
rect 5813 14903 5871 14909
rect 5994 14900 6000 14912
rect 6052 14900 6058 14952
rect 6564 14940 6592 15107
rect 10042 15104 10048 15156
rect 10100 15144 10106 15156
rect 10229 15147 10287 15153
rect 10229 15144 10241 15147
rect 10100 15116 10241 15144
rect 10100 15104 10106 15116
rect 10229 15113 10241 15116
rect 10275 15144 10287 15147
rect 10321 15147 10379 15153
rect 10321 15144 10333 15147
rect 10275 15116 10333 15144
rect 10275 15113 10287 15116
rect 10229 15107 10287 15113
rect 10321 15113 10333 15116
rect 10367 15113 10379 15147
rect 11974 15144 11980 15156
rect 11935 15116 11980 15144
rect 10321 15107 10379 15113
rect 11974 15104 11980 15116
rect 12032 15104 12038 15156
rect 17402 15144 17408 15156
rect 17363 15116 17408 15144
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 17865 15147 17923 15153
rect 17865 15113 17877 15147
rect 17911 15144 17923 15147
rect 17954 15144 17960 15156
rect 17911 15116 17960 15144
rect 17911 15113 17923 15116
rect 17865 15107 17923 15113
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 12342 15036 12348 15088
rect 12400 15076 12406 15088
rect 13081 15079 13139 15085
rect 13081 15076 13093 15079
rect 12400 15048 13093 15076
rect 12400 15036 12406 15048
rect 13081 15045 13093 15048
rect 13127 15045 13139 15079
rect 13081 15039 13139 15045
rect 17770 15036 17776 15088
rect 17828 15076 17834 15088
rect 21361 15079 21419 15085
rect 21361 15076 21373 15079
rect 17828 15048 21373 15076
rect 17828 15036 17834 15048
rect 21361 15045 21373 15048
rect 21407 15045 21419 15079
rect 21361 15039 21419 15045
rect 9398 14968 9404 15020
rect 9456 15008 9462 15020
rect 10505 15011 10563 15017
rect 10505 15008 10517 15011
rect 9456 14980 10517 15008
rect 9456 14968 9462 14980
rect 10505 14977 10517 14980
rect 10551 15008 10563 15011
rect 11054 15008 11060 15020
rect 10551 14980 11060 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 12529 15011 12587 15017
rect 12529 14977 12541 15011
rect 12575 15008 12587 15011
rect 13262 15008 13268 15020
rect 12575 14980 13268 15008
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 18138 15008 18144 15020
rect 18099 14980 18144 15008
rect 18138 14968 18144 14980
rect 18196 14968 18202 15020
rect 18414 15008 18420 15020
rect 18375 14980 18420 15008
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 19153 15011 19211 15017
rect 19153 14977 19165 15011
rect 19199 15008 19211 15011
rect 19794 15008 19800 15020
rect 19199 14980 19800 15008
rect 19199 14977 19211 14980
rect 19153 14971 19211 14977
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6564 14912 6837 14940
rect 6825 14909 6837 14912
rect 6871 14940 6883 14943
rect 7561 14943 7619 14949
rect 7561 14940 7573 14943
rect 6871 14912 7573 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 7561 14909 7573 14912
rect 7607 14940 7619 14943
rect 7650 14940 7656 14952
rect 7607 14912 7656 14940
rect 7607 14909 7619 14912
rect 7561 14903 7619 14909
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 7926 14940 7932 14952
rect 7887 14912 7932 14940
rect 7926 14900 7932 14912
rect 7984 14900 7990 14952
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 8389 14943 8447 14949
rect 8389 14940 8401 14943
rect 8352 14912 8401 14940
rect 8352 14900 8358 14912
rect 8389 14909 8401 14912
rect 8435 14909 8447 14943
rect 8754 14940 8760 14952
rect 8715 14912 8760 14940
rect 8389 14903 8447 14909
rect 3006 14875 3064 14881
rect 3006 14872 3018 14875
rect 2608 14844 3018 14872
rect 2608 14816 2636 14844
rect 3006 14841 3018 14844
rect 3052 14872 3064 14875
rect 3418 14872 3424 14884
rect 3052 14844 3424 14872
rect 3052 14841 3064 14844
rect 3006 14835 3064 14841
rect 3418 14832 3424 14844
rect 3476 14832 3482 14884
rect 5350 14832 5356 14884
rect 5408 14872 5414 14884
rect 5408 14844 7052 14872
rect 5408 14832 5414 14844
rect 7024 14816 7052 14844
rect 1394 14804 1400 14816
rect 1355 14776 1400 14804
rect 1394 14764 1400 14776
rect 1452 14764 1458 14816
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 2590 14804 2596 14816
rect 2551 14776 2596 14804
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 3602 14804 3608 14816
rect 3563 14776 3608 14804
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 4062 14804 4068 14816
rect 4023 14776 4068 14804
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 4522 14804 4528 14816
rect 4483 14776 4528 14804
rect 4522 14764 4528 14776
rect 4580 14764 4586 14816
rect 6270 14804 6276 14816
rect 6231 14776 6276 14804
rect 6270 14764 6276 14776
rect 6328 14764 6334 14816
rect 7006 14804 7012 14816
rect 6919 14776 7012 14804
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 8404 14804 8432 14903
rect 8754 14900 8760 14912
rect 8812 14900 8818 14952
rect 9122 14940 9128 14952
rect 9083 14912 9128 14940
rect 9122 14900 9128 14912
rect 9180 14900 9186 14952
rect 14461 14943 14519 14949
rect 14461 14940 14473 14943
rect 14292 14912 14473 14940
rect 9401 14875 9459 14881
rect 9401 14841 9413 14875
rect 9447 14872 9459 14875
rect 10686 14872 10692 14884
rect 9447 14844 10692 14872
rect 9447 14841 9459 14844
rect 9401 14835 9459 14841
rect 10686 14832 10692 14844
rect 10744 14832 10750 14884
rect 12621 14875 12679 14881
rect 12621 14841 12633 14875
rect 12667 14872 12679 14875
rect 12894 14872 12900 14884
rect 12667 14844 12900 14872
rect 12667 14841 12679 14844
rect 12621 14835 12679 14841
rect 9677 14807 9735 14813
rect 9677 14804 9689 14807
rect 8404 14776 9689 14804
rect 9677 14773 9689 14776
rect 9723 14804 9735 14807
rect 9766 14804 9772 14816
rect 9723 14776 9772 14804
rect 9723 14773 9735 14776
rect 9677 14767 9735 14773
rect 9766 14764 9772 14776
rect 9824 14764 9830 14816
rect 10229 14807 10287 14813
rect 10229 14773 10241 14807
rect 10275 14804 10287 14807
rect 10870 14804 10876 14816
rect 10275 14776 10876 14804
rect 10275 14773 10287 14776
rect 10229 14767 10287 14773
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 11425 14807 11483 14813
rect 11425 14773 11437 14807
rect 11471 14804 11483 14807
rect 12636 14804 12664 14835
rect 12894 14832 12900 14844
rect 12952 14832 12958 14884
rect 14292 14816 14320 14912
rect 14461 14909 14473 14912
rect 14507 14909 14519 14943
rect 14461 14903 14519 14909
rect 14826 14900 14832 14952
rect 14884 14940 14890 14952
rect 14921 14943 14979 14949
rect 14921 14940 14933 14943
rect 14884 14912 14933 14940
rect 14884 14900 14890 14912
rect 14921 14909 14933 14912
rect 14967 14909 14979 14943
rect 14921 14903 14979 14909
rect 15197 14943 15255 14949
rect 15197 14909 15209 14943
rect 15243 14940 15255 14943
rect 16025 14943 16083 14949
rect 16025 14940 16037 14943
rect 15243 14912 16037 14940
rect 15243 14909 15255 14912
rect 15197 14903 15255 14909
rect 16025 14909 16037 14912
rect 16071 14940 16083 14943
rect 16482 14940 16488 14952
rect 16071 14912 16488 14940
rect 16071 14909 16083 14912
rect 16025 14903 16083 14909
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 16945 14943 17003 14949
rect 16945 14909 16957 14943
rect 16991 14909 17003 14943
rect 16945 14903 17003 14909
rect 16346 14875 16404 14881
rect 16346 14841 16358 14875
rect 16392 14841 16404 14875
rect 16960 14872 16988 14903
rect 18138 14872 18144 14884
rect 16960 14844 18144 14872
rect 16346 14835 16404 14841
rect 13538 14804 13544 14816
rect 11471 14776 12664 14804
rect 13499 14776 13544 14804
rect 11471 14773 11483 14776
rect 11425 14767 11483 14773
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 14274 14804 14280 14816
rect 14235 14776 14280 14804
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 15470 14804 15476 14816
rect 15431 14776 15476 14804
rect 15470 14764 15476 14776
rect 15528 14804 15534 14816
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 15528 14776 15853 14804
rect 15528 14764 15534 14776
rect 15841 14773 15853 14776
rect 15887 14804 15899 14807
rect 16361 14804 16389 14835
rect 18138 14832 18144 14844
rect 18196 14872 18202 14884
rect 18233 14875 18291 14881
rect 18233 14872 18245 14875
rect 18196 14844 18245 14872
rect 18196 14832 18202 14844
rect 18233 14841 18245 14844
rect 18279 14841 18291 14875
rect 18233 14835 18291 14841
rect 18322 14832 18328 14884
rect 18380 14872 18386 14884
rect 19168 14872 19196 14971
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 19978 15008 19984 15020
rect 19939 14980 19984 15008
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 21174 14940 21180 14952
rect 21135 14912 21180 14940
rect 21174 14900 21180 14912
rect 21232 14940 21238 14952
rect 21637 14943 21695 14949
rect 21637 14940 21649 14943
rect 21232 14912 21649 14940
rect 21232 14900 21238 14912
rect 21637 14909 21649 14912
rect 21683 14909 21695 14943
rect 21637 14903 21695 14909
rect 18380 14844 19196 14872
rect 18380 14832 18386 14844
rect 19518 14832 19524 14884
rect 19576 14872 19582 14884
rect 19705 14875 19763 14881
rect 19705 14872 19717 14875
rect 19576 14844 19717 14872
rect 19576 14832 19582 14844
rect 19705 14841 19717 14844
rect 19751 14841 19763 14875
rect 19705 14835 19763 14841
rect 19794 14832 19800 14884
rect 19852 14872 19858 14884
rect 19852 14844 19897 14872
rect 19852 14832 19858 14844
rect 19426 14804 19432 14816
rect 15887 14776 16389 14804
rect 19339 14776 19432 14804
rect 15887 14773 15899 14776
rect 15841 14767 15899 14773
rect 19426 14764 19432 14776
rect 19484 14804 19490 14816
rect 20254 14804 20260 14816
rect 19484 14776 20260 14804
rect 19484 14764 19490 14776
rect 20254 14764 20260 14776
rect 20312 14764 20318 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 2409 14603 2467 14609
rect 2409 14600 2421 14603
rect 2004 14572 2421 14600
rect 2004 14560 2010 14572
rect 2409 14569 2421 14572
rect 2455 14569 2467 14603
rect 2409 14563 2467 14569
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14600 3295 14603
rect 3602 14600 3608 14612
rect 3283 14572 3608 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 3602 14560 3608 14572
rect 3660 14560 3666 14612
rect 4246 14560 4252 14612
rect 4304 14600 4310 14612
rect 4709 14603 4767 14609
rect 4709 14600 4721 14603
rect 4304 14572 4721 14600
rect 4304 14560 4310 14572
rect 4709 14569 4721 14572
rect 4755 14569 4767 14603
rect 6178 14600 6184 14612
rect 6139 14572 6184 14600
rect 4709 14563 4767 14569
rect 6178 14560 6184 14572
rect 6236 14560 6242 14612
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 9732 14572 10149 14600
rect 9732 14560 9738 14572
rect 10137 14569 10149 14572
rect 10183 14569 10195 14603
rect 11790 14600 11796 14612
rect 10137 14563 10195 14569
rect 10565 14572 11796 14600
rect 1851 14535 1909 14541
rect 1851 14501 1863 14535
rect 1897 14532 1909 14535
rect 2590 14532 2596 14544
rect 1897 14504 2596 14532
rect 1897 14501 1909 14504
rect 1851 14495 1909 14501
rect 2590 14492 2596 14504
rect 2648 14492 2654 14544
rect 2777 14535 2835 14541
rect 2777 14501 2789 14535
rect 2823 14532 2835 14535
rect 4522 14532 4528 14544
rect 2823 14504 4528 14532
rect 2823 14501 2835 14504
rect 2777 14495 2835 14501
rect 1489 14467 1547 14473
rect 1489 14433 1501 14467
rect 1535 14464 1547 14467
rect 2792 14464 2820 14495
rect 4522 14492 4528 14504
rect 4580 14492 4586 14544
rect 8573 14535 8631 14541
rect 8573 14501 8585 14535
rect 8619 14532 8631 14535
rect 10565 14532 10593 14572
rect 11790 14560 11796 14572
rect 11848 14600 11854 14612
rect 11885 14603 11943 14609
rect 11885 14600 11897 14603
rect 11848 14572 11897 14600
rect 11848 14560 11854 14572
rect 11885 14569 11897 14572
rect 11931 14569 11943 14603
rect 11885 14563 11943 14569
rect 14553 14603 14611 14609
rect 14553 14569 14565 14603
rect 14599 14600 14611 14603
rect 14826 14600 14832 14612
rect 14599 14572 14832 14600
rect 14599 14569 14611 14572
rect 14553 14563 14611 14569
rect 14826 14560 14832 14572
rect 14884 14560 14890 14612
rect 16482 14600 16488 14612
rect 16443 14572 16488 14600
rect 16482 14560 16488 14572
rect 16540 14560 16546 14612
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 18233 14603 18291 14609
rect 18233 14600 18245 14603
rect 18196 14572 18245 14600
rect 18196 14560 18202 14572
rect 18233 14569 18245 14572
rect 18279 14600 18291 14603
rect 18414 14600 18420 14612
rect 18279 14572 18420 14600
rect 18279 14569 18291 14572
rect 18233 14563 18291 14569
rect 18414 14560 18420 14572
rect 18472 14600 18478 14612
rect 20070 14600 20076 14612
rect 18472 14572 20076 14600
rect 18472 14560 18478 14572
rect 20070 14560 20076 14572
rect 20128 14560 20134 14612
rect 8619 14504 10593 14532
rect 8619 14501 8631 14504
rect 8573 14495 8631 14501
rect 10870 14492 10876 14544
rect 10928 14532 10934 14544
rect 11010 14535 11068 14541
rect 11010 14532 11022 14535
rect 10928 14504 11022 14532
rect 10928 14492 10934 14504
rect 11010 14501 11022 14504
rect 11056 14501 11068 14535
rect 11010 14495 11068 14501
rect 12250 14492 12256 14544
rect 12308 14532 12314 14544
rect 12618 14532 12624 14544
rect 12308 14504 12624 14532
rect 12308 14492 12314 14504
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 13173 14535 13231 14541
rect 13173 14501 13185 14535
rect 13219 14532 13231 14535
rect 13262 14532 13268 14544
rect 13219 14504 13268 14532
rect 13219 14501 13231 14504
rect 13173 14495 13231 14501
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 15470 14492 15476 14544
rect 15528 14532 15534 14544
rect 15610 14535 15668 14541
rect 15610 14532 15622 14535
rect 15528 14504 15622 14532
rect 15528 14492 15534 14504
rect 15610 14501 15622 14504
rect 15656 14501 15668 14535
rect 17218 14532 17224 14544
rect 17179 14504 17224 14532
rect 15610 14495 15668 14501
rect 17218 14492 17224 14504
rect 17276 14492 17282 14544
rect 17313 14535 17371 14541
rect 17313 14501 17325 14535
rect 17359 14532 17371 14535
rect 17402 14532 17408 14544
rect 17359 14504 17408 14532
rect 17359 14501 17371 14504
rect 17313 14495 17371 14501
rect 17402 14492 17408 14504
rect 17460 14492 17466 14544
rect 17862 14532 17868 14544
rect 17823 14504 17868 14532
rect 17862 14492 17868 14504
rect 17920 14492 17926 14544
rect 18046 14492 18052 14544
rect 18104 14532 18110 14544
rect 18785 14535 18843 14541
rect 18785 14532 18797 14535
rect 18104 14504 18797 14532
rect 18104 14492 18110 14504
rect 18785 14501 18797 14504
rect 18831 14501 18843 14535
rect 18785 14495 18843 14501
rect 18874 14492 18880 14544
rect 18932 14532 18938 14544
rect 18932 14504 18977 14532
rect 18932 14492 18938 14504
rect 19242 14492 19248 14544
rect 19300 14532 19306 14544
rect 19978 14532 19984 14544
rect 19300 14504 19984 14532
rect 19300 14492 19306 14504
rect 19978 14492 19984 14504
rect 20036 14492 20042 14544
rect 1535 14436 2820 14464
rect 1535 14433 1547 14436
rect 1489 14427 1547 14433
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 4212 14436 4445 14464
rect 4212 14424 4218 14436
rect 4433 14433 4445 14436
rect 4479 14433 4491 14467
rect 4433 14427 4491 14433
rect 4614 14424 4620 14476
rect 4672 14464 4678 14476
rect 4893 14467 4951 14473
rect 4893 14464 4905 14467
rect 4672 14436 4905 14464
rect 4672 14424 4678 14436
rect 4893 14433 4905 14436
rect 4939 14433 4951 14467
rect 4893 14427 4951 14433
rect 5445 14467 5503 14473
rect 5445 14433 5457 14467
rect 5491 14464 5503 14467
rect 5534 14464 5540 14476
rect 5491 14436 5540 14464
rect 5491 14433 5503 14436
rect 5445 14427 5503 14433
rect 4341 14399 4399 14405
rect 4341 14396 4353 14399
rect 4126 14368 4353 14396
rect 3142 14288 3148 14340
rect 3200 14328 3206 14340
rect 3786 14328 3792 14340
rect 3200 14300 3792 14328
rect 3200 14288 3206 14300
rect 3786 14288 3792 14300
rect 3844 14328 3850 14340
rect 4126 14328 4154 14368
rect 4341 14365 4353 14368
rect 4387 14396 4399 14399
rect 5460 14396 5488 14427
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 5813 14467 5871 14473
rect 5813 14433 5825 14467
rect 5859 14464 5871 14467
rect 5994 14464 6000 14476
rect 5859 14436 6000 14464
rect 5859 14433 5871 14436
rect 5813 14427 5871 14433
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6822 14464 6828 14476
rect 6783 14436 6828 14464
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 9582 14464 9588 14476
rect 9171 14436 9588 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 9582 14424 9588 14436
rect 9640 14464 9646 14476
rect 9712 14467 9770 14473
rect 9712 14464 9724 14467
rect 9640 14436 9724 14464
rect 9640 14424 9646 14436
rect 9712 14433 9724 14436
rect 9758 14433 9770 14467
rect 9712 14427 9770 14433
rect 9815 14467 9873 14473
rect 9815 14433 9827 14467
rect 9861 14464 9873 14467
rect 11790 14464 11796 14476
rect 9861 14436 11796 14464
rect 9861 14433 9873 14436
rect 9815 14427 9873 14433
rect 11790 14424 11796 14436
rect 11848 14424 11854 14476
rect 13998 14464 14004 14476
rect 13962 14436 14004 14464
rect 13998 14424 14004 14436
rect 14056 14473 14062 14476
rect 14056 14467 14110 14473
rect 14056 14433 14064 14467
rect 14098 14464 14110 14467
rect 14734 14464 14740 14476
rect 14098 14436 14740 14464
rect 14098 14433 14110 14436
rect 14056 14427 14110 14433
rect 14056 14424 14062 14427
rect 14734 14424 14740 14436
rect 14792 14424 14798 14476
rect 20806 14464 20812 14476
rect 20767 14436 20812 14464
rect 20806 14424 20812 14436
rect 20864 14464 20870 14476
rect 24581 14467 24639 14473
rect 24581 14464 24593 14467
rect 20864 14436 24593 14464
rect 20864 14424 20870 14436
rect 24581 14433 24593 14436
rect 24627 14464 24639 14467
rect 25038 14464 25044 14476
rect 24627 14436 25044 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 25038 14424 25044 14436
rect 25096 14424 25102 14476
rect 4387 14368 5488 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 6270 14356 6276 14408
rect 6328 14396 6334 14408
rect 6733 14399 6791 14405
rect 6733 14396 6745 14399
rect 6328 14368 6745 14396
rect 6328 14356 6334 14368
rect 6733 14365 6745 14368
rect 6779 14365 6791 14399
rect 6733 14359 6791 14365
rect 7926 14356 7932 14408
rect 7984 14396 7990 14408
rect 8297 14399 8355 14405
rect 8297 14396 8309 14399
rect 7984 14368 8309 14396
rect 7984 14356 7990 14368
rect 8297 14365 8309 14368
rect 8343 14396 8355 14399
rect 8754 14396 8760 14408
rect 8343 14368 8760 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 10686 14396 10692 14408
rect 10647 14368 10692 14396
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 12529 14399 12587 14405
rect 12529 14365 12541 14399
rect 12575 14396 12587 14399
rect 13449 14399 13507 14405
rect 13449 14396 13461 14399
rect 12575 14368 13461 14396
rect 12575 14365 12587 14368
rect 12529 14359 12587 14365
rect 13449 14365 13461 14368
rect 13495 14396 13507 14399
rect 14139 14399 14197 14405
rect 14139 14396 14151 14399
rect 13495 14368 14151 14396
rect 13495 14365 13507 14368
rect 13449 14359 13507 14365
rect 14139 14365 14151 14368
rect 14185 14365 14197 14399
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 14139 14359 14197 14365
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 18138 14356 18144 14408
rect 18196 14396 18202 14408
rect 18509 14399 18567 14405
rect 18509 14396 18521 14399
rect 18196 14368 18521 14396
rect 18196 14356 18202 14368
rect 18509 14365 18521 14368
rect 18555 14365 18567 14399
rect 18509 14359 18567 14365
rect 19061 14399 19119 14405
rect 19061 14365 19073 14399
rect 19107 14365 19119 14399
rect 19061 14359 19119 14365
rect 3844 14300 4154 14328
rect 3844 14288 3850 14300
rect 4246 14288 4252 14340
rect 4304 14328 4310 14340
rect 5074 14328 5080 14340
rect 4304 14300 5080 14328
rect 4304 14288 4310 14300
rect 5074 14288 5080 14300
rect 5132 14288 5138 14340
rect 11609 14331 11667 14337
rect 11609 14297 11621 14331
rect 11655 14328 11667 14331
rect 12618 14328 12624 14340
rect 11655 14300 12624 14328
rect 11655 14297 11667 14300
rect 11609 14291 11667 14297
rect 12618 14288 12624 14300
rect 12676 14288 12682 14340
rect 18230 14288 18236 14340
rect 18288 14328 18294 14340
rect 19076 14328 19104 14359
rect 19242 14328 19248 14340
rect 18288 14300 19248 14328
rect 18288 14288 18294 14300
rect 19242 14288 19248 14300
rect 19300 14288 19306 14340
rect 24762 14328 24768 14340
rect 24723 14300 24768 14328
rect 24762 14288 24768 14300
rect 24820 14288 24826 14340
rect 3881 14263 3939 14269
rect 3881 14229 3893 14263
rect 3927 14260 3939 14263
rect 6086 14260 6092 14272
rect 3927 14232 6092 14260
rect 3927 14229 3939 14232
rect 3881 14223 3939 14229
rect 6086 14220 6092 14232
rect 6144 14220 6150 14272
rect 6638 14260 6644 14272
rect 6599 14232 6644 14260
rect 6638 14220 6644 14232
rect 6696 14220 6702 14272
rect 7466 14220 7472 14272
rect 7524 14260 7530 14272
rect 7929 14263 7987 14269
rect 7929 14260 7941 14263
rect 7524 14232 7941 14260
rect 7524 14220 7530 14232
rect 7929 14229 7941 14232
rect 7975 14260 7987 14263
rect 8294 14260 8300 14272
rect 7975 14232 8300 14260
rect 7975 14229 7987 14232
rect 7929 14223 7987 14229
rect 8294 14220 8300 14232
rect 8352 14220 8358 14272
rect 9306 14220 9312 14272
rect 9364 14260 9370 14272
rect 9401 14263 9459 14269
rect 9401 14260 9413 14263
rect 9364 14232 9413 14260
rect 9364 14220 9370 14232
rect 9401 14229 9413 14232
rect 9447 14260 9459 14263
rect 10502 14260 10508 14272
rect 9447 14232 10508 14260
rect 9447 14229 9459 14232
rect 9401 14223 9459 14229
rect 10502 14220 10508 14232
rect 10560 14260 10566 14272
rect 10778 14260 10784 14272
rect 10560 14232 10784 14260
rect 10560 14220 10566 14232
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 12345 14263 12403 14269
rect 12345 14229 12357 14263
rect 12391 14260 12403 14263
rect 12526 14260 12532 14272
rect 12391 14232 12532 14260
rect 12391 14229 12403 14232
rect 12345 14223 12403 14229
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 16209 14263 16267 14269
rect 16209 14229 16221 14263
rect 16255 14260 16267 14263
rect 17402 14260 17408 14272
rect 16255 14232 17408 14260
rect 16255 14229 16267 14232
rect 16209 14223 16267 14229
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 19518 14220 19524 14272
rect 19576 14260 19582 14272
rect 19794 14260 19800 14272
rect 19576 14232 19800 14260
rect 19576 14220 19582 14232
rect 19794 14220 19800 14232
rect 19852 14220 19858 14272
rect 20162 14220 20168 14272
rect 20220 14260 20226 14272
rect 21039 14263 21097 14269
rect 21039 14260 21051 14263
rect 20220 14232 21051 14260
rect 20220 14220 20226 14232
rect 21039 14229 21051 14232
rect 21085 14229 21097 14263
rect 21039 14223 21097 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1946 14016 1952 14068
rect 2004 14056 2010 14068
rect 2222 14056 2228 14068
rect 2004 14028 2228 14056
rect 2004 14016 2010 14028
rect 2222 14016 2228 14028
rect 2280 14056 2286 14068
rect 2961 14059 3019 14065
rect 2961 14056 2973 14059
rect 2280 14028 2973 14056
rect 2280 14016 2286 14028
rect 2961 14025 2973 14028
rect 3007 14025 3019 14059
rect 2961 14019 3019 14025
rect 3786 14016 3792 14068
rect 3844 14056 3850 14068
rect 3970 14056 3976 14068
rect 3844 14028 3976 14056
rect 3844 14016 3850 14028
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 4525 14059 4583 14065
rect 4525 14025 4537 14059
rect 4571 14056 4583 14059
rect 4614 14056 4620 14068
rect 4571 14028 4620 14056
rect 4571 14025 4583 14028
rect 4525 14019 4583 14025
rect 4614 14016 4620 14028
rect 4672 14056 4678 14068
rect 4893 14059 4951 14065
rect 4893 14056 4905 14059
rect 4672 14028 4905 14056
rect 4672 14016 4678 14028
rect 4893 14025 4905 14028
rect 4939 14025 4951 14059
rect 6270 14056 6276 14068
rect 6231 14028 6276 14056
rect 4893 14019 4951 14025
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 1854 13920 1860 13932
rect 1719 13892 1860 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 1854 13880 1860 13892
rect 1912 13920 1918 13932
rect 3050 13920 3056 13932
rect 1912 13892 3056 13920
rect 1912 13880 1918 13892
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 4908 13920 4936 14019
rect 6270 14016 6276 14028
rect 6328 14016 6334 14068
rect 8754 14016 8760 14068
rect 8812 14056 8818 14068
rect 9674 14056 9680 14068
rect 8812 14028 9680 14056
rect 8812 14016 8818 14028
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 10686 14016 10692 14068
rect 10744 14056 10750 14068
rect 11609 14059 11667 14065
rect 11609 14056 11621 14059
rect 10744 14028 11621 14056
rect 10744 14016 10750 14028
rect 11609 14025 11621 14028
rect 11655 14025 11667 14059
rect 12250 14056 12256 14068
rect 12211 14028 12256 14056
rect 11609 14019 11667 14025
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 13725 14059 13783 14065
rect 13725 14025 13737 14059
rect 13771 14056 13783 14059
rect 14826 14056 14832 14068
rect 13771 14028 14832 14056
rect 13771 14025 13783 14028
rect 13725 14019 13783 14025
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 17221 14059 17279 14065
rect 17221 14025 17233 14059
rect 17267 14056 17279 14059
rect 17402 14056 17408 14068
rect 17267 14028 17408 14056
rect 17267 14025 17279 14028
rect 17221 14019 17279 14025
rect 17402 14016 17408 14028
rect 17460 14056 17466 14068
rect 17865 14059 17923 14065
rect 17865 14056 17877 14059
rect 17460 14028 17877 14056
rect 17460 14016 17466 14028
rect 17865 14025 17877 14028
rect 17911 14056 17923 14059
rect 18322 14056 18328 14068
rect 17911 14028 18328 14056
rect 17911 14025 17923 14028
rect 17865 14019 17923 14025
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 18874 14016 18880 14068
rect 18932 14056 18938 14068
rect 19061 14059 19119 14065
rect 19061 14056 19073 14059
rect 18932 14028 19073 14056
rect 18932 14016 18938 14028
rect 19061 14025 19073 14028
rect 19107 14025 19119 14059
rect 19061 14019 19119 14025
rect 19794 14016 19800 14068
rect 19852 14056 19858 14068
rect 24719 14059 24777 14065
rect 24719 14056 24731 14059
rect 19852 14028 24731 14056
rect 19852 14016 19858 14028
rect 24719 14025 24731 14028
rect 24765 14025 24777 14059
rect 25038 14056 25044 14068
rect 24999 14028 25044 14056
rect 24719 14019 24777 14025
rect 25038 14016 25044 14028
rect 25096 14016 25102 14068
rect 5074 13948 5080 14000
rect 5132 13988 5138 14000
rect 5994 13988 6000 14000
rect 5132 13960 6000 13988
rect 5132 13948 5138 13960
rect 5994 13948 6000 13960
rect 6052 13988 6058 14000
rect 6641 13991 6699 13997
rect 6641 13988 6653 13991
rect 6052 13960 6653 13988
rect 6052 13948 6058 13960
rect 6641 13957 6653 13960
rect 6687 13988 6699 13991
rect 8938 13988 8944 14000
rect 6687 13960 8944 13988
rect 6687 13957 6699 13960
rect 6641 13951 6699 13957
rect 8938 13948 8944 13960
rect 8996 13948 9002 14000
rect 4908 13892 6776 13920
rect 3970 13812 3976 13864
rect 4028 13852 4034 13864
rect 4709 13855 4767 13861
rect 4709 13852 4721 13855
rect 4028 13824 4721 13852
rect 4028 13812 4034 13824
rect 4709 13821 4721 13824
rect 4755 13821 4767 13855
rect 5534 13852 5540 13864
rect 5495 13824 5540 13852
rect 4709 13815 4767 13821
rect 1670 13744 1676 13796
rect 1728 13784 1734 13796
rect 1765 13787 1823 13793
rect 1765 13784 1777 13787
rect 1728 13756 1777 13784
rect 1728 13744 1734 13756
rect 1765 13753 1777 13756
rect 1811 13784 1823 13787
rect 1946 13784 1952 13796
rect 1811 13756 1952 13784
rect 1811 13753 1823 13756
rect 1765 13747 1823 13753
rect 1946 13744 1952 13756
rect 2004 13744 2010 13796
rect 2314 13784 2320 13796
rect 2227 13756 2320 13784
rect 2314 13744 2320 13756
rect 2372 13784 2378 13796
rect 3237 13787 3295 13793
rect 3237 13784 3249 13787
rect 2372 13756 3249 13784
rect 2372 13744 2378 13756
rect 3237 13753 3249 13756
rect 3283 13753 3295 13787
rect 3237 13747 3295 13753
rect 3329 13787 3387 13793
rect 3329 13753 3341 13787
rect 3375 13784 3387 13787
rect 3510 13784 3516 13796
rect 3375 13756 3516 13784
rect 3375 13753 3387 13756
rect 3329 13747 3387 13753
rect 2590 13716 2596 13728
rect 2551 13688 2596 13716
rect 2590 13676 2596 13688
rect 2648 13676 2654 13728
rect 3252 13716 3280 13747
rect 3510 13744 3516 13756
rect 3568 13744 3574 13796
rect 3878 13784 3884 13796
rect 3839 13756 3884 13784
rect 3878 13744 3884 13756
rect 3936 13744 3942 13796
rect 3418 13716 3424 13728
rect 3252 13688 3424 13716
rect 3418 13676 3424 13688
rect 3476 13676 3482 13728
rect 4724 13716 4752 13815
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 5721 13855 5779 13861
rect 5721 13821 5733 13855
rect 5767 13852 5779 13855
rect 6270 13852 6276 13864
rect 5767 13824 6276 13852
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 6270 13812 6276 13824
rect 6328 13812 6334 13864
rect 6748 13852 6776 13892
rect 7558 13880 7564 13932
rect 7616 13920 7622 13932
rect 9398 13920 9404 13932
rect 7616 13892 7880 13920
rect 7616 13880 7622 13892
rect 7852 13864 7880 13892
rect 8680 13892 9260 13920
rect 9359 13892 9404 13920
rect 7466 13852 7472 13864
rect 6748 13824 7472 13852
rect 7466 13812 7472 13824
rect 7524 13852 7530 13864
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7524 13824 7757 13852
rect 7524 13812 7530 13824
rect 7745 13821 7757 13824
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 7834 13812 7840 13864
rect 7892 13852 7898 13864
rect 7929 13855 7987 13861
rect 7929 13852 7941 13855
rect 7892 13824 7941 13852
rect 7892 13812 7898 13824
rect 7929 13821 7941 13824
rect 7975 13821 7987 13855
rect 7929 13815 7987 13821
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 8352 13824 8401 13852
rect 8352 13812 8358 13824
rect 8389 13821 8401 13824
rect 8435 13821 8447 13855
rect 8389 13815 8447 13821
rect 6822 13784 6828 13796
rect 5828 13756 6828 13784
rect 5169 13719 5227 13725
rect 5169 13716 5181 13719
rect 4724 13688 5181 13716
rect 5169 13685 5181 13688
rect 5215 13716 5227 13719
rect 5828 13716 5856 13756
rect 6822 13744 6828 13756
rect 6880 13784 6886 13796
rect 7377 13787 7435 13793
rect 7377 13784 7389 13787
rect 6880 13756 7389 13784
rect 6880 13744 6886 13756
rect 7377 13753 7389 13756
rect 7423 13784 7435 13787
rect 8680 13784 8708 13892
rect 8757 13855 8815 13861
rect 8757 13821 8769 13855
rect 8803 13821 8815 13855
rect 8757 13815 8815 13821
rect 7423 13756 8708 13784
rect 7423 13753 7435 13756
rect 7377 13747 7435 13753
rect 5215 13688 5856 13716
rect 5905 13719 5963 13725
rect 5215 13685 5227 13688
rect 5169 13679 5227 13685
rect 5905 13685 5917 13719
rect 5951 13716 5963 13719
rect 6178 13716 6184 13728
rect 5951 13688 6184 13716
rect 5951 13685 5963 13688
rect 5905 13679 5963 13685
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 6917 13719 6975 13725
rect 6917 13685 6929 13719
rect 6963 13716 6975 13719
rect 7834 13716 7840 13728
rect 6963 13688 7840 13716
rect 6963 13685 6975 13688
rect 6917 13679 6975 13685
rect 7834 13676 7840 13688
rect 7892 13676 7898 13728
rect 7926 13676 7932 13728
rect 7984 13716 7990 13728
rect 8772 13716 8800 13815
rect 8938 13812 8944 13864
rect 8996 13852 9002 13864
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 8996 13824 9137 13852
rect 8996 13812 9002 13824
rect 9125 13821 9137 13824
rect 9171 13821 9183 13855
rect 9232 13852 9260 13892
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 9692 13920 9720 14016
rect 9953 13991 10011 13997
rect 9953 13957 9965 13991
rect 9999 13988 10011 13991
rect 10134 13988 10140 14000
rect 9999 13960 10140 13988
rect 9999 13957 10011 13960
rect 9953 13951 10011 13957
rect 10134 13948 10140 13960
rect 10192 13988 10198 14000
rect 10321 13991 10379 13997
rect 10321 13988 10333 13991
rect 10192 13960 10333 13988
rect 10192 13948 10198 13960
rect 10321 13957 10333 13960
rect 10367 13957 10379 13991
rect 10321 13951 10379 13957
rect 10870 13948 10876 14000
rect 10928 13988 10934 14000
rect 11241 13991 11299 13997
rect 11241 13988 11253 13991
rect 10928 13960 11253 13988
rect 10928 13948 10934 13960
rect 11241 13957 11253 13960
rect 11287 13957 11299 13991
rect 13998 13988 14004 14000
rect 13959 13960 14004 13988
rect 11241 13951 11299 13957
rect 13998 13948 14004 13960
rect 14056 13948 14062 14000
rect 20806 13948 20812 14000
rect 20864 13988 20870 14000
rect 21453 13991 21511 13997
rect 21453 13988 21465 13991
rect 20864 13960 21465 13988
rect 20864 13948 20870 13960
rect 21453 13957 21465 13960
rect 21499 13957 21511 13991
rect 21453 13951 21511 13957
rect 24663 13960 25544 13988
rect 13173 13923 13231 13929
rect 9692 13892 10272 13920
rect 10244 13861 10272 13892
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13262 13920 13268 13932
rect 13219 13892 13268 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 14366 13880 14372 13932
rect 14424 13920 14430 13932
rect 15105 13923 15163 13929
rect 14424 13892 14504 13920
rect 14424 13880 14430 13892
rect 9953 13855 10011 13861
rect 9953 13852 9965 13855
rect 9232 13824 9965 13852
rect 9125 13815 9183 13821
rect 9953 13821 9965 13824
rect 9999 13852 10011 13855
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 9999 13824 10057 13852
rect 9999 13821 10011 13824
rect 9953 13815 10011 13821
rect 10045 13821 10057 13824
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 10229 13855 10287 13861
rect 10229 13821 10241 13855
rect 10275 13821 10287 13855
rect 10502 13852 10508 13864
rect 10463 13824 10508 13852
rect 10229 13815 10287 13821
rect 10502 13812 10508 13824
rect 10560 13812 10566 13864
rect 14476 13861 14504 13892
rect 15105 13889 15117 13923
rect 15151 13920 15163 13923
rect 15286 13920 15292 13932
rect 15151 13892 15292 13920
rect 15151 13889 15163 13892
rect 15105 13883 15163 13889
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15396 13892 15853 13920
rect 14461 13855 14519 13861
rect 14461 13821 14473 13855
rect 14507 13821 14519 13855
rect 14461 13815 14519 13821
rect 14826 13812 14832 13864
rect 14884 13852 14890 13864
rect 14921 13855 14979 13861
rect 14921 13852 14933 13855
rect 14884 13824 14933 13852
rect 14884 13812 14890 13824
rect 14921 13821 14933 13824
rect 14967 13852 14979 13855
rect 15396 13852 15424 13892
rect 15841 13889 15853 13892
rect 15887 13920 15899 13923
rect 15887 13892 16436 13920
rect 15887 13889 15899 13892
rect 15841 13883 15899 13889
rect 16408 13864 16436 13892
rect 18230 13880 18236 13932
rect 18288 13920 18294 13932
rect 18417 13923 18475 13929
rect 18417 13920 18429 13923
rect 18288 13892 18429 13920
rect 18288 13880 18294 13892
rect 18417 13889 18429 13892
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 15930 13852 15936 13864
rect 14967 13824 15424 13852
rect 15891 13824 15936 13852
rect 14967 13821 14979 13824
rect 14921 13815 14979 13821
rect 15930 13812 15936 13824
rect 15988 13812 15994 13864
rect 16390 13812 16396 13864
rect 16448 13852 16454 13864
rect 16485 13855 16543 13861
rect 16485 13852 16497 13855
rect 16448 13824 16497 13852
rect 16448 13812 16454 13824
rect 16485 13821 16497 13824
rect 16531 13852 16543 13855
rect 17770 13852 17776 13864
rect 16531 13824 17776 13852
rect 16531 13821 16543 13824
rect 16485 13815 16543 13821
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 19680 13855 19738 13861
rect 19680 13821 19692 13855
rect 19726 13852 19738 13855
rect 20070 13852 20076 13864
rect 19726 13824 20076 13852
rect 19726 13821 19738 13824
rect 19680 13815 19738 13821
rect 20070 13812 20076 13824
rect 20128 13852 20134 13864
rect 24663 13861 24691 13960
rect 20660 13855 20718 13861
rect 20660 13852 20672 13855
rect 20128 13824 20672 13852
rect 20128 13812 20134 13824
rect 20660 13821 20672 13824
rect 20706 13852 20718 13855
rect 21085 13855 21143 13861
rect 21085 13852 21097 13855
rect 20706 13824 21097 13852
rect 20706 13821 20718 13824
rect 20660 13815 20718 13821
rect 21085 13821 21097 13824
rect 21131 13821 21143 13855
rect 21085 13815 21143 13821
rect 24648 13855 24706 13861
rect 24648 13821 24660 13855
rect 24694 13821 24706 13855
rect 24648 13815 24706 13821
rect 10962 13784 10968 13796
rect 10923 13756 10968 13784
rect 10962 13744 10968 13756
rect 11020 13744 11026 13796
rect 12158 13744 12164 13796
rect 12216 13784 12222 13796
rect 12526 13784 12532 13796
rect 12216 13756 12532 13784
rect 12216 13744 12222 13756
rect 12526 13744 12532 13756
rect 12584 13744 12590 13796
rect 12618 13744 12624 13796
rect 12676 13784 12682 13796
rect 13538 13784 13544 13796
rect 12676 13756 13544 13784
rect 12676 13744 12682 13756
rect 13538 13744 13544 13756
rect 13596 13744 13602 13796
rect 18138 13784 18144 13796
rect 18051 13756 18144 13784
rect 18138 13744 18144 13756
rect 18196 13744 18202 13796
rect 18233 13787 18291 13793
rect 18233 13753 18245 13787
rect 18279 13784 18291 13787
rect 18322 13784 18328 13796
rect 18279 13756 18328 13784
rect 18279 13753 18291 13756
rect 18233 13747 18291 13753
rect 18322 13744 18328 13756
rect 18380 13744 18386 13796
rect 25516 13793 25544 13960
rect 25501 13787 25559 13793
rect 25501 13784 25513 13787
rect 18432 13756 19656 13784
rect 25411 13756 25513 13784
rect 7984 13688 8800 13716
rect 7984 13676 7990 13688
rect 14826 13676 14832 13728
rect 14884 13716 14890 13728
rect 15381 13719 15439 13725
rect 15381 13716 15393 13719
rect 14884 13688 15393 13716
rect 14884 13676 14890 13688
rect 15381 13685 15393 13688
rect 15427 13716 15439 13719
rect 15470 13716 15476 13728
rect 15427 13688 15476 13716
rect 15427 13685 15439 13688
rect 15381 13679 15439 13685
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 15838 13676 15844 13728
rect 15896 13716 15902 13728
rect 16025 13719 16083 13725
rect 16025 13716 16037 13719
rect 15896 13688 16037 13716
rect 15896 13676 15902 13688
rect 16025 13685 16037 13688
rect 16071 13685 16083 13719
rect 18156 13716 18184 13744
rect 18432 13716 18460 13756
rect 19426 13716 19432 13728
rect 18156 13688 18460 13716
rect 19387 13688 19432 13716
rect 16025 13679 16083 13685
rect 19426 13676 19432 13688
rect 19484 13676 19490 13728
rect 19628 13716 19656 13756
rect 25501 13753 25513 13756
rect 25547 13784 25559 13787
rect 26234 13784 26240 13796
rect 25547 13756 26240 13784
rect 25547 13753 25559 13756
rect 25501 13747 25559 13753
rect 26234 13744 26240 13756
rect 26292 13744 26298 13796
rect 19751 13719 19809 13725
rect 19751 13716 19763 13719
rect 19628 13688 19763 13716
rect 19751 13685 19763 13688
rect 19797 13685 19809 13719
rect 19751 13679 19809 13685
rect 20070 13676 20076 13728
rect 20128 13716 20134 13728
rect 20763 13719 20821 13725
rect 20763 13716 20775 13719
rect 20128 13688 20775 13716
rect 20128 13676 20134 13688
rect 20763 13685 20775 13688
rect 20809 13685 20821 13719
rect 20763 13679 20821 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 3237 13515 3295 13521
rect 3237 13512 3249 13515
rect 3108 13484 3249 13512
rect 3108 13472 3114 13484
rect 3237 13481 3249 13484
rect 3283 13481 3295 13515
rect 3237 13475 3295 13481
rect 3418 13472 3424 13524
rect 3476 13512 3482 13524
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 3476 13484 5825 13512
rect 3476 13472 3482 13484
rect 5813 13481 5825 13484
rect 5859 13481 5871 13515
rect 7558 13512 7564 13524
rect 7519 13484 7564 13512
rect 5813 13475 5871 13481
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 7742 13472 7748 13524
rect 7800 13512 7806 13524
rect 8294 13512 8300 13524
rect 7800 13484 8300 13512
rect 7800 13472 7806 13484
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 9674 13472 9680 13524
rect 9732 13512 9738 13524
rect 10229 13515 10287 13521
rect 10229 13512 10241 13515
rect 9732 13484 10241 13512
rect 9732 13472 9738 13484
rect 10229 13481 10241 13484
rect 10275 13481 10287 13515
rect 10229 13475 10287 13481
rect 10551 13515 10609 13521
rect 10551 13481 10563 13515
rect 10597 13512 10609 13515
rect 12158 13512 12164 13524
rect 10597 13484 12164 13512
rect 10597 13481 10609 13484
rect 10551 13475 10609 13481
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 12529 13515 12587 13521
rect 12529 13481 12541 13515
rect 12575 13512 12587 13515
rect 12618 13512 12624 13524
rect 12575 13484 12624 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 12986 13472 12992 13524
rect 13044 13512 13050 13524
rect 14366 13512 14372 13524
rect 13044 13484 13124 13512
rect 14327 13484 14372 13512
rect 13044 13472 13050 13484
rect 1670 13444 1676 13456
rect 1631 13416 1676 13444
rect 1670 13404 1676 13416
rect 1728 13404 1734 13456
rect 2222 13444 2228 13456
rect 2183 13416 2228 13444
rect 2222 13404 2228 13416
rect 2280 13404 2286 13456
rect 4062 13444 4068 13456
rect 4023 13416 4068 13444
rect 4062 13404 4068 13416
rect 4120 13404 4126 13456
rect 5074 13444 5080 13456
rect 5035 13416 5080 13444
rect 5074 13404 5080 13416
rect 5132 13404 5138 13456
rect 9306 13444 9312 13456
rect 7024 13416 9312 13444
rect 7024 13388 7052 13416
rect 3510 13336 3516 13388
rect 3568 13376 3574 13388
rect 4157 13379 4215 13385
rect 4157 13376 4169 13379
rect 3568 13348 4169 13376
rect 3568 13336 3574 13348
rect 4157 13345 4169 13348
rect 4203 13345 4215 13379
rect 4157 13339 4215 13345
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 6181 13379 6239 13385
rect 6181 13376 6193 13379
rect 5592 13348 6193 13376
rect 5592 13336 5598 13348
rect 6181 13345 6193 13348
rect 6227 13376 6239 13379
rect 6362 13376 6368 13388
rect 6227 13348 6368 13376
rect 6227 13345 6239 13348
rect 6181 13339 6239 13345
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 6454 13336 6460 13388
rect 6512 13376 6518 13388
rect 7006 13376 7012 13388
rect 6512 13348 7012 13376
rect 6512 13336 6518 13348
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 7926 13336 7932 13388
rect 7984 13376 7990 13388
rect 8312 13385 8340 13416
rect 9306 13404 9312 13416
rect 9364 13444 9370 13456
rect 9401 13447 9459 13453
rect 9401 13444 9413 13447
rect 9364 13416 9413 13444
rect 9364 13404 9370 13416
rect 9401 13413 9413 13416
rect 9447 13413 9459 13447
rect 11606 13444 11612 13456
rect 11567 13416 11612 13444
rect 9401 13407 9459 13413
rect 11606 13404 11612 13416
rect 11664 13404 11670 13456
rect 13096 13453 13124 13484
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 15105 13515 15163 13521
rect 15105 13481 15117 13515
rect 15151 13512 15163 13515
rect 15286 13512 15292 13524
rect 15151 13484 15292 13512
rect 15151 13481 15163 13484
rect 15105 13475 15163 13481
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 15930 13472 15936 13524
rect 15988 13512 15994 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 15988 13484 16313 13512
rect 15988 13472 15994 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 17218 13512 17224 13524
rect 17179 13484 17224 13512
rect 16301 13475 16359 13481
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 17451 13515 17509 13521
rect 17451 13481 17463 13515
rect 17497 13512 17509 13515
rect 18046 13512 18052 13524
rect 17497 13484 18052 13512
rect 17497 13481 17509 13484
rect 17451 13475 17509 13481
rect 18046 13472 18052 13484
rect 18104 13512 18110 13524
rect 19426 13512 19432 13524
rect 18104 13484 19432 13512
rect 18104 13472 18110 13484
rect 19426 13472 19432 13484
rect 19484 13472 19490 13524
rect 13081 13447 13139 13453
rect 13081 13413 13093 13447
rect 13127 13413 13139 13447
rect 13081 13407 13139 13413
rect 13173 13447 13231 13453
rect 13173 13413 13185 13447
rect 13219 13444 13231 13447
rect 13538 13444 13544 13456
rect 13219 13416 13544 13444
rect 13219 13413 13231 13416
rect 13173 13407 13231 13413
rect 13538 13404 13544 13416
rect 13596 13404 13602 13456
rect 16022 13444 16028 13456
rect 15983 13416 16028 13444
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 18230 13404 18236 13456
rect 18288 13444 18294 13456
rect 18506 13444 18512 13456
rect 18288 13416 18512 13444
rect 18288 13404 18294 13416
rect 18506 13404 18512 13416
rect 18564 13404 18570 13456
rect 19061 13447 19119 13453
rect 19061 13413 19073 13447
rect 19107 13444 19119 13447
rect 19242 13444 19248 13456
rect 19107 13416 19248 13444
rect 19107 13413 19119 13416
rect 19061 13407 19119 13413
rect 19242 13404 19248 13416
rect 19300 13404 19306 13456
rect 8021 13379 8079 13385
rect 8021 13376 8033 13379
rect 7984 13348 8033 13376
rect 7984 13336 7990 13348
rect 8021 13345 8033 13348
rect 8067 13345 8079 13379
rect 8021 13339 8079 13345
rect 8297 13379 8355 13385
rect 8297 13345 8309 13379
rect 8343 13345 8355 13379
rect 8297 13339 8355 13345
rect 10318 13336 10324 13388
rect 10376 13376 10382 13388
rect 10448 13379 10506 13385
rect 10448 13376 10460 13379
rect 10376 13348 10460 13376
rect 10376 13336 10382 13348
rect 10448 13345 10460 13348
rect 10494 13345 10506 13379
rect 10448 13339 10506 13345
rect 14090 13336 14096 13388
rect 14148 13376 14154 13388
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 14148 13348 15301 13376
rect 14148 13336 14154 13348
rect 15289 13345 15301 13348
rect 15335 13345 15347 13379
rect 15289 13339 15347 13345
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13376 15899 13379
rect 15930 13376 15936 13388
rect 15887 13348 15936 13376
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 15930 13336 15936 13348
rect 15988 13376 15994 13388
rect 16390 13376 16396 13388
rect 15988 13348 16396 13376
rect 15988 13336 15994 13348
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 17310 13376 17316 13388
rect 17271 13348 17316 13376
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 20806 13336 20812 13388
rect 20864 13376 20870 13388
rect 20936 13379 20994 13385
rect 20936 13376 20948 13379
rect 20864 13348 20948 13376
rect 20864 13336 20870 13348
rect 20936 13345 20948 13348
rect 20982 13345 20994 13379
rect 20936 13339 20994 13345
rect 23636 13379 23694 13385
rect 23636 13345 23648 13379
rect 23682 13376 23694 13379
rect 23842 13376 23848 13388
rect 23682 13348 23848 13376
rect 23682 13345 23694 13348
rect 23636 13339 23694 13345
rect 23842 13336 23848 13348
rect 23900 13336 23906 13388
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 1581 13311 1639 13317
rect 1581 13308 1593 13311
rect 1452 13280 1593 13308
rect 1452 13268 1458 13280
rect 1581 13277 1593 13280
rect 1627 13308 1639 13311
rect 2869 13311 2927 13317
rect 2869 13308 2881 13311
rect 1627 13280 2881 13308
rect 1627 13277 1639 13280
rect 1581 13271 1639 13277
rect 2869 13277 2881 13280
rect 2915 13277 2927 13311
rect 2869 13271 2927 13277
rect 3881 13311 3939 13317
rect 3881 13277 3893 13311
rect 3927 13308 3939 13311
rect 4706 13308 4712 13320
rect 3927 13280 4712 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13308 6975 13311
rect 7466 13308 7472 13320
rect 6963 13280 7472 13308
rect 6963 13277 6975 13280
rect 6917 13271 6975 13277
rect 7466 13268 7472 13280
rect 7524 13268 7530 13320
rect 8478 13308 8484 13320
rect 8439 13280 8484 13308
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 9858 13308 9864 13320
rect 9088 13280 9864 13308
rect 9088 13268 9094 13280
rect 9858 13268 9864 13280
rect 9916 13268 9922 13320
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 11882 13308 11888 13320
rect 11563 13280 11888 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 11882 13268 11888 13280
rect 11940 13308 11946 13320
rect 13354 13308 13360 13320
rect 11940 13280 12388 13308
rect 13315 13280 13360 13308
rect 11940 13268 11946 13280
rect 1486 13200 1492 13252
rect 1544 13240 1550 13252
rect 2593 13243 2651 13249
rect 2593 13240 2605 13243
rect 1544 13212 2605 13240
rect 1544 13200 1550 13212
rect 2593 13209 2605 13212
rect 2639 13240 2651 13243
rect 4522 13240 4528 13252
rect 2639 13212 4528 13240
rect 2639 13209 2651 13212
rect 2593 13203 2651 13209
rect 4522 13200 4528 13212
rect 4580 13240 4586 13252
rect 5445 13243 5503 13249
rect 5445 13240 5457 13243
rect 4580 13212 5457 13240
rect 4580 13200 4586 13212
rect 5445 13209 5457 13212
rect 5491 13209 5503 13243
rect 5445 13203 5503 13209
rect 6178 13200 6184 13252
rect 6236 13240 6242 13252
rect 6273 13243 6331 13249
rect 6273 13240 6285 13243
rect 6236 13212 6285 13240
rect 6236 13200 6242 13212
rect 6273 13209 6285 13212
rect 6319 13209 6331 13243
rect 6273 13203 6331 13209
rect 8113 13243 8171 13249
rect 8113 13209 8125 13243
rect 8159 13209 8171 13243
rect 8113 13203 8171 13209
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 5074 13172 5080 13184
rect 3384 13144 5080 13172
rect 3384 13132 3390 13144
rect 5074 13132 5080 13144
rect 5132 13132 5138 13184
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 7800 13144 7849 13172
rect 7800 13132 7806 13144
rect 7837 13141 7849 13144
rect 7883 13172 7895 13175
rect 8128 13172 8156 13203
rect 11790 13200 11796 13252
rect 11848 13240 11854 13252
rect 12069 13243 12127 13249
rect 12069 13240 12081 13243
rect 11848 13212 12081 13240
rect 11848 13200 11854 13212
rect 12069 13209 12081 13212
rect 12115 13209 12127 13243
rect 12360 13240 12388 13280
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 18233 13311 18291 13317
rect 18233 13308 18245 13311
rect 13786 13280 18245 13308
rect 13786 13240 13814 13280
rect 18233 13277 18245 13280
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 18417 13311 18475 13317
rect 18417 13277 18429 13311
rect 18463 13308 18475 13311
rect 19426 13308 19432 13320
rect 18463 13280 19432 13308
rect 18463 13277 18475 13280
rect 18417 13271 18475 13277
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 12360 13212 13814 13240
rect 12069 13203 12127 13209
rect 16482 13200 16488 13252
rect 16540 13240 16546 13252
rect 16761 13243 16819 13249
rect 16761 13240 16773 13243
rect 16540 13212 16773 13240
rect 16540 13200 16546 13212
rect 16761 13209 16773 13212
rect 16807 13240 16819 13243
rect 21039 13243 21097 13249
rect 21039 13240 21051 13243
rect 16807 13212 21051 13240
rect 16807 13209 16819 13212
rect 16761 13203 16819 13209
rect 21039 13209 21051 13212
rect 21085 13209 21097 13243
rect 21039 13203 21097 13209
rect 9122 13172 9128 13184
rect 7883 13144 8156 13172
rect 9083 13144 9128 13172
rect 7883 13141 7895 13144
rect 7837 13135 7895 13141
rect 9122 13132 9128 13144
rect 9180 13132 9186 13184
rect 10870 13172 10876 13184
rect 10831 13144 10876 13172
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 12526 13132 12532 13184
rect 12584 13172 12590 13184
rect 12805 13175 12863 13181
rect 12805 13172 12817 13175
rect 12584 13144 12817 13172
rect 12584 13132 12590 13144
rect 12805 13141 12817 13144
rect 12851 13141 12863 13175
rect 18138 13172 18144 13184
rect 18099 13144 18144 13172
rect 12805 13135 12863 13141
rect 18138 13132 18144 13144
rect 18196 13132 18202 13184
rect 18233 13175 18291 13181
rect 18233 13141 18245 13175
rect 18279 13172 18291 13175
rect 20162 13172 20168 13184
rect 18279 13144 20168 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 20162 13132 20168 13144
rect 20220 13132 20226 13184
rect 23707 13175 23765 13181
rect 23707 13141 23719 13175
rect 23753 13172 23765 13175
rect 24026 13172 24032 13184
rect 23753 13144 24032 13172
rect 23753 13141 23765 13144
rect 23707 13135 23765 13141
rect 24026 13132 24032 13144
rect 24084 13132 24090 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 2409 12971 2467 12977
rect 2409 12968 2421 12971
rect 1728 12940 2421 12968
rect 1728 12928 1734 12940
rect 2409 12937 2421 12940
rect 2455 12937 2467 12971
rect 2409 12931 2467 12937
rect 6362 12928 6368 12980
rect 6420 12968 6426 12980
rect 6549 12971 6607 12977
rect 6549 12968 6561 12971
rect 6420 12940 6561 12968
rect 6420 12928 6426 12940
rect 6549 12937 6561 12940
rect 6595 12937 6607 12971
rect 10318 12968 10324 12980
rect 10279 12940 10324 12968
rect 6549 12931 6607 12937
rect 10318 12928 10324 12940
rect 10376 12968 10382 12980
rect 12894 12968 12900 12980
rect 10376 12940 12900 12968
rect 10376 12928 10382 12940
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 12986 12928 12992 12980
rect 13044 12968 13050 12980
rect 13817 12971 13875 12977
rect 13817 12968 13829 12971
rect 13044 12940 13829 12968
rect 13044 12928 13050 12940
rect 13817 12937 13829 12940
rect 13863 12937 13875 12971
rect 14274 12968 14280 12980
rect 14235 12940 14280 12968
rect 13817 12931 13875 12937
rect 14274 12928 14280 12940
rect 14332 12968 14338 12980
rect 15930 12968 15936 12980
rect 14332 12940 14964 12968
rect 15891 12940 15936 12968
rect 14332 12928 14338 12940
rect 1489 12903 1547 12909
rect 1489 12869 1501 12903
rect 1535 12900 1547 12903
rect 2222 12900 2228 12912
rect 1535 12872 2228 12900
rect 1535 12869 1547 12872
rect 1489 12863 1547 12869
rect 2222 12860 2228 12872
rect 2280 12900 2286 12912
rect 3973 12903 4031 12909
rect 3973 12900 3985 12903
rect 2280 12872 3985 12900
rect 2280 12860 2286 12872
rect 3973 12869 3985 12872
rect 4019 12900 4031 12903
rect 4617 12903 4675 12909
rect 4617 12900 4629 12903
rect 4019 12872 4629 12900
rect 4019 12869 4031 12872
rect 3973 12863 4031 12869
rect 4617 12869 4629 12872
rect 4663 12869 4675 12903
rect 4617 12863 4675 12869
rect 5905 12903 5963 12909
rect 5905 12869 5917 12903
rect 5951 12900 5963 12903
rect 6454 12900 6460 12912
rect 5951 12872 6460 12900
rect 5951 12869 5963 12872
rect 5905 12863 5963 12869
rect 6454 12860 6460 12872
rect 6512 12860 6518 12912
rect 9953 12903 10011 12909
rect 9953 12869 9965 12903
rect 9999 12900 10011 12903
rect 10778 12900 10784 12912
rect 9999 12872 10784 12900
rect 9999 12869 10011 12872
rect 9953 12863 10011 12869
rect 10778 12860 10784 12872
rect 10836 12860 10842 12912
rect 11333 12903 11391 12909
rect 11333 12869 11345 12903
rect 11379 12869 11391 12903
rect 11333 12863 11391 12869
rect 14 12792 20 12844
rect 72 12832 78 12844
rect 72 12804 1716 12832
rect 72 12792 78 12804
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 1486 12764 1492 12776
rect 1443 12736 1492 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1486 12724 1492 12736
rect 1544 12724 1550 12776
rect 1688 12773 1716 12804
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4430 12832 4436 12844
rect 4304 12804 4436 12832
rect 4304 12792 4310 12804
rect 4430 12792 4436 12804
rect 4488 12792 4494 12844
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 10413 12835 10471 12841
rect 10413 12832 10425 12835
rect 9631 12804 10425 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 10413 12801 10425 12804
rect 10459 12832 10471 12835
rect 10870 12832 10876 12844
rect 10459 12804 10876 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11348 12832 11376 12863
rect 11790 12860 11796 12912
rect 11848 12900 11854 12912
rect 13081 12903 13139 12909
rect 13081 12900 13093 12903
rect 11848 12872 13093 12900
rect 11848 12860 11854 12872
rect 13081 12869 13093 12872
rect 13127 12869 13139 12903
rect 13081 12863 13139 12869
rect 14090 12860 14096 12912
rect 14148 12900 14154 12912
rect 14645 12903 14703 12909
rect 14645 12900 14657 12903
rect 14148 12872 14657 12900
rect 14148 12860 14154 12872
rect 14645 12869 14657 12872
rect 14691 12869 14703 12903
rect 14645 12863 14703 12869
rect 11606 12832 11612 12844
rect 11348 12804 11612 12832
rect 11606 12792 11612 12804
rect 11664 12832 11670 12844
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 11664 12804 11713 12832
rect 11664 12792 11670 12804
rect 11701 12801 11713 12804
rect 11747 12832 11759 12835
rect 13630 12832 13636 12844
rect 11747 12804 13636 12832
rect 11747 12801 11759 12804
rect 11701 12795 11759 12801
rect 13630 12792 13636 12804
rect 13688 12792 13694 12844
rect 14936 12841 14964 12940
rect 15930 12928 15936 12940
rect 15988 12928 15994 12980
rect 18506 12928 18512 12980
rect 18564 12968 18570 12980
rect 19061 12971 19119 12977
rect 19061 12968 19073 12971
rect 18564 12940 19073 12968
rect 18564 12928 18570 12940
rect 19061 12937 19073 12940
rect 19107 12937 19119 12971
rect 19426 12968 19432 12980
rect 19387 12940 19432 12968
rect 19061 12931 19119 12937
rect 19426 12928 19432 12940
rect 19484 12968 19490 12980
rect 19751 12971 19809 12977
rect 19751 12968 19763 12971
rect 19484 12940 19763 12968
rect 19484 12928 19490 12940
rect 19751 12937 19763 12940
rect 19797 12937 19809 12971
rect 19751 12931 19809 12937
rect 20806 12928 20812 12980
rect 20864 12968 20870 12980
rect 21085 12971 21143 12977
rect 21085 12968 21097 12971
rect 20864 12940 21097 12968
rect 20864 12928 20870 12940
rect 21085 12937 21097 12940
rect 21131 12937 21143 12971
rect 23842 12968 23848 12980
rect 23803 12940 23848 12968
rect 21085 12931 21143 12937
rect 23842 12928 23848 12940
rect 23900 12928 23906 12980
rect 17402 12860 17408 12912
rect 17460 12900 17466 12912
rect 17460 12872 20806 12900
rect 17460 12860 17466 12872
rect 14921 12835 14979 12841
rect 14921 12801 14933 12835
rect 14967 12801 14979 12835
rect 16482 12832 16488 12844
rect 16443 12804 16488 12832
rect 14921 12795 14979 12801
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 18138 12832 18144 12844
rect 18051 12804 18144 12832
rect 18138 12792 18144 12804
rect 18196 12832 18202 12844
rect 18966 12832 18972 12844
rect 18196 12804 18972 12832
rect 18196 12792 18202 12804
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 19150 12792 19156 12844
rect 19208 12832 19214 12844
rect 20778 12841 20806 12872
rect 20763 12835 20821 12841
rect 19208 12804 20275 12832
rect 19208 12792 19214 12804
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12764 1731 12767
rect 1854 12764 1860 12776
rect 1719 12736 1860 12764
rect 1719 12733 1731 12736
rect 1673 12727 1731 12733
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 4522 12764 4528 12776
rect 4483 12736 4528 12764
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 4801 12767 4859 12773
rect 4801 12733 4813 12767
rect 4847 12733 4859 12767
rect 4801 12727 4859 12733
rect 2130 12696 2136 12708
rect 2091 12668 2136 12696
rect 2130 12656 2136 12668
rect 2188 12656 2194 12708
rect 3050 12696 3056 12708
rect 3011 12668 3056 12696
rect 3050 12656 3056 12668
rect 3108 12656 3114 12708
rect 3145 12699 3203 12705
rect 3145 12665 3157 12699
rect 3191 12665 3203 12699
rect 3145 12659 3203 12665
rect 3697 12699 3755 12705
rect 3697 12665 3709 12699
rect 3743 12696 3755 12699
rect 3878 12696 3884 12708
rect 3743 12668 3884 12696
rect 3743 12665 3755 12668
rect 3697 12659 3755 12665
rect 2866 12628 2872 12640
rect 2827 12600 2872 12628
rect 2866 12588 2872 12600
rect 2924 12628 2930 12640
rect 3160 12628 3188 12659
rect 3878 12656 3884 12668
rect 3936 12656 3942 12708
rect 2924 12600 3188 12628
rect 2924 12588 2930 12600
rect 4246 12588 4252 12640
rect 4304 12628 4310 12640
rect 4341 12631 4399 12637
rect 4341 12628 4353 12631
rect 4304 12600 4353 12628
rect 4304 12588 4310 12600
rect 4341 12597 4353 12600
rect 4387 12628 4399 12631
rect 4816 12628 4844 12727
rect 4890 12724 4896 12776
rect 4948 12764 4954 12776
rect 7190 12764 7196 12776
rect 4948 12736 7196 12764
rect 4948 12724 4954 12736
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 8202 12764 8208 12776
rect 8163 12736 8208 12764
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12733 8631 12767
rect 9030 12764 9036 12776
rect 8991 12736 9036 12764
rect 8573 12727 8631 12733
rect 7561 12699 7619 12705
rect 7561 12696 7573 12699
rect 6196 12668 7573 12696
rect 6196 12640 6224 12668
rect 7561 12665 7573 12668
rect 7607 12696 7619 12699
rect 7742 12696 7748 12708
rect 7607 12668 7748 12696
rect 7607 12665 7619 12668
rect 7561 12659 7619 12665
rect 7742 12656 7748 12668
rect 7800 12696 7806 12708
rect 8588 12696 8616 12727
rect 9030 12724 9036 12736
rect 9088 12724 9094 12776
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 9122 12696 9128 12708
rect 7800 12668 8616 12696
rect 8909 12668 9128 12696
rect 7800 12656 7806 12668
rect 4982 12628 4988 12640
rect 4387 12600 4844 12628
rect 4943 12600 4988 12628
rect 4387 12597 4399 12600
rect 4341 12591 4399 12597
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 6178 12628 6184 12640
rect 6139 12600 6184 12628
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 6825 12631 6883 12637
rect 6825 12597 6837 12631
rect 6871 12628 6883 12631
rect 6914 12628 6920 12640
rect 6871 12600 6920 12628
rect 6871 12597 6883 12600
rect 6825 12591 6883 12597
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 7926 12628 7932 12640
rect 7887 12600 7932 12628
rect 7926 12588 7932 12600
rect 7984 12588 7990 12640
rect 8570 12588 8576 12640
rect 8628 12628 8634 12640
rect 8909 12628 8937 12668
rect 9122 12656 9128 12668
rect 9180 12696 9186 12708
rect 9324 12696 9352 12727
rect 17126 12724 17132 12776
rect 17184 12764 17190 12776
rect 17954 12764 17960 12776
rect 17184 12736 17960 12764
rect 17184 12724 17190 12736
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 19680 12767 19738 12773
rect 19680 12733 19692 12767
rect 19726 12764 19738 12767
rect 20247 12764 20275 12804
rect 20763 12801 20775 12835
rect 20809 12801 20821 12835
rect 20763 12795 20821 12801
rect 20676 12767 20734 12773
rect 20676 12764 20688 12767
rect 19726 12736 20208 12764
rect 20247 12736 20688 12764
rect 19726 12733 19738 12736
rect 19680 12727 19738 12733
rect 12526 12696 12532 12708
rect 9180 12668 9352 12696
rect 12487 12668 12532 12696
rect 9180 12656 9186 12668
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 12621 12699 12679 12705
rect 12621 12665 12633 12699
rect 12667 12665 12679 12699
rect 15010 12696 15016 12708
rect 14971 12668 15016 12696
rect 12621 12659 12679 12665
rect 10778 12628 10784 12640
rect 8628 12600 8937 12628
rect 10739 12600 10784 12628
rect 8628 12588 8634 12600
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 12250 12628 12256 12640
rect 12163 12600 12256 12628
rect 12250 12588 12256 12600
rect 12308 12628 12314 12640
rect 12636 12628 12664 12659
rect 15010 12656 15016 12668
rect 15068 12656 15074 12708
rect 15565 12699 15623 12705
rect 15565 12665 15577 12699
rect 15611 12696 15623 12699
rect 15654 12696 15660 12708
rect 15611 12668 15660 12696
rect 15611 12665 15623 12668
rect 15565 12659 15623 12665
rect 15654 12656 15660 12668
rect 15712 12656 15718 12708
rect 16577 12699 16635 12705
rect 16577 12665 16589 12699
rect 16623 12665 16635 12699
rect 18230 12696 18236 12708
rect 16577 12659 16635 12665
rect 17788 12668 18236 12696
rect 12308 12600 12664 12628
rect 13541 12631 13599 12637
rect 12308 12588 12314 12600
rect 13541 12597 13553 12631
rect 13587 12628 13599 12631
rect 13630 12628 13636 12640
rect 13587 12600 13636 12628
rect 13587 12597 13599 12600
rect 13541 12591 13599 12597
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 16206 12628 16212 12640
rect 16167 12600 16212 12628
rect 16206 12588 16212 12600
rect 16264 12628 16270 12640
rect 16592 12628 16620 12659
rect 17402 12628 17408 12640
rect 16264 12600 16620 12628
rect 17363 12600 17408 12628
rect 16264 12588 16270 12600
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 17494 12588 17500 12640
rect 17552 12628 17558 12640
rect 17788 12637 17816 12668
rect 18230 12656 18236 12668
rect 18288 12656 18294 12708
rect 18785 12699 18843 12705
rect 18785 12665 18797 12699
rect 18831 12665 18843 12699
rect 18785 12659 18843 12665
rect 17773 12631 17831 12637
rect 17773 12628 17785 12631
rect 17552 12600 17785 12628
rect 17552 12588 17558 12600
rect 17773 12597 17785 12600
rect 17819 12597 17831 12631
rect 17773 12591 17831 12597
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 18800 12628 18828 12659
rect 20180 12640 20208 12736
rect 20676 12733 20688 12736
rect 20722 12764 20734 12767
rect 21453 12767 21511 12773
rect 21453 12764 21465 12767
rect 20722 12736 21465 12764
rect 20722 12733 20734 12736
rect 20676 12727 20734 12733
rect 21453 12733 21465 12736
rect 21499 12733 21511 12767
rect 21453 12727 21511 12733
rect 20162 12628 20168 12640
rect 18012 12600 18828 12628
rect 20123 12600 20168 12628
rect 18012 12588 18018 12600
rect 20162 12588 20168 12600
rect 20220 12588 20226 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1854 12424 1860 12436
rect 1815 12396 1860 12424
rect 1854 12384 1860 12396
rect 1912 12384 1918 12436
rect 2866 12424 2872 12436
rect 2827 12396 2872 12424
rect 2866 12384 2872 12396
rect 2924 12384 2930 12436
rect 3510 12424 3516 12436
rect 3471 12396 3516 12424
rect 3510 12384 3516 12396
rect 3568 12384 3574 12436
rect 3786 12424 3792 12436
rect 3747 12396 3792 12424
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4212 12396 4257 12424
rect 4212 12384 4218 12396
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 7009 12427 7067 12433
rect 7009 12424 7021 12427
rect 6052 12396 7021 12424
rect 6052 12384 6058 12396
rect 7009 12393 7021 12396
rect 7055 12424 7067 12427
rect 8570 12424 8576 12436
rect 7055 12396 8576 12424
rect 7055 12393 7067 12396
rect 7009 12387 7067 12393
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 8938 12384 8944 12436
rect 8996 12424 9002 12436
rect 9398 12424 9404 12436
rect 8996 12396 9404 12424
rect 8996 12384 9002 12396
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 9766 12424 9772 12436
rect 9727 12396 9772 12424
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 11882 12424 11888 12436
rect 11843 12396 11888 12424
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 12066 12384 12072 12436
rect 12124 12424 12130 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 12124 12396 13093 12424
rect 12124 12384 12130 12396
rect 13081 12393 13093 12396
rect 13127 12424 13139 12427
rect 13354 12424 13360 12436
rect 13127 12396 13360 12424
rect 13127 12393 13139 12396
rect 13081 12387 13139 12393
rect 13354 12384 13360 12396
rect 13412 12384 13418 12436
rect 14921 12427 14979 12433
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 15010 12424 15016 12436
rect 14967 12396 15016 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 15010 12384 15016 12396
rect 15068 12424 15074 12436
rect 15378 12424 15384 12436
rect 15068 12396 15384 12424
rect 15068 12384 15074 12396
rect 15378 12384 15384 12396
rect 15436 12424 15442 12436
rect 17494 12424 17500 12436
rect 15436 12396 17500 12424
rect 15436 12384 15442 12396
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 17586 12384 17592 12436
rect 17644 12424 17650 12436
rect 17644 12396 19288 12424
rect 17644 12384 17650 12396
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 2866 12288 2872 12300
rect 2827 12260 2872 12288
rect 2866 12248 2872 12260
rect 2924 12248 2930 12300
rect 3804 12288 3832 12384
rect 7374 12316 7380 12368
rect 7432 12356 7438 12368
rect 9416 12356 9444 12384
rect 7432 12328 8754 12356
rect 9416 12328 10916 12356
rect 7432 12316 7438 12328
rect 4341 12291 4399 12297
rect 4341 12288 4353 12291
rect 3804 12260 4353 12288
rect 4341 12257 4353 12260
rect 4387 12257 4399 12291
rect 4798 12288 4804 12300
rect 4759 12260 4804 12288
rect 4341 12251 4399 12257
rect 4356 12220 4384 12251
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 4985 12291 5043 12297
rect 4985 12257 4997 12291
rect 5031 12257 5043 12291
rect 4985 12251 5043 12257
rect 5000 12220 5028 12251
rect 5074 12248 5080 12300
rect 5132 12288 5138 12300
rect 5261 12291 5319 12297
rect 5261 12288 5273 12291
rect 5132 12260 5273 12288
rect 5132 12248 5138 12260
rect 5261 12257 5273 12260
rect 5307 12257 5319 12291
rect 5261 12251 5319 12257
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12288 6883 12291
rect 7561 12291 7619 12297
rect 7561 12288 7573 12291
rect 6871 12260 7573 12288
rect 6871 12257 6883 12260
rect 6825 12251 6883 12257
rect 7561 12257 7573 12260
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 5442 12220 5448 12232
rect 4356 12192 4752 12220
rect 5000 12192 5448 12220
rect 4724 12164 4752 12192
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 7576 12220 7604 12251
rect 7650 12248 7656 12300
rect 7708 12288 7714 12300
rect 8312 12297 8340 12328
rect 7745 12291 7803 12297
rect 7745 12288 7757 12291
rect 7708 12260 7757 12288
rect 7708 12248 7714 12260
rect 7745 12257 7757 12260
rect 7791 12257 7803 12291
rect 7745 12251 7803 12257
rect 8297 12291 8355 12297
rect 8297 12257 8309 12291
rect 8343 12257 8355 12291
rect 8570 12288 8576 12300
rect 8531 12260 8576 12288
rect 8297 12251 8355 12257
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 8726 12288 8754 12328
rect 9858 12288 9864 12300
rect 8726 12260 9864 12288
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 9953 12291 10011 12297
rect 9953 12257 9965 12291
rect 9999 12257 10011 12291
rect 9953 12251 10011 12257
rect 8018 12220 8024 12232
rect 7576 12192 8024 12220
rect 8018 12180 8024 12192
rect 8076 12220 8082 12232
rect 9968 12220 9996 12251
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 10137 12291 10195 12297
rect 10137 12288 10149 12291
rect 10100 12260 10149 12288
rect 10100 12248 10106 12260
rect 10137 12257 10149 12260
rect 10183 12257 10195 12291
rect 10502 12288 10508 12300
rect 10463 12260 10508 12288
rect 10137 12251 10195 12257
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 10888 12297 10916 12328
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 12161 12359 12219 12365
rect 12161 12356 12173 12359
rect 11572 12328 12173 12356
rect 11572 12316 11578 12328
rect 12161 12325 12173 12328
rect 12207 12325 12219 12359
rect 12161 12319 12219 12325
rect 15930 12316 15936 12368
rect 15988 12356 15994 12368
rect 16254 12359 16312 12365
rect 16254 12356 16266 12359
rect 15988 12328 16266 12356
rect 15988 12316 15994 12328
rect 16254 12325 16266 12328
rect 16300 12325 16312 12359
rect 17770 12356 17776 12368
rect 17731 12328 17776 12356
rect 16254 12319 16312 12325
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 17862 12316 17868 12368
rect 17920 12356 17926 12368
rect 17920 12328 17965 12356
rect 17920 12316 17926 12328
rect 19260 12300 19288 12396
rect 10873 12291 10931 12297
rect 10873 12257 10885 12291
rect 10919 12288 10931 12291
rect 10962 12288 10968 12300
rect 10919 12260 10968 12288
rect 10919 12257 10931 12260
rect 10873 12251 10931 12257
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 13630 12288 13636 12300
rect 13591 12260 13636 12288
rect 13630 12248 13636 12260
rect 13688 12248 13694 12300
rect 19242 12288 19248 12300
rect 19155 12260 19248 12288
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 19426 12248 19432 12300
rect 19484 12288 19490 12300
rect 19705 12291 19763 12297
rect 19705 12288 19717 12291
rect 19484 12260 19717 12288
rect 19484 12248 19490 12260
rect 19705 12257 19717 12260
rect 19751 12257 19763 12291
rect 19705 12251 19763 12257
rect 20968 12291 21026 12297
rect 20968 12257 20980 12291
rect 21014 12288 21026 12291
rect 21450 12288 21456 12300
rect 21014 12260 21456 12288
rect 21014 12257 21026 12260
rect 20968 12251 21026 12257
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 23636 12291 23694 12297
rect 23636 12257 23648 12291
rect 23682 12288 23694 12291
rect 23842 12288 23848 12300
rect 23682 12260 23848 12288
rect 23682 12257 23694 12260
rect 23636 12251 23694 12257
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 11422 12220 11428 12232
rect 8076 12192 11428 12220
rect 8076 12180 8082 12192
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 12066 12220 12072 12232
rect 12027 12192 12072 12220
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 12250 12180 12256 12232
rect 12308 12220 12314 12232
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 12308 12192 13553 12220
rect 12308 12180 12314 12192
rect 13541 12189 13553 12192
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12189 15991 12223
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 15933 12183 15991 12189
rect 17880 12192 19809 12220
rect 1581 12155 1639 12161
rect 1581 12121 1593 12155
rect 1627 12152 1639 12155
rect 4614 12152 4620 12164
rect 1627 12124 4620 12152
rect 1627 12121 1639 12124
rect 1581 12115 1639 12121
rect 4614 12112 4620 12124
rect 4672 12112 4678 12164
rect 4706 12112 4712 12164
rect 4764 12152 4770 12164
rect 5905 12155 5963 12161
rect 5905 12152 5917 12155
rect 4764 12124 5917 12152
rect 4764 12112 4770 12124
rect 5905 12121 5917 12124
rect 5951 12152 5963 12155
rect 8662 12152 8668 12164
rect 5951 12124 8248 12152
rect 8623 12124 8668 12152
rect 5951 12121 5963 12124
rect 5905 12115 5963 12121
rect 8220 12096 8248 12124
rect 8662 12112 8668 12124
rect 8720 12112 8726 12164
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 10502 12152 10508 12164
rect 9916 12124 10508 12152
rect 9916 12112 9922 12124
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 12618 12152 12624 12164
rect 12579 12124 12624 12152
rect 12618 12112 12624 12124
rect 12676 12112 12682 12164
rect 15948 12152 15976 12183
rect 16574 12152 16580 12164
rect 15948 12124 16580 12152
rect 16574 12112 16580 12124
rect 16632 12152 16638 12164
rect 17880 12152 17908 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 16632 12124 17908 12152
rect 18325 12155 18383 12161
rect 16632 12112 16638 12124
rect 18325 12121 18337 12155
rect 18371 12152 18383 12155
rect 18506 12152 18512 12164
rect 18371 12124 18512 12152
rect 18371 12121 18383 12124
rect 18325 12115 18383 12121
rect 18506 12112 18512 12124
rect 18564 12112 18570 12164
rect 2222 12084 2228 12096
rect 2183 12056 2228 12084
rect 2222 12044 2228 12056
rect 2280 12044 2286 12096
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 6181 12087 6239 12093
rect 6181 12084 6193 12087
rect 6052 12056 6193 12084
rect 6052 12044 6058 12056
rect 6181 12053 6193 12056
rect 6227 12053 6239 12087
rect 6181 12047 6239 12053
rect 6454 12044 6460 12096
rect 6512 12084 6518 12096
rect 7009 12087 7067 12093
rect 7009 12084 7021 12087
rect 6512 12056 7021 12084
rect 6512 12044 6518 12056
rect 7009 12053 7021 12056
rect 7055 12084 7067 12087
rect 7101 12087 7159 12093
rect 7101 12084 7113 12087
rect 7055 12056 7113 12084
rect 7055 12053 7067 12056
rect 7009 12047 7067 12053
rect 7101 12053 7113 12056
rect 7147 12053 7159 12087
rect 7101 12047 7159 12053
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 9033 12087 9091 12093
rect 9033 12084 9045 12087
rect 8260 12056 9045 12084
rect 8260 12044 8266 12056
rect 9033 12053 9045 12056
rect 9079 12053 9091 12087
rect 9033 12047 9091 12053
rect 10410 12044 10416 12096
rect 10468 12084 10474 12096
rect 11425 12087 11483 12093
rect 11425 12084 11437 12087
rect 10468 12056 11437 12084
rect 10468 12044 10474 12056
rect 11425 12053 11437 12056
rect 11471 12053 11483 12087
rect 11425 12047 11483 12053
rect 16853 12087 16911 12093
rect 16853 12053 16865 12087
rect 16899 12084 16911 12087
rect 16942 12084 16948 12096
rect 16899 12056 16948 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 16942 12044 16948 12056
rect 17000 12044 17006 12096
rect 17218 12084 17224 12096
rect 17131 12056 17224 12084
rect 17218 12044 17224 12056
rect 17276 12084 17282 12096
rect 18414 12084 18420 12096
rect 17276 12056 18420 12084
rect 17276 12044 17282 12056
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 18782 12084 18788 12096
rect 18743 12056 18788 12084
rect 18782 12044 18788 12056
rect 18840 12044 18846 12096
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 21039 12087 21097 12093
rect 21039 12084 21051 12087
rect 18932 12056 21051 12084
rect 18932 12044 18938 12056
rect 21039 12053 21051 12056
rect 21085 12053 21097 12087
rect 21039 12047 21097 12053
rect 23707 12087 23765 12093
rect 23707 12053 23719 12087
rect 23753 12084 23765 12087
rect 24118 12084 24124 12096
rect 23753 12056 24124 12084
rect 23753 12053 23765 12056
rect 23707 12047 23765 12053
rect 24118 12044 24124 12056
rect 24176 12044 24182 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 4890 11840 4896 11892
rect 4948 11880 4954 11892
rect 6178 11880 6184 11892
rect 4948 11852 6184 11880
rect 4948 11840 4954 11852
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 7009 11883 7067 11889
rect 7009 11849 7021 11883
rect 7055 11880 7067 11883
rect 7926 11880 7932 11892
rect 7055 11852 7932 11880
rect 7055 11849 7067 11852
rect 7009 11843 7067 11849
rect 7926 11840 7932 11852
rect 7984 11840 7990 11892
rect 9858 11880 9864 11892
rect 9819 11852 9864 11880
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 10321 11883 10379 11889
rect 10321 11849 10333 11883
rect 10367 11880 10379 11883
rect 10778 11880 10784 11892
rect 10367 11852 10784 11880
rect 10367 11849 10379 11852
rect 10321 11843 10379 11849
rect 10778 11840 10784 11852
rect 10836 11880 10842 11892
rect 13630 11880 13636 11892
rect 10836 11852 13492 11880
rect 13591 11852 13636 11880
rect 10836 11840 10842 11852
rect 2130 11772 2136 11824
rect 2188 11812 2194 11824
rect 6641 11815 6699 11821
rect 2188 11784 4154 11812
rect 2188 11772 2194 11784
rect 1535 11747 1593 11753
rect 1535 11713 1547 11747
rect 1581 11744 1593 11747
rect 3050 11744 3056 11756
rect 1581 11716 3056 11744
rect 1581 11713 1593 11716
rect 1535 11707 1593 11713
rect 3050 11704 3056 11716
rect 3108 11704 3114 11756
rect 4126 11744 4154 11784
rect 6641 11781 6653 11815
rect 6687 11812 6699 11815
rect 7650 11812 7656 11824
rect 6687 11784 7656 11812
rect 6687 11781 6699 11784
rect 6641 11775 6699 11781
rect 7650 11772 7656 11784
rect 7708 11772 7714 11824
rect 7834 11772 7840 11824
rect 7892 11812 7898 11824
rect 12342 11812 12348 11824
rect 7892 11784 12348 11812
rect 7892 11772 7898 11784
rect 12342 11772 12348 11784
rect 12400 11812 12406 11824
rect 13464 11812 13492 11852
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 15378 11880 15384 11892
rect 15339 11852 15384 11880
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 18782 11840 18788 11892
rect 18840 11880 18846 11892
rect 20763 11883 20821 11889
rect 20763 11880 20775 11883
rect 18840 11852 20775 11880
rect 18840 11840 18846 11852
rect 20763 11849 20775 11852
rect 20809 11849 20821 11883
rect 23842 11880 23848 11892
rect 23803 11852 23848 11880
rect 20763 11843 20821 11849
rect 23842 11840 23848 11852
rect 23900 11840 23906 11892
rect 24762 11880 24768 11892
rect 24723 11852 24768 11880
rect 24762 11840 24768 11852
rect 24820 11840 24826 11892
rect 14277 11815 14335 11821
rect 14277 11812 14289 11815
rect 12400 11784 12572 11812
rect 13464 11784 14289 11812
rect 12400 11772 12406 11784
rect 7374 11744 7380 11756
rect 4126 11716 6868 11744
rect 7335 11716 7380 11744
rect 1210 11636 1216 11688
rect 1268 11676 1274 11688
rect 1432 11679 1490 11685
rect 1432 11676 1444 11679
rect 1268 11648 1444 11676
rect 1268 11636 1274 11648
rect 1432 11645 1444 11648
rect 1478 11676 1490 11679
rect 1857 11679 1915 11685
rect 1857 11676 1869 11679
rect 1478 11648 1869 11676
rect 1478 11645 1490 11648
rect 1432 11639 1490 11645
rect 1857 11645 1869 11648
rect 1903 11645 1915 11679
rect 1857 11639 1915 11645
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11676 2743 11679
rect 2774 11676 2780 11688
rect 2731 11648 2780 11676
rect 2731 11645 2743 11648
rect 2685 11639 2743 11645
rect 2774 11636 2780 11648
rect 2832 11676 2838 11688
rect 4154 11676 4160 11688
rect 2832 11648 4160 11676
rect 2832 11636 2838 11648
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 4706 11676 4712 11688
rect 4667 11648 4712 11676
rect 4706 11636 4712 11648
rect 4764 11636 4770 11688
rect 4890 11676 4896 11688
rect 4851 11648 4896 11676
rect 4890 11636 4896 11648
rect 4948 11636 4954 11688
rect 5442 11676 5448 11688
rect 5355 11648 5448 11676
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 5813 11679 5871 11685
rect 5813 11676 5825 11679
rect 5592 11648 5825 11676
rect 5592 11636 5598 11648
rect 5813 11645 5825 11648
rect 5859 11676 5871 11679
rect 5994 11676 6000 11688
rect 5859 11648 6000 11676
rect 5859 11645 5871 11648
rect 5813 11639 5871 11645
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 6840 11685 6868 11716
rect 7374 11704 7380 11716
rect 7432 11704 7438 11756
rect 9030 11744 9036 11756
rect 8956 11716 9036 11744
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 7653 11679 7711 11685
rect 7653 11676 7665 11679
rect 6871 11648 7665 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 7653 11645 7665 11648
rect 7699 11645 7711 11679
rect 8202 11676 8208 11688
rect 8163 11648 8208 11676
rect 7653 11639 7711 11645
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8956 11685 8984 11716
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11744 9643 11747
rect 10410 11744 10416 11756
rect 9631 11716 10416 11744
rect 9631 11713 9643 11716
rect 9585 11707 9643 11713
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 12250 11744 12256 11756
rect 12211 11716 12256 11744
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 12544 11753 12572 11784
rect 14277 11781 14289 11784
rect 14323 11781 14335 11815
rect 14277 11775 14335 11781
rect 12529 11747 12587 11753
rect 12529 11713 12541 11747
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11744 13231 11747
rect 13354 11744 13360 11756
rect 13219 11716 13360 11744
rect 13219 11713 13231 11716
rect 13173 11707 13231 11713
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 14292 11744 14320 11775
rect 14826 11744 14832 11756
rect 14292 11716 14832 11744
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 15654 11704 15660 11756
rect 15712 11744 15718 11756
rect 16485 11747 16543 11753
rect 16485 11744 16497 11747
rect 15712 11716 16497 11744
rect 15712 11704 15718 11716
rect 16485 11713 16497 11716
rect 16531 11744 16543 11747
rect 17218 11744 17224 11756
rect 16531 11716 17224 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 18141 11747 18199 11753
rect 18141 11713 18153 11747
rect 18187 11744 18199 11747
rect 18800 11744 18828 11840
rect 18966 11772 18972 11824
rect 19024 11812 19030 11824
rect 19751 11815 19809 11821
rect 19751 11812 19763 11815
rect 19024 11784 19763 11812
rect 19024 11772 19030 11784
rect 19751 11781 19763 11784
rect 19797 11781 19809 11815
rect 19751 11775 19809 11781
rect 19242 11744 19248 11756
rect 18187 11716 18828 11744
rect 19203 11716 19248 11744
rect 18187 11713 18199 11716
rect 18141 11707 18199 11713
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11645 8631 11679
rect 8573 11639 8631 11645
rect 8941 11679 8999 11685
rect 8941 11645 8953 11679
rect 8987 11645 8999 11679
rect 9398 11676 9404 11688
rect 9359 11648 9404 11676
rect 8941 11639 8999 11645
rect 2590 11608 2596 11620
rect 2503 11580 2596 11608
rect 2590 11568 2596 11580
rect 2648 11608 2654 11620
rect 3006 11611 3064 11617
rect 3006 11608 3018 11611
rect 2648 11580 3018 11608
rect 2648 11568 2654 11580
rect 3006 11577 3018 11580
rect 3052 11608 3064 11611
rect 3510 11608 3516 11620
rect 3052 11580 3516 11608
rect 3052 11577 3064 11580
rect 3006 11571 3064 11577
rect 3510 11568 3516 11580
rect 3568 11568 3574 11620
rect 3602 11540 3608 11552
rect 3563 11512 3608 11540
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 4157 11543 4215 11549
rect 4157 11509 4169 11543
rect 4203 11540 4215 11543
rect 5074 11540 5080 11552
rect 4203 11512 5080 11540
rect 4203 11509 4215 11512
rect 4157 11503 4215 11509
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 5166 11500 5172 11552
rect 5224 11540 5230 11552
rect 5460 11540 5488 11636
rect 5905 11611 5963 11617
rect 5905 11577 5917 11611
rect 5951 11608 5963 11611
rect 6086 11608 6092 11620
rect 5951 11580 6092 11608
rect 5951 11577 5963 11580
rect 5905 11571 5963 11577
rect 6086 11568 6092 11580
rect 6144 11568 6150 11620
rect 7742 11568 7748 11620
rect 7800 11608 7806 11620
rect 8588 11608 8616 11639
rect 9398 11636 9404 11648
rect 9456 11636 9462 11688
rect 7800 11580 8616 11608
rect 12268 11608 12296 11704
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 13924 11648 14473 11676
rect 12621 11611 12679 11617
rect 12621 11608 12633 11611
rect 12268 11580 12633 11608
rect 7800 11568 7806 11580
rect 12621 11577 12633 11580
rect 12667 11577 12679 11611
rect 12621 11571 12679 11577
rect 13924 11552 13952 11648
rect 14461 11645 14473 11648
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 14844 11676 14872 11704
rect 15930 11676 15936 11688
rect 14844 11648 15936 11676
rect 14844 11617 14872 11648
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 18966 11636 18972 11688
rect 19024 11676 19030 11688
rect 19648 11679 19706 11685
rect 19648 11676 19660 11679
rect 19024 11648 19660 11676
rect 19024 11636 19030 11648
rect 19648 11645 19660 11648
rect 19694 11676 19706 11679
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 19694 11648 20085 11676
rect 19694 11645 19706 11648
rect 19648 11639 19706 11645
rect 20073 11645 20085 11648
rect 20119 11645 20131 11679
rect 20073 11639 20131 11645
rect 20692 11679 20750 11685
rect 20692 11645 20704 11679
rect 20738 11645 20750 11679
rect 20692 11639 20750 11645
rect 14823 11611 14881 11617
rect 14823 11577 14835 11611
rect 14869 11577 14881 11611
rect 14823 11571 14881 11577
rect 16577 11611 16635 11617
rect 16577 11577 16589 11611
rect 16623 11608 16635 11611
rect 16850 11608 16856 11620
rect 16623 11580 16856 11608
rect 16623 11577 16635 11580
rect 16577 11571 16635 11577
rect 16850 11568 16856 11580
rect 16908 11568 16914 11620
rect 17129 11611 17187 11617
rect 17129 11577 17141 11611
rect 17175 11608 17187 11611
rect 17310 11608 17316 11620
rect 17175 11580 17316 11608
rect 17175 11577 17187 11580
rect 17129 11571 17187 11577
rect 17310 11568 17316 11580
rect 17368 11568 17374 11620
rect 17402 11568 17408 11620
rect 17460 11608 17466 11620
rect 18230 11608 18236 11620
rect 17460 11580 18000 11608
rect 18191 11580 18236 11608
rect 17460 11568 17466 11580
rect 7374 11540 7380 11552
rect 5224 11512 7380 11540
rect 5224 11500 5230 11512
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 10778 11540 10784 11552
rect 10739 11512 10784 11540
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 11330 11540 11336 11552
rect 11291 11512 11336 11540
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 11514 11500 11520 11552
rect 11572 11540 11578 11552
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11572 11512 11805 11540
rect 11572 11500 11578 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 13906 11540 13912 11552
rect 13867 11512 13912 11540
rect 11793 11503 11851 11509
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 17681 11543 17739 11549
rect 17681 11540 17693 11543
rect 16264 11512 17693 11540
rect 16264 11500 16270 11512
rect 17681 11509 17693 11512
rect 17727 11540 17739 11543
rect 17862 11540 17868 11552
rect 17727 11512 17868 11540
rect 17727 11509 17739 11512
rect 17681 11503 17739 11509
rect 17862 11500 17868 11512
rect 17920 11500 17926 11552
rect 17972 11540 18000 11580
rect 18230 11568 18236 11580
rect 18288 11568 18294 11620
rect 18506 11568 18512 11620
rect 18564 11608 18570 11620
rect 18785 11611 18843 11617
rect 18785 11608 18797 11611
rect 18564 11580 18797 11608
rect 18564 11568 18570 11580
rect 18785 11577 18797 11580
rect 18831 11577 18843 11611
rect 20707 11608 20735 11639
rect 24118 11636 24124 11688
rect 24176 11676 24182 11688
rect 24581 11679 24639 11685
rect 24581 11676 24593 11679
rect 24176 11648 24593 11676
rect 24176 11636 24182 11648
rect 24581 11645 24593 11648
rect 24627 11676 24639 11679
rect 25133 11679 25191 11685
rect 25133 11676 25145 11679
rect 24627 11648 25145 11676
rect 24627 11645 24639 11648
rect 24581 11639 24639 11645
rect 25133 11645 25145 11648
rect 25179 11645 25191 11679
rect 25133 11639 25191 11645
rect 21177 11611 21235 11617
rect 21177 11608 21189 11611
rect 18785 11571 18843 11577
rect 18984 11580 21189 11608
rect 18984 11540 19012 11580
rect 21177 11577 21189 11580
rect 21223 11608 21235 11611
rect 25498 11608 25504 11620
rect 21223 11580 25504 11608
rect 21223 11577 21235 11580
rect 21177 11571 21235 11577
rect 25498 11568 25504 11580
rect 25556 11568 25562 11620
rect 21450 11540 21456 11552
rect 17972 11512 19012 11540
rect 21411 11512 21456 11540
rect 21450 11500 21456 11512
rect 21508 11500 21514 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 1854 11336 1860 11348
rect 1452 11308 1860 11336
rect 1452 11296 1458 11308
rect 1854 11296 1860 11308
rect 1912 11336 1918 11348
rect 2409 11339 2467 11345
rect 2409 11336 2421 11339
rect 1912 11308 2421 11336
rect 1912 11296 1918 11308
rect 2409 11305 2421 11308
rect 2455 11305 2467 11339
rect 2866 11336 2872 11348
rect 2827 11308 2872 11336
rect 2409 11299 2467 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 3881 11339 3939 11345
rect 3191 11308 3832 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 2884 11268 2912 11296
rect 3513 11271 3571 11277
rect 3513 11268 3525 11271
rect 2884 11240 3525 11268
rect 3513 11237 3525 11240
rect 3559 11268 3571 11271
rect 3602 11268 3608 11280
rect 3559 11240 3608 11268
rect 3559 11237 3571 11240
rect 3513 11231 3571 11237
rect 3602 11228 3608 11240
rect 3660 11228 3666 11280
rect 3804 11268 3832 11308
rect 3881 11305 3893 11339
rect 3927 11336 3939 11339
rect 4890 11336 4896 11348
rect 3927 11308 4896 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 4890 11296 4896 11308
rect 4948 11296 4954 11348
rect 4985 11339 5043 11345
rect 4985 11305 4997 11339
rect 5031 11336 5043 11339
rect 5166 11336 5172 11348
rect 5031 11308 5172 11336
rect 5031 11305 5043 11308
rect 4985 11299 5043 11305
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5442 11336 5448 11348
rect 5403 11308 5448 11336
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 7650 11296 7656 11348
rect 7708 11336 7714 11348
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 7708 11308 9413 11336
rect 7708 11296 7714 11308
rect 9401 11305 9413 11308
rect 9447 11336 9459 11339
rect 10042 11336 10048 11348
rect 9447 11308 10048 11336
rect 9447 11305 9459 11308
rect 9401 11299 9459 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 10962 11336 10968 11348
rect 10923 11308 10968 11336
rect 10962 11296 10968 11308
rect 11020 11296 11026 11348
rect 11422 11336 11428 11348
rect 11383 11308 11428 11336
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 12529 11339 12587 11345
rect 12529 11336 12541 11339
rect 12400 11308 12541 11336
rect 12400 11296 12406 11308
rect 12529 11305 12541 11308
rect 12575 11305 12587 11339
rect 16574 11336 16580 11348
rect 16535 11308 16580 11336
rect 12529 11299 12587 11305
rect 16574 11296 16580 11308
rect 16632 11296 16638 11348
rect 18141 11339 18199 11345
rect 18141 11305 18153 11339
rect 18187 11336 18199 11339
rect 18230 11336 18236 11348
rect 18187 11308 18236 11336
rect 18187 11305 18199 11308
rect 18141 11299 18199 11305
rect 18230 11296 18236 11308
rect 18288 11296 18294 11348
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 19613 11339 19671 11345
rect 19613 11336 19625 11339
rect 19484 11308 19625 11336
rect 19484 11296 19490 11308
rect 19613 11305 19625 11308
rect 19659 11336 19671 11339
rect 24762 11336 24768 11348
rect 19659 11308 19840 11336
rect 24723 11308 24768 11336
rect 19659 11305 19671 11308
rect 19613 11299 19671 11305
rect 19812 11280 19840 11308
rect 24762 11296 24768 11308
rect 24820 11296 24826 11348
rect 3804 11240 4568 11268
rect 1762 11200 1768 11212
rect 1723 11172 1768 11200
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 2961 11203 3019 11209
rect 2961 11169 2973 11203
rect 3007 11200 3019 11203
rect 3418 11200 3424 11212
rect 3007 11172 3424 11200
rect 3007 11169 3019 11172
rect 2961 11163 3019 11169
rect 3418 11160 3424 11172
rect 3476 11160 3482 11212
rect 4540 11209 4568 11240
rect 4614 11228 4620 11280
rect 4672 11268 4678 11280
rect 6638 11268 6644 11280
rect 4672 11240 6644 11268
rect 4672 11228 4678 11240
rect 6638 11228 6644 11240
rect 6696 11228 6702 11280
rect 7006 11268 7012 11280
rect 6967 11240 7012 11268
rect 7006 11228 7012 11240
rect 7064 11228 7070 11280
rect 7558 11268 7564 11280
rect 7519 11240 7564 11268
rect 7558 11228 7564 11240
rect 7616 11228 7622 11280
rect 7742 11228 7748 11280
rect 7800 11268 7806 11280
rect 8205 11271 8263 11277
rect 8205 11268 8217 11271
rect 7800 11240 8217 11268
rect 7800 11228 7806 11240
rect 8205 11237 8217 11240
rect 8251 11237 8263 11271
rect 8205 11231 8263 11237
rect 11330 11228 11336 11280
rect 11388 11268 11394 11280
rect 11701 11271 11759 11277
rect 11701 11268 11713 11271
rect 11388 11240 11713 11268
rect 11388 11228 11394 11240
rect 11701 11237 11713 11240
rect 11747 11237 11759 11271
rect 14182 11268 14188 11280
rect 11701 11231 11759 11237
rect 13924 11240 14188 11268
rect 4111 11203 4169 11209
rect 4111 11169 4123 11203
rect 4157 11169 4169 11203
rect 4111 11163 4169 11169
rect 4525 11203 4583 11209
rect 4525 11169 4537 11203
rect 4571 11200 4583 11203
rect 5166 11200 5172 11212
rect 4571 11172 5172 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 4126 11132 4154 11163
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 8110 11160 8116 11212
rect 8168 11200 8174 11212
rect 8570 11200 8576 11212
rect 8628 11209 8634 11212
rect 8628 11203 8666 11209
rect 8168 11172 8576 11200
rect 8168 11160 8174 11172
rect 8570 11160 8576 11172
rect 8654 11169 8666 11203
rect 8628 11163 8666 11169
rect 8628 11160 8634 11163
rect 9214 11160 9220 11212
rect 9272 11200 9278 11212
rect 9950 11200 9956 11212
rect 9272 11172 9956 11200
rect 9272 11160 9278 11172
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 10410 11200 10416 11212
rect 10371 11172 10416 11200
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 13924 11209 13952 11240
rect 14182 11228 14188 11240
rect 14240 11228 14246 11280
rect 15651 11271 15709 11277
rect 15651 11237 15663 11271
rect 15697 11268 15709 11271
rect 15930 11268 15936 11280
rect 15697 11240 15936 11268
rect 15697 11237 15709 11240
rect 15651 11231 15709 11237
rect 15930 11228 15936 11240
rect 15988 11228 15994 11280
rect 16942 11228 16948 11280
rect 17000 11268 17006 11280
rect 17221 11271 17279 11277
rect 17221 11268 17233 11271
rect 17000 11240 17233 11268
rect 17000 11228 17006 11240
rect 17221 11237 17233 11240
rect 17267 11237 17279 11271
rect 17221 11231 17279 11237
rect 17770 11228 17776 11280
rect 17828 11268 17834 11280
rect 18417 11271 18475 11277
rect 18417 11268 18429 11271
rect 17828 11240 18429 11268
rect 17828 11228 17834 11240
rect 18417 11237 18429 11240
rect 18463 11237 18475 11271
rect 18417 11231 18475 11237
rect 18785 11271 18843 11277
rect 18785 11237 18797 11271
rect 18831 11268 18843 11271
rect 19058 11268 19064 11280
rect 18831 11240 19064 11268
rect 18831 11237 18843 11240
rect 18785 11231 18843 11237
rect 19058 11228 19064 11240
rect 19116 11228 19122 11280
rect 19794 11228 19800 11280
rect 19852 11228 19858 11280
rect 13909 11203 13967 11209
rect 13909 11169 13921 11203
rect 13955 11169 13967 11203
rect 13909 11163 13967 11169
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 14093 11203 14151 11209
rect 14093 11200 14105 11203
rect 14056 11172 14105 11200
rect 14056 11160 14062 11172
rect 14093 11169 14105 11172
rect 14139 11169 14151 11203
rect 14093 11163 14151 11169
rect 20254 11160 20260 11212
rect 20312 11200 20318 11212
rect 21358 11200 21364 11212
rect 20312 11172 21364 11200
rect 20312 11160 20318 11172
rect 21358 11160 21364 11172
rect 21416 11160 21422 11212
rect 24026 11160 24032 11212
rect 24084 11200 24090 11212
rect 24581 11203 24639 11209
rect 24581 11200 24593 11203
rect 24084 11172 24593 11200
rect 24084 11160 24090 11172
rect 24581 11169 24593 11172
rect 24627 11200 24639 11203
rect 24670 11200 24676 11212
rect 24627 11172 24676 11200
rect 24627 11169 24639 11172
rect 24581 11163 24639 11169
rect 24670 11160 24676 11172
rect 24728 11160 24734 11212
rect 4706 11132 4712 11144
rect 4126 11104 4712 11132
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 6086 11132 6092 11144
rect 5123 11104 6092 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6914 11132 6920 11144
rect 6875 11104 6920 11132
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 10686 11132 10692 11144
rect 10647 11104 10692 11132
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 11609 11135 11667 11141
rect 11609 11101 11621 11135
rect 11655 11132 11667 11135
rect 11790 11132 11796 11144
rect 11655 11104 11796 11132
rect 11655 11101 11667 11104
rect 11609 11095 11667 11101
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11132 11943 11135
rect 12618 11132 12624 11144
rect 11931 11104 12624 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 3694 11024 3700 11076
rect 3752 11064 3758 11076
rect 4203 11067 4261 11073
rect 4203 11064 4215 11067
rect 3752 11036 4215 11064
rect 3752 11024 3758 11036
rect 4203 11033 4215 11036
rect 4249 11064 4261 11067
rect 6273 11067 6331 11073
rect 6273 11064 6285 11067
rect 4249 11036 6285 11064
rect 4249 11033 4261 11036
rect 4203 11027 4261 11033
rect 6273 11033 6285 11036
rect 6319 11033 6331 11067
rect 6273 11027 6331 11033
rect 11422 11024 11428 11076
rect 11480 11064 11486 11076
rect 11900 11064 11928 11095
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 14366 11132 14372 11144
rect 14327 11104 14372 11132
rect 14366 11092 14372 11104
rect 14424 11132 14430 11144
rect 15289 11135 15347 11141
rect 15289 11132 15301 11135
rect 14424 11104 15301 11132
rect 14424 11092 14430 11104
rect 15289 11101 15301 11104
rect 15335 11101 15347 11135
rect 17126 11132 17132 11144
rect 17087 11104 17132 11132
rect 15289 11095 15347 11101
rect 17126 11092 17132 11104
rect 17184 11132 17190 11144
rect 18690 11132 18696 11144
rect 17184 11104 18000 11132
rect 18651 11104 18696 11132
rect 17184 11092 17190 11104
rect 11480 11036 11928 11064
rect 11480 11024 11486 11036
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 17681 11067 17739 11073
rect 17681 11064 17693 11067
rect 17368 11036 17693 11064
rect 17368 11024 17374 11036
rect 17681 11033 17693 11036
rect 17727 11033 17739 11067
rect 17972 11064 18000 11104
rect 18690 11092 18696 11104
rect 18748 11092 18754 11144
rect 18969 11135 19027 11141
rect 18969 11101 18981 11135
rect 19015 11101 19027 11135
rect 18969 11095 19027 11101
rect 18984 11064 19012 11095
rect 17972 11036 19012 11064
rect 17681 11027 17739 11033
rect 1670 10996 1676 11008
rect 1631 10968 1676 10996
rect 1670 10956 1676 10968
rect 1728 10956 1734 11008
rect 5350 10956 5356 11008
rect 5408 10996 5414 11008
rect 5994 10996 6000 11008
rect 5408 10968 6000 10996
rect 5408 10956 5414 10968
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 8711 10999 8769 11005
rect 8711 10965 8723 10999
rect 8757 10996 8769 10999
rect 8938 10996 8944 11008
rect 8757 10968 8944 10996
rect 8757 10965 8769 10968
rect 8711 10959 8769 10965
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 9122 10996 9128 11008
rect 9083 10968 9128 10996
rect 9122 10956 9128 10968
rect 9180 10956 9186 11008
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 12897 10999 12955 11005
rect 12897 10996 12909 10999
rect 12768 10968 12909 10996
rect 12768 10956 12774 10968
rect 12897 10965 12909 10968
rect 12943 10965 12955 10999
rect 12897 10959 12955 10965
rect 14826 10956 14832 11008
rect 14884 10996 14890 11008
rect 14921 10999 14979 11005
rect 14921 10996 14933 10999
rect 14884 10968 14933 10996
rect 14884 10956 14890 10968
rect 14921 10965 14933 10968
rect 14967 10965 14979 10999
rect 16206 10996 16212 11008
rect 16167 10968 16212 10996
rect 14921 10959 14979 10965
rect 16206 10956 16212 10968
rect 16264 10956 16270 11008
rect 16850 10996 16856 11008
rect 16811 10968 16856 10996
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 17696 10996 17724 11027
rect 17862 10996 17868 11008
rect 17696 10968 17868 10996
rect 17862 10956 17868 10968
rect 17920 10996 17926 11008
rect 19150 10996 19156 11008
rect 17920 10968 19156 10996
rect 17920 10956 17926 10968
rect 19150 10956 19156 10968
rect 19208 10956 19214 11008
rect 21545 10999 21603 11005
rect 21545 10965 21557 10999
rect 21591 10996 21603 10999
rect 22186 10996 22192 11008
rect 21591 10968 22192 10996
rect 21591 10965 21603 10968
rect 21545 10959 21603 10965
rect 22186 10956 22192 10968
rect 22244 10956 22250 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 2406 10792 2412 10804
rect 1820 10764 2412 10792
rect 1820 10752 1826 10764
rect 2406 10752 2412 10764
rect 2464 10792 2470 10804
rect 2501 10795 2559 10801
rect 2501 10792 2513 10795
rect 2464 10764 2513 10792
rect 2464 10752 2470 10764
rect 2501 10761 2513 10764
rect 2547 10761 2559 10795
rect 4246 10792 4252 10804
rect 2501 10755 2559 10761
rect 3252 10764 4252 10792
rect 1302 10616 1308 10668
rect 1360 10656 1366 10668
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 1360 10628 1593 10656
rect 1360 10616 1366 10628
rect 1581 10625 1593 10628
rect 1627 10656 1639 10659
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 1627 10628 2881 10656
rect 1627 10625 1639 10628
rect 1581 10619 1639 10625
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 1486 10588 1492 10600
rect 1447 10560 1492 10588
rect 1486 10548 1492 10560
rect 1544 10548 1550 10600
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 3252 10597 3280 10764
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 4525 10795 4583 10801
rect 4525 10761 4537 10795
rect 4571 10792 4583 10795
rect 5077 10795 5135 10801
rect 5077 10792 5089 10795
rect 4571 10764 5089 10792
rect 4571 10761 4583 10764
rect 4525 10755 4583 10761
rect 5077 10761 5089 10764
rect 5123 10792 5135 10795
rect 5442 10792 5448 10804
rect 5123 10764 5448 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 6273 10795 6331 10801
rect 6273 10761 6285 10795
rect 6319 10792 6331 10795
rect 6914 10792 6920 10804
rect 6319 10764 6920 10792
rect 6319 10761 6331 10764
rect 6273 10755 6331 10761
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 8202 10792 8208 10804
rect 8163 10764 8208 10792
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 8570 10792 8576 10804
rect 8531 10764 8576 10792
rect 8570 10752 8576 10764
rect 8628 10752 8634 10804
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 11388 10764 11805 10792
rect 11388 10752 11394 10764
rect 11793 10761 11805 10764
rect 11839 10761 11851 10795
rect 14366 10792 14372 10804
rect 14327 10764 14372 10792
rect 11793 10755 11851 10761
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 15930 10792 15936 10804
rect 15891 10764 15936 10792
rect 15930 10752 15936 10764
rect 15988 10752 15994 10804
rect 16853 10795 16911 10801
rect 16853 10761 16865 10795
rect 16899 10792 16911 10795
rect 16942 10792 16948 10804
rect 16899 10764 16948 10792
rect 16899 10761 16911 10764
rect 16853 10755 16911 10761
rect 16942 10752 16948 10764
rect 17000 10752 17006 10804
rect 18690 10752 18696 10804
rect 18748 10792 18754 10804
rect 19429 10795 19487 10801
rect 19429 10792 19441 10795
rect 18748 10764 19441 10792
rect 18748 10752 18754 10764
rect 19429 10761 19441 10764
rect 19475 10761 19487 10795
rect 19794 10792 19800 10804
rect 19755 10764 19800 10792
rect 19429 10755 19487 10761
rect 19794 10752 19800 10764
rect 19852 10752 19858 10804
rect 21358 10792 21364 10804
rect 21319 10764 21364 10792
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 24670 10792 24676 10804
rect 24631 10764 24676 10792
rect 24670 10752 24676 10764
rect 24728 10752 24734 10804
rect 4706 10724 4712 10736
rect 4667 10696 4712 10724
rect 4706 10684 4712 10696
rect 4764 10684 4770 10736
rect 5813 10727 5871 10733
rect 5813 10693 5825 10727
rect 5859 10724 5871 10727
rect 7558 10724 7564 10736
rect 5859 10696 7564 10724
rect 5859 10693 5871 10696
rect 5813 10687 5871 10693
rect 7558 10684 7564 10696
rect 7616 10684 7622 10736
rect 7650 10684 7656 10736
rect 7708 10724 7714 10736
rect 13633 10727 13691 10733
rect 13633 10724 13645 10727
rect 7708 10696 13645 10724
rect 7708 10684 7714 10696
rect 13633 10693 13645 10696
rect 13679 10724 13691 10727
rect 14182 10724 14188 10736
rect 13679 10696 14188 10724
rect 13679 10693 13691 10696
rect 13633 10687 13691 10693
rect 14182 10684 14188 10696
rect 14240 10684 14246 10736
rect 19058 10724 19064 10736
rect 19019 10696 19064 10724
rect 19058 10684 19064 10696
rect 19116 10684 19122 10736
rect 3694 10656 3700 10668
rect 3655 10628 3700 10656
rect 3694 10616 3700 10628
rect 3752 10616 3758 10668
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3936 10628 3985 10656
rect 3936 10616 3942 10628
rect 3973 10625 3985 10628
rect 4019 10656 4031 10659
rect 6641 10659 6699 10665
rect 4019 10628 5120 10656
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1728 10560 1777 10588
rect 1728 10548 1734 10560
rect 1765 10557 1777 10560
rect 1811 10588 1823 10591
rect 3237 10591 3295 10597
rect 3237 10588 3249 10591
rect 1811 10560 3249 10588
rect 1811 10557 1823 10560
rect 1765 10551 1823 10557
rect 3237 10557 3249 10560
rect 3283 10557 3295 10591
rect 3237 10551 3295 10557
rect 2225 10523 2283 10529
rect 2225 10489 2237 10523
rect 2271 10520 2283 10523
rect 3418 10520 3424 10532
rect 2271 10492 3424 10520
rect 2271 10489 2283 10492
rect 2225 10483 2283 10489
rect 3418 10480 3424 10492
rect 3476 10480 3482 10532
rect 3694 10480 3700 10532
rect 3752 10520 3758 10532
rect 3789 10523 3847 10529
rect 3789 10520 3801 10523
rect 3752 10492 3801 10520
rect 3752 10480 3758 10492
rect 3789 10489 3801 10492
rect 3835 10489 3847 10523
rect 5092 10520 5120 10628
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 6825 10659 6883 10665
rect 6825 10656 6837 10659
rect 6687 10628 6837 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 6825 10625 6837 10628
rect 6871 10656 6883 10659
rect 7006 10656 7012 10668
rect 6871 10628 7012 10656
rect 6871 10625 6883 10628
rect 6825 10619 6883 10625
rect 7006 10616 7012 10628
rect 7064 10616 7070 10668
rect 11514 10656 11520 10668
rect 11475 10628 11520 10656
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10656 12587 10659
rect 12710 10656 12716 10668
rect 12575 10628 12716 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 14826 10656 14832 10668
rect 13786 10628 14832 10656
rect 5994 10548 6000 10600
rect 6052 10588 6058 10600
rect 6917 10591 6975 10597
rect 6917 10588 6929 10591
rect 6052 10560 6929 10588
rect 6052 10548 6058 10560
rect 6917 10557 6929 10560
rect 6963 10588 6975 10591
rect 7098 10588 7104 10600
rect 6963 10560 7104 10588
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 8941 10591 8999 10597
rect 8941 10557 8953 10591
rect 8987 10557 8999 10591
rect 8941 10551 8999 10557
rect 5258 10520 5264 10532
rect 5092 10492 5264 10520
rect 3789 10483 3847 10489
rect 5258 10480 5264 10492
rect 5316 10480 5322 10532
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 8956 10520 8984 10551
rect 9122 10548 9128 10600
rect 9180 10588 9186 10600
rect 9401 10591 9459 10597
rect 9401 10588 9413 10591
rect 9180 10560 9413 10588
rect 9180 10548 9186 10560
rect 9401 10557 9413 10560
rect 9447 10588 9459 10591
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 9447 10560 10333 10588
rect 9447 10557 9459 10560
rect 9401 10551 9459 10557
rect 10321 10557 10333 10560
rect 10367 10588 10379 10591
rect 10410 10588 10416 10600
rect 10367 10560 10416 10588
rect 10367 10557 10379 10560
rect 10321 10551 10379 10557
rect 10410 10548 10416 10560
rect 10468 10548 10474 10600
rect 11330 10588 11336 10600
rect 11291 10560 11336 10588
rect 11330 10548 11336 10560
rect 11388 10548 11394 10600
rect 13173 10591 13231 10597
rect 13173 10557 13185 10591
rect 13219 10588 13231 10591
rect 13262 10588 13268 10600
rect 13219 10560 13268 10588
rect 13219 10557 13231 10560
rect 13173 10551 13231 10557
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 9030 10520 9036 10532
rect 5408 10492 5453 10520
rect 6840 10492 9036 10520
rect 5408 10480 5414 10492
rect 3510 10412 3516 10464
rect 3568 10452 3574 10464
rect 4525 10455 4583 10461
rect 4525 10452 4537 10455
rect 3568 10424 4537 10452
rect 3568 10412 3574 10424
rect 4525 10421 4537 10424
rect 4571 10421 4583 10455
rect 4525 10415 4583 10421
rect 4614 10412 4620 10464
rect 4672 10452 4678 10464
rect 6840 10452 6868 10492
rect 9030 10480 9036 10492
rect 9088 10480 9094 10532
rect 9674 10520 9680 10532
rect 9635 10492 9680 10520
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 12621 10523 12679 10529
rect 12621 10489 12633 10523
rect 12667 10489 12679 10523
rect 13786 10520 13814 10628
rect 14826 10616 14832 10628
rect 14884 10656 14890 10668
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 14884 10628 15025 10656
rect 14884 10616 14890 10628
rect 15013 10625 15025 10628
rect 15059 10625 15071 10659
rect 15654 10656 15660 10668
rect 15615 10628 15660 10656
rect 15013 10619 15071 10625
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 17788 10628 18153 10656
rect 12621 10483 12679 10489
rect 13280 10492 13814 10520
rect 14829 10523 14887 10529
rect 4672 10424 6868 10452
rect 4672 10412 4678 10424
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 9950 10452 9956 10464
rect 7064 10424 9956 10452
rect 7064 10412 7070 10424
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 11974 10412 11980 10464
rect 12032 10452 12038 10464
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 12032 10424 12173 10452
rect 12032 10412 12038 10424
rect 12161 10421 12173 10424
rect 12207 10452 12219 10455
rect 12636 10452 12664 10483
rect 12207 10424 12664 10452
rect 12207 10421 12219 10424
rect 12161 10415 12219 10421
rect 12802 10412 12808 10464
rect 12860 10452 12866 10464
rect 13280 10452 13308 10492
rect 14829 10489 14841 10523
rect 14875 10520 14887 10523
rect 15105 10523 15163 10529
rect 15105 10520 15117 10523
rect 14875 10492 15117 10520
rect 14875 10489 14887 10492
rect 14829 10483 14887 10489
rect 15105 10489 15117 10492
rect 15151 10520 15163 10523
rect 16206 10520 16212 10532
rect 15151 10492 16212 10520
rect 15151 10489 15163 10492
rect 15105 10483 15163 10489
rect 16206 10480 16212 10492
rect 16264 10480 16270 10532
rect 17788 10529 17816 10628
rect 18141 10625 18153 10628
rect 18187 10625 18199 10659
rect 18414 10656 18420 10668
rect 18375 10628 18420 10656
rect 18141 10619 18199 10625
rect 18414 10616 18420 10628
rect 18472 10616 18478 10668
rect 19426 10548 19432 10600
rect 19484 10588 19490 10600
rect 19613 10591 19671 10597
rect 19613 10588 19625 10591
rect 19484 10560 19625 10588
rect 19484 10548 19490 10560
rect 19613 10557 19625 10560
rect 19659 10588 19671 10591
rect 20073 10591 20131 10597
rect 20073 10588 20085 10591
rect 19659 10560 20085 10588
rect 19659 10557 19671 10560
rect 19613 10551 19671 10557
rect 20073 10557 20085 10560
rect 20119 10557 20131 10591
rect 20073 10551 20131 10557
rect 16945 10523 17003 10529
rect 16945 10489 16957 10523
rect 16991 10520 17003 10523
rect 17773 10523 17831 10529
rect 17773 10520 17785 10523
rect 16991 10492 17785 10520
rect 16991 10489 17003 10492
rect 16945 10483 17003 10489
rect 17773 10489 17785 10492
rect 17819 10489 17831 10523
rect 18230 10520 18236 10532
rect 18191 10492 18236 10520
rect 17773 10483 17831 10489
rect 18230 10480 18236 10492
rect 18288 10480 18294 10532
rect 13998 10452 14004 10464
rect 12860 10424 13308 10452
rect 13959 10424 14004 10452
rect 12860 10412 12866 10424
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 17497 10455 17555 10461
rect 17497 10421 17509 10455
rect 17543 10452 17555 10455
rect 17954 10452 17960 10464
rect 17543 10424 17960 10452
rect 17543 10421 17555 10424
rect 17497 10415 17555 10421
rect 17954 10412 17960 10424
rect 18012 10412 18018 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 2409 10251 2467 10257
rect 2409 10248 2421 10251
rect 1544 10220 2421 10248
rect 1544 10208 1550 10220
rect 2409 10217 2421 10220
rect 2455 10217 2467 10251
rect 2774 10248 2780 10260
rect 2735 10220 2780 10248
rect 2409 10211 2467 10217
rect 2774 10208 2780 10220
rect 2832 10208 2838 10260
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 3418 10248 3424 10260
rect 3379 10220 3424 10248
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 4249 10251 4307 10257
rect 4249 10217 4261 10251
rect 4295 10248 4307 10251
rect 4430 10248 4436 10260
rect 4295 10220 4436 10248
rect 4295 10217 4307 10220
rect 4249 10211 4307 10217
rect 4430 10208 4436 10220
rect 4488 10208 4494 10260
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 5350 10248 5356 10260
rect 4663 10220 5356 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 6086 10248 6092 10260
rect 6047 10220 6092 10248
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 7098 10248 7104 10260
rect 7059 10220 7104 10248
rect 7098 10208 7104 10220
rect 7156 10208 7162 10260
rect 9030 10248 9036 10260
rect 8991 10220 9036 10248
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 9861 10251 9919 10257
rect 9861 10248 9873 10251
rect 9732 10220 9873 10248
rect 9732 10208 9738 10220
rect 9861 10217 9873 10220
rect 9907 10217 9919 10251
rect 9861 10211 9919 10217
rect 11330 10208 11336 10260
rect 11388 10248 11394 10260
rect 11425 10251 11483 10257
rect 11425 10248 11437 10251
rect 11388 10220 11437 10248
rect 11388 10208 11394 10220
rect 11425 10217 11437 10220
rect 11471 10217 11483 10251
rect 11790 10248 11796 10260
rect 11751 10220 11796 10248
rect 11425 10211 11483 10217
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 13906 10248 13912 10260
rect 13867 10220 13912 10248
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 15930 10248 15936 10260
rect 15891 10220 15936 10248
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 16485 10251 16543 10257
rect 16485 10217 16497 10251
rect 16531 10248 16543 10251
rect 16850 10248 16856 10260
rect 16531 10220 16856 10248
rect 16531 10217 16543 10220
rect 16485 10211 16543 10217
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 17126 10248 17132 10260
rect 17087 10220 17132 10248
rect 17126 10208 17132 10220
rect 17184 10208 17190 10260
rect 17678 10248 17684 10260
rect 17639 10220 17684 10248
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 18012 10220 18245 10248
rect 18012 10208 18018 10220
rect 18233 10217 18245 10220
rect 18279 10248 18291 10251
rect 18322 10248 18328 10260
rect 18279 10220 18328 10248
rect 18279 10217 18291 10220
rect 18233 10211 18291 10217
rect 18322 10208 18328 10220
rect 18380 10248 18386 10260
rect 19058 10248 19064 10260
rect 18380 10220 19064 10248
rect 18380 10208 18386 10220
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 2133 10183 2191 10189
rect 2133 10149 2145 10183
rect 2179 10180 2191 10183
rect 2222 10180 2228 10192
rect 2179 10152 2228 10180
rect 2179 10149 2191 10152
rect 2133 10143 2191 10149
rect 2222 10140 2228 10152
rect 2280 10140 2286 10192
rect 4982 10180 4988 10192
rect 2976 10152 4988 10180
rect 1302 10072 1308 10124
rect 1360 10112 1366 10124
rect 1489 10115 1547 10121
rect 1489 10112 1501 10115
rect 1360 10084 1501 10112
rect 1360 10072 1366 10084
rect 1489 10081 1501 10084
rect 1535 10081 1547 10115
rect 1489 10075 1547 10081
rect 2866 10072 2872 10124
rect 2924 10112 2930 10124
rect 2976 10121 3004 10152
rect 4982 10140 4988 10152
rect 5040 10140 5046 10192
rect 5258 10140 5264 10192
rect 5316 10180 5322 10192
rect 6457 10183 6515 10189
rect 6457 10180 6469 10183
rect 5316 10152 6469 10180
rect 5316 10140 5322 10152
rect 6457 10149 6469 10152
rect 6503 10149 6515 10183
rect 8294 10180 8300 10192
rect 6457 10143 6515 10149
rect 8128 10152 8300 10180
rect 8128 10124 8156 10152
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 8386 10140 8392 10192
rect 8444 10180 8450 10192
rect 10229 10183 10287 10189
rect 10229 10180 10241 10183
rect 8444 10152 10241 10180
rect 8444 10140 8450 10152
rect 10229 10149 10241 10152
rect 10275 10180 10287 10183
rect 10505 10183 10563 10189
rect 10505 10180 10517 10183
rect 10275 10152 10517 10180
rect 10275 10149 10287 10152
rect 10229 10143 10287 10149
rect 10505 10149 10517 10152
rect 10551 10149 10563 10183
rect 10505 10143 10563 10149
rect 10597 10183 10655 10189
rect 10597 10149 10609 10183
rect 10643 10180 10655 10183
rect 10962 10180 10968 10192
rect 10643 10152 10968 10180
rect 10643 10149 10655 10152
rect 10597 10143 10655 10149
rect 10962 10140 10968 10152
rect 11020 10140 11026 10192
rect 12161 10183 12219 10189
rect 12161 10149 12173 10183
rect 12207 10180 12219 10183
rect 12342 10180 12348 10192
rect 12207 10152 12348 10180
rect 12207 10149 12219 10152
rect 12161 10143 12219 10149
rect 12342 10140 12348 10152
rect 12400 10140 12406 10192
rect 14274 10180 14280 10192
rect 13924 10152 14280 10180
rect 2961 10115 3019 10121
rect 2961 10112 2973 10115
rect 2924 10084 2973 10112
rect 2924 10072 2930 10084
rect 2961 10081 2973 10084
rect 3007 10081 3019 10115
rect 4062 10112 4068 10124
rect 4023 10084 4068 10112
rect 2961 10075 3019 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 5074 10112 5080 10124
rect 5035 10084 5080 10112
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10081 5411 10115
rect 5353 10075 5411 10081
rect 5813 10115 5871 10121
rect 5813 10081 5825 10115
rect 5859 10112 5871 10115
rect 6641 10115 6699 10121
rect 6641 10112 6653 10115
rect 5859 10084 6653 10112
rect 5859 10081 5871 10084
rect 5813 10075 5871 10081
rect 6641 10081 6653 10084
rect 6687 10112 6699 10115
rect 7098 10112 7104 10124
rect 6687 10084 7104 10112
rect 6687 10081 6699 10084
rect 6641 10075 6699 10081
rect 4982 10004 4988 10056
rect 5040 10044 5046 10056
rect 5368 10044 5396 10075
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 8110 10112 8116 10124
rect 8023 10084 8116 10112
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 8481 10115 8539 10121
rect 8481 10112 8493 10115
rect 8260 10084 8493 10112
rect 8260 10072 8266 10084
rect 8481 10081 8493 10084
rect 8527 10081 8539 10115
rect 8481 10075 8539 10081
rect 13722 10072 13728 10124
rect 13780 10112 13786 10124
rect 13924 10121 13952 10152
rect 14274 10140 14280 10152
rect 14332 10140 14338 10192
rect 18690 10140 18696 10192
rect 18748 10180 18754 10192
rect 19199 10183 19257 10189
rect 19199 10180 19211 10183
rect 18748 10152 19211 10180
rect 18748 10140 18754 10152
rect 19199 10149 19211 10152
rect 19245 10149 19257 10183
rect 19199 10143 19257 10149
rect 13909 10115 13967 10121
rect 13909 10112 13921 10115
rect 13780 10084 13921 10112
rect 13780 10072 13786 10084
rect 13909 10081 13921 10084
rect 13955 10081 13967 10115
rect 13909 10075 13967 10081
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 14056 10084 14105 10112
rect 14056 10072 14062 10084
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 19112 10115 19170 10121
rect 19112 10081 19124 10115
rect 19158 10112 19170 10115
rect 19158 10081 19196 10112
rect 19112 10075 19196 10081
rect 5040 10016 5396 10044
rect 8757 10047 8815 10053
rect 5040 10004 5046 10016
rect 8757 10013 8769 10047
rect 8803 10044 8815 10047
rect 10134 10044 10140 10056
rect 8803 10016 10140 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 12066 10044 12072 10056
rect 12027 10016 12072 10044
rect 12066 10004 12072 10016
rect 12124 10004 12130 10056
rect 12710 10044 12716 10056
rect 12671 10016 12716 10044
rect 12710 10004 12716 10016
rect 12768 10004 12774 10056
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 15565 10047 15623 10053
rect 15565 10044 15577 10047
rect 15436 10016 15577 10044
rect 15436 10004 15442 10016
rect 15565 10013 15577 10016
rect 15611 10013 15623 10047
rect 17310 10044 17316 10056
rect 17271 10016 17316 10044
rect 15565 10007 15623 10013
rect 17310 10004 17316 10016
rect 17368 10004 17374 10056
rect 19168 10044 19196 10075
rect 19242 10044 19248 10056
rect 19168 10016 19248 10044
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 3881 9979 3939 9985
rect 3881 9945 3893 9979
rect 3927 9976 3939 9979
rect 3970 9976 3976 9988
rect 3927 9948 3976 9976
rect 3927 9945 3939 9948
rect 3881 9939 3939 9945
rect 3970 9936 3976 9948
rect 4028 9976 4034 9988
rect 4154 9976 4160 9988
rect 4028 9948 4160 9976
rect 4028 9936 4034 9948
rect 4154 9936 4160 9948
rect 4212 9936 4218 9988
rect 5169 9979 5227 9985
rect 5169 9945 5181 9979
rect 5215 9976 5227 9979
rect 5258 9976 5264 9988
rect 5215 9948 5264 9976
rect 5215 9945 5227 9948
rect 5169 9939 5227 9945
rect 5258 9936 5264 9948
rect 5316 9936 5322 9988
rect 11057 9979 11115 9985
rect 11057 9945 11069 9979
rect 11103 9976 11115 9979
rect 12728 9976 12756 10004
rect 11103 9948 12756 9976
rect 11103 9945 11115 9948
rect 11057 9939 11115 9945
rect 4985 9911 5043 9917
rect 4985 9877 4997 9911
rect 5031 9908 5043 9911
rect 5534 9908 5540 9920
rect 5031 9880 5540 9908
rect 5031 9877 5043 9880
rect 4985 9871 5043 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 6730 9868 6736 9920
rect 6788 9908 6794 9920
rect 6825 9911 6883 9917
rect 6825 9908 6837 9911
rect 6788 9880 6837 9908
rect 6788 9868 6794 9880
rect 6825 9877 6837 9880
rect 6871 9908 6883 9911
rect 7650 9908 7656 9920
rect 6871 9880 7656 9908
rect 6871 9877 6883 9880
rect 6825 9871 6883 9877
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 7834 9908 7840 9920
rect 7795 9880 7840 9908
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 13354 9868 13360 9920
rect 13412 9908 13418 9920
rect 14645 9911 14703 9917
rect 14645 9908 14657 9911
rect 13412 9880 14657 9908
rect 13412 9868 13418 9880
rect 14645 9877 14657 9880
rect 14691 9877 14703 9911
rect 14645 9871 14703 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 2406 9704 2412 9716
rect 2367 9676 2412 9704
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 8202 9664 8208 9716
rect 8260 9704 8266 9716
rect 8260 9676 8845 9704
rect 8260 9664 8266 9676
rect 2777 9639 2835 9645
rect 2777 9636 2789 9639
rect 1504 9608 2789 9636
rect 1302 9528 1308 9580
rect 1360 9568 1366 9580
rect 1504 9577 1532 9608
rect 2777 9605 2789 9608
rect 2823 9636 2835 9639
rect 3145 9639 3203 9645
rect 3145 9636 3157 9639
rect 2823 9608 3157 9636
rect 2823 9605 2835 9608
rect 2777 9599 2835 9605
rect 3145 9605 3157 9608
rect 3191 9605 3203 9639
rect 6730 9636 6736 9648
rect 3145 9599 3203 9605
rect 4126 9608 6736 9636
rect 1489 9571 1547 9577
rect 1489 9568 1501 9571
rect 1360 9540 1501 9568
rect 1360 9528 1366 9540
rect 1489 9537 1501 9540
rect 1535 9537 1547 9571
rect 1854 9568 1860 9580
rect 1815 9540 1860 9568
rect 1489 9531 1547 9537
rect 1854 9528 1860 9540
rect 1912 9528 1918 9580
rect 4126 9568 4154 9608
rect 6730 9596 6736 9608
rect 6788 9596 6794 9648
rect 7009 9639 7067 9645
rect 7009 9605 7021 9639
rect 7055 9636 7067 9639
rect 8294 9636 8300 9648
rect 7055 9608 8300 9636
rect 7055 9605 7067 9608
rect 7009 9599 7067 9605
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 8817 9636 8845 9676
rect 8938 9664 8944 9716
rect 8996 9704 9002 9716
rect 11241 9707 11299 9713
rect 11241 9704 11253 9707
rect 8996 9676 11253 9704
rect 8996 9664 9002 9676
rect 11241 9673 11253 9676
rect 11287 9704 11299 9707
rect 12066 9704 12072 9716
rect 11287 9676 12072 9704
rect 11287 9673 11299 9676
rect 11241 9667 11299 9673
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 13722 9704 13728 9716
rect 13683 9676 13728 9704
rect 13722 9664 13728 9676
rect 13780 9664 13786 9716
rect 13906 9664 13912 9716
rect 13964 9704 13970 9716
rect 15289 9707 15347 9713
rect 15289 9704 15301 9707
rect 13964 9676 15301 9704
rect 13964 9664 13970 9676
rect 15289 9673 15301 9676
rect 15335 9704 15347 9707
rect 15565 9707 15623 9713
rect 15565 9704 15577 9707
rect 15335 9676 15577 9704
rect 15335 9673 15347 9676
rect 15289 9667 15347 9673
rect 15565 9673 15577 9676
rect 15611 9704 15623 9707
rect 15930 9704 15936 9716
rect 15611 9676 15936 9704
rect 15611 9673 15623 9676
rect 15565 9667 15623 9673
rect 15930 9664 15936 9676
rect 15988 9664 15994 9716
rect 17865 9707 17923 9713
rect 17865 9673 17877 9707
rect 17911 9704 17923 9707
rect 18322 9704 18328 9716
rect 17911 9676 18328 9704
rect 17911 9673 17923 9676
rect 17865 9667 17923 9673
rect 18322 9664 18328 9676
rect 18380 9664 18386 9716
rect 19242 9704 19248 9716
rect 19203 9676 19248 9704
rect 19242 9664 19248 9676
rect 19300 9664 19306 9716
rect 9122 9636 9128 9648
rect 8817 9608 9128 9636
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 3896 9540 4154 9568
rect 4341 9571 4399 9577
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 2406 9500 2412 9512
rect 1719 9472 2412 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 3896 9509 3924 9540
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 7834 9568 7840 9580
rect 4387 9540 7840 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 7834 9528 7840 9540
rect 7892 9568 7898 9580
rect 7929 9571 7987 9577
rect 7929 9568 7941 9571
rect 7892 9540 7941 9568
rect 7892 9528 7898 9540
rect 7929 9537 7941 9540
rect 7975 9537 7987 9571
rect 9401 9571 9459 9577
rect 9401 9568 9413 9571
rect 7929 9531 7987 9537
rect 8404 9540 9413 9568
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3752 9472 3893 9500
rect 3752 9460 3758 9472
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 4065 9503 4123 9509
rect 4065 9500 4077 9503
rect 4028 9472 4077 9500
rect 4028 9460 4034 9472
rect 4065 9469 4077 9472
rect 4111 9469 4123 9503
rect 4065 9463 4123 9469
rect 4709 9503 4767 9509
rect 4709 9469 4721 9503
rect 4755 9500 4767 9503
rect 4982 9500 4988 9512
rect 4755 9472 4988 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5169 9503 5227 9509
rect 5169 9469 5181 9503
rect 5215 9469 5227 9503
rect 5169 9463 5227 9469
rect 5184 9432 5212 9463
rect 5258 9460 5264 9512
rect 5316 9500 5322 9512
rect 5445 9503 5503 9509
rect 5316 9472 5361 9500
rect 5316 9460 5322 9472
rect 5445 9469 5457 9503
rect 5491 9500 5503 9503
rect 5994 9500 6000 9512
rect 5491 9472 6000 9500
rect 5491 9469 5503 9472
rect 5445 9463 5503 9469
rect 5994 9460 6000 9472
rect 6052 9500 6058 9512
rect 6549 9503 6607 9509
rect 6549 9500 6561 9503
rect 6052 9472 6561 9500
rect 6052 9460 6058 9472
rect 6549 9469 6561 9472
rect 6595 9469 6607 9503
rect 6549 9463 6607 9469
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 6871 9472 7328 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 5534 9432 5540 9444
rect 5184 9404 5540 9432
rect 5534 9392 5540 9404
rect 5592 9392 5598 9444
rect 5905 9435 5963 9441
rect 5905 9401 5917 9435
rect 5951 9432 5963 9435
rect 6730 9432 6736 9444
rect 5951 9404 6736 9432
rect 5951 9401 5963 9404
rect 5905 9395 5963 9401
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 7300 9376 7328 9472
rect 8404 9444 8432 9540
rect 9401 9537 9413 9540
rect 9447 9568 9459 9571
rect 9493 9571 9551 9577
rect 9493 9568 9505 9571
rect 9447 9540 9505 9568
rect 9447 9537 9459 9540
rect 9401 9531 9459 9537
rect 9493 9537 9505 9540
rect 9539 9537 9551 9571
rect 9674 9568 9680 9580
rect 9635 9540 9680 9568
rect 9493 9531 9551 9537
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 13262 9528 13268 9580
rect 13320 9568 13326 9580
rect 14369 9571 14427 9577
rect 14369 9568 14381 9571
rect 13320 9540 14381 9568
rect 13320 9528 13326 9540
rect 14369 9537 14381 9540
rect 14415 9537 14427 9571
rect 15948 9568 15976 9664
rect 15948 9540 16297 9568
rect 14369 9531 14427 9537
rect 11977 9503 12035 9509
rect 11977 9500 11989 9503
rect 8864 9472 11989 9500
rect 7742 9432 7748 9444
rect 7703 9404 7748 9432
rect 7742 9392 7748 9404
rect 7800 9432 7806 9444
rect 8250 9435 8308 9441
rect 8250 9432 8262 9435
rect 7800 9404 8262 9432
rect 7800 9392 7806 9404
rect 8250 9401 8262 9404
rect 8296 9432 8308 9435
rect 8386 9432 8392 9444
rect 8296 9404 8392 9432
rect 8296 9401 8308 9404
rect 8250 9395 8308 9401
rect 8386 9392 8392 9404
rect 8444 9392 8450 9444
rect 8864 9376 8892 9472
rect 11977 9469 11989 9472
rect 12023 9500 12035 9503
rect 12342 9500 12348 9512
rect 12023 9472 12348 9500
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 15930 9500 15936 9512
rect 15891 9472 15936 9500
rect 15930 9460 15936 9472
rect 15988 9460 15994 9512
rect 16269 9500 16297 9540
rect 17218 9528 17224 9580
rect 17276 9568 17282 9580
rect 18506 9568 18512 9580
rect 17276 9540 18512 9568
rect 17276 9528 17282 9540
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 17313 9503 17371 9509
rect 17313 9500 17325 9503
rect 16269 9472 17325 9500
rect 10042 9441 10048 9444
rect 9401 9435 9459 9441
rect 9401 9401 9413 9435
rect 9447 9432 9459 9435
rect 9998 9435 10048 9441
rect 9998 9432 10010 9435
rect 9447 9404 10010 9432
rect 9447 9401 9459 9404
rect 9401 9395 9459 9401
rect 9998 9401 10010 9404
rect 10044 9401 10048 9435
rect 9998 9395 10048 9401
rect 10042 9392 10048 9395
rect 10100 9392 10106 9444
rect 11701 9435 11759 9441
rect 11701 9401 11713 9435
rect 11747 9432 11759 9435
rect 12529 9435 12587 9441
rect 12529 9432 12541 9435
rect 11747 9404 12541 9432
rect 11747 9401 11759 9404
rect 11701 9395 11759 9401
rect 12529 9401 12541 9404
rect 12575 9401 12587 9435
rect 12529 9395 12587 9401
rect 4522 9324 4528 9376
rect 4580 9364 4586 9376
rect 4985 9367 5043 9373
rect 4985 9364 4997 9367
rect 4580 9336 4997 9364
rect 4580 9324 4586 9336
rect 4985 9333 4997 9336
rect 5031 9364 5043 9367
rect 5074 9364 5080 9376
rect 5031 9336 5080 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 6178 9364 6184 9376
rect 6139 9336 6184 9364
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 7282 9364 7288 9376
rect 7243 9336 7288 9364
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 8846 9364 8852 9376
rect 8807 9336 8852 9364
rect 8846 9324 8852 9336
rect 8904 9324 8910 9376
rect 10597 9367 10655 9373
rect 10597 9333 10609 9367
rect 10643 9364 10655 9367
rect 10962 9364 10968 9376
rect 10643 9336 10968 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12544 9364 12572 9395
rect 12618 9392 12624 9444
rect 12676 9432 12682 9444
rect 13173 9435 13231 9441
rect 12676 9404 12721 9432
rect 12676 9392 12682 9404
rect 13173 9401 13185 9435
rect 13219 9432 13231 9435
rect 13354 9432 13360 9444
rect 13219 9404 13360 9432
rect 13219 9401 13231 9404
rect 13173 9395 13231 9401
rect 13354 9392 13360 9404
rect 13412 9432 13418 9444
rect 14093 9435 14151 9441
rect 14093 9432 14105 9435
rect 13412 9404 14105 9432
rect 13412 9392 13418 9404
rect 14093 9401 14105 9404
rect 14139 9401 14151 9435
rect 14093 9395 14151 9401
rect 14182 9392 14188 9444
rect 14240 9432 14246 9444
rect 16269 9441 16297 9472
rect 17313 9469 17325 9472
rect 17359 9500 17371 9503
rect 17678 9500 17684 9512
rect 17359 9472 17684 9500
rect 17359 9469 17371 9472
rect 17313 9463 17371 9469
rect 17678 9460 17684 9472
rect 17736 9460 17742 9512
rect 16254 9435 16312 9441
rect 14240 9404 14285 9432
rect 14240 9392 14246 9404
rect 16254 9401 16266 9435
rect 16300 9401 16312 9435
rect 18230 9432 18236 9444
rect 18191 9404 18236 9432
rect 16254 9395 16312 9401
rect 18230 9392 18236 9404
rect 18288 9392 18294 9444
rect 18322 9392 18328 9444
rect 18380 9432 18386 9444
rect 18380 9404 18425 9432
rect 18380 9392 18386 9404
rect 16850 9364 16856 9376
rect 12492 9336 12572 9364
rect 16811 9336 16856 9364
rect 12492 9324 12498 9336
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2866 9160 2872 9172
rect 2827 9132 2872 9160
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 3145 9163 3203 9169
rect 3145 9129 3157 9163
rect 3191 9160 3203 9163
rect 3326 9160 3332 9172
rect 3191 9132 3332 9160
rect 3191 9129 3203 9132
rect 3145 9123 3203 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 3694 9160 3700 9172
rect 3655 9132 3700 9160
rect 3694 9120 3700 9132
rect 3752 9120 3758 9172
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 6638 9160 6644 9172
rect 4120 9132 4384 9160
rect 4120 9120 4126 9132
rect 1394 9092 1400 9104
rect 1355 9064 1400 9092
rect 1394 9052 1400 9064
rect 1452 9092 1458 9104
rect 2409 9095 2467 9101
rect 2409 9092 2421 9095
rect 1452 9064 2421 9092
rect 1452 9052 1458 9064
rect 2409 9061 2421 9064
rect 2455 9061 2467 9095
rect 2409 9055 2467 9061
rect 1486 9024 1492 9036
rect 1447 8996 1492 9024
rect 1486 8984 1492 8996
rect 1544 8984 1550 9036
rect 2958 9024 2964 9036
rect 2919 8996 2964 9024
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 4356 8965 4384 9132
rect 5552 9132 6644 9160
rect 5552 9104 5580 9132
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 7098 9160 7104 9172
rect 7059 9132 7104 9160
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 7837 9163 7895 9169
rect 7837 9129 7849 9163
rect 7883 9160 7895 9163
rect 8110 9160 8116 9172
rect 7883 9132 8116 9160
rect 7883 9129 7895 9132
rect 7837 9123 7895 9129
rect 8110 9120 8116 9132
rect 8168 9160 8174 9172
rect 9861 9163 9919 9169
rect 9861 9160 9873 9163
rect 8168 9132 9873 9160
rect 8168 9120 8174 9132
rect 9861 9129 9873 9132
rect 9907 9129 9919 9163
rect 11974 9160 11980 9172
rect 11935 9132 11980 9160
rect 9861 9123 9919 9129
rect 5261 9095 5319 9101
rect 5261 9061 5273 9095
rect 5307 9092 5319 9095
rect 5534 9092 5540 9104
rect 5307 9064 5540 9092
rect 5307 9061 5319 9064
rect 5261 9055 5319 9061
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 5994 9052 6000 9104
rect 6052 9092 6058 9104
rect 6052 9064 6408 9092
rect 6052 9052 6058 9064
rect 4522 8984 4528 9036
rect 4580 9024 4586 9036
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 4580 8996 4629 9024
rect 4580 8984 4586 8996
rect 4617 8993 4629 8996
rect 4663 9024 4675 9027
rect 6086 9024 6092 9036
rect 4663 8996 6092 9024
rect 4663 8993 4675 8996
rect 4617 8987 4675 8993
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6380 9033 6408 9064
rect 7926 9052 7932 9104
rect 7984 9092 7990 9104
rect 8202 9092 8208 9104
rect 7984 9064 8208 9092
rect 7984 9052 7990 9064
rect 8202 9052 8208 9064
rect 8260 9092 8266 9104
rect 8260 9064 8524 9092
rect 8260 9052 8266 9064
rect 6365 9027 6423 9033
rect 6365 8993 6377 9027
rect 6411 8993 6423 9027
rect 8294 9024 8300 9036
rect 8255 8996 8300 9024
rect 6365 8987 6423 8993
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 8496 9033 8524 9064
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 8993 8539 9027
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 8481 8987 8539 8993
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8956 4399 8959
rect 6549 8959 6607 8965
rect 6549 8956 6561 8959
rect 4387 8928 6561 8956
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 6549 8925 6561 8928
rect 6595 8925 6607 8959
rect 8570 8956 8576 8968
rect 8531 8928 8576 8956
rect 6549 8919 6607 8925
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 6178 8888 6184 8900
rect 5552 8860 6184 8888
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 5258 8820 5264 8832
rect 5132 8792 5264 8820
rect 5132 8780 5138 8792
rect 5258 8780 5264 8792
rect 5316 8820 5322 8832
rect 5552 8829 5580 8860
rect 6178 8848 6184 8860
rect 6236 8848 6242 8900
rect 9876 8888 9904 9123
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12342 9120 12348 9172
rect 12400 9160 12406 9172
rect 12437 9163 12495 9169
rect 12437 9160 12449 9163
rect 12400 9132 12449 9160
rect 12400 9120 12406 9132
rect 12437 9129 12449 9132
rect 12483 9160 12495 9163
rect 12618 9160 12624 9172
rect 12483 9132 12624 9160
rect 12483 9129 12495 9132
rect 12437 9123 12495 9129
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 13725 9163 13783 9169
rect 13725 9129 13737 9163
rect 13771 9160 13783 9163
rect 14182 9160 14188 9172
rect 13771 9132 14188 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 14182 9120 14188 9132
rect 14240 9160 14246 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 14240 9132 14381 9160
rect 14240 9120 14246 9132
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 14369 9123 14427 9129
rect 15930 9120 15936 9172
rect 15988 9160 15994 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 15988 9132 16681 9160
rect 15988 9120 15994 9132
rect 16669 9129 16681 9132
rect 16715 9129 16727 9163
rect 16669 9123 16727 9129
rect 18230 9120 18236 9172
rect 18288 9160 18294 9172
rect 18509 9163 18567 9169
rect 18509 9160 18521 9163
rect 18288 9132 18521 9160
rect 18288 9120 18294 9132
rect 18509 9129 18521 9132
rect 18555 9160 18567 9163
rect 18831 9163 18889 9169
rect 18831 9160 18843 9163
rect 18555 9132 18843 9160
rect 18555 9129 18567 9132
rect 18509 9123 18567 9129
rect 18831 9129 18843 9132
rect 18877 9129 18889 9163
rect 18831 9123 18889 9129
rect 10042 9052 10048 9104
rect 10100 9092 10106 9104
rect 11378 9095 11436 9101
rect 11378 9092 11390 9095
rect 10100 9064 11390 9092
rect 10100 9052 10106 9064
rect 11378 9061 11390 9064
rect 11424 9092 11436 9095
rect 11514 9092 11520 9104
rect 11424 9064 11520 9092
rect 11424 9061 11436 9064
rect 11378 9055 11436 9061
rect 11514 9052 11520 9064
rect 11572 9092 11578 9104
rect 13126 9095 13184 9101
rect 13126 9092 13138 9095
rect 11572 9064 13138 9092
rect 11572 9052 11578 9064
rect 13126 9061 13138 9064
rect 13172 9092 13184 9095
rect 13906 9092 13912 9104
rect 13172 9064 13912 9092
rect 13172 9061 13184 9064
rect 13126 9055 13184 9061
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 13998 9052 14004 9104
rect 14056 9092 14062 9104
rect 14093 9095 14151 9101
rect 14093 9092 14105 9095
rect 14056 9064 14105 9092
rect 14056 9052 14062 9064
rect 14093 9061 14105 9064
rect 14139 9092 14151 9095
rect 14139 9064 15884 9092
rect 14139 9061 14151 9064
rect 14093 9055 14151 9061
rect 10134 8984 10140 9036
rect 10192 9024 10198 9036
rect 11057 9027 11115 9033
rect 11057 9024 11069 9027
rect 10192 8996 11069 9024
rect 10192 8984 10198 8996
rect 11057 8993 11069 8996
rect 11103 9024 11115 9027
rect 11238 9024 11244 9036
rect 11103 8996 11244 9024
rect 11103 8993 11115 8996
rect 11057 8987 11115 8993
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 14550 8984 14556 9036
rect 14608 9024 14614 9036
rect 15286 9024 15292 9036
rect 14608 8996 15292 9024
rect 14608 8984 14614 8996
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 15856 9033 15884 9064
rect 16850 9052 16856 9104
rect 16908 9092 16914 9104
rect 17313 9095 17371 9101
rect 17313 9092 17325 9095
rect 16908 9064 17325 9092
rect 16908 9052 16914 9064
rect 17313 9061 17325 9064
rect 17359 9061 17371 9095
rect 17862 9092 17868 9104
rect 17823 9064 17868 9092
rect 17313 9055 17371 9061
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 15841 9027 15899 9033
rect 15841 8993 15853 9027
rect 15887 9024 15899 9027
rect 16298 9024 16304 9036
rect 15887 8996 16304 9024
rect 15887 8993 15899 8996
rect 15841 8987 15899 8993
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 18693 9027 18751 9033
rect 18693 8993 18705 9027
rect 18739 9024 18751 9027
rect 18782 9024 18788 9036
rect 18739 8996 18788 9024
rect 18739 8993 18751 8996
rect 18693 8987 18751 8993
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 10744 8928 12817 8956
rect 10744 8916 10750 8928
rect 12805 8925 12817 8928
rect 12851 8956 12863 8959
rect 13630 8956 13636 8968
rect 12851 8928 13636 8956
rect 12851 8925 12863 8928
rect 12805 8919 12863 8925
rect 13630 8916 13636 8928
rect 13688 8916 13694 8968
rect 16025 8959 16083 8965
rect 16025 8925 16037 8959
rect 16071 8956 16083 8959
rect 17218 8956 17224 8968
rect 16071 8928 16297 8956
rect 17179 8928 17224 8956
rect 16071 8925 16083 8928
rect 16025 8919 16083 8925
rect 14090 8888 14096 8900
rect 9876 8860 14096 8888
rect 14090 8848 14096 8860
rect 14148 8888 14154 8900
rect 15746 8888 15752 8900
rect 14148 8860 15752 8888
rect 14148 8848 14154 8860
rect 15746 8848 15752 8860
rect 15804 8848 15810 8900
rect 16269 8888 16297 8928
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 18141 8959 18199 8965
rect 18141 8956 18153 8959
rect 17368 8928 18153 8956
rect 17368 8916 17374 8928
rect 18141 8925 18153 8928
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 17328 8888 17356 8916
rect 16269 8860 17356 8888
rect 5537 8823 5595 8829
rect 5537 8820 5549 8823
rect 5316 8792 5549 8820
rect 5316 8780 5322 8792
rect 5537 8789 5549 8792
rect 5583 8789 5595 8823
rect 5994 8820 6000 8832
rect 5955 8792 6000 8820
rect 5537 8783 5595 8789
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 10594 8820 10600 8832
rect 10555 8792 10600 8820
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 10962 8820 10968 8832
rect 10923 8792 10968 8820
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 15105 8823 15163 8829
rect 15105 8789 15117 8823
rect 15151 8820 15163 8823
rect 15378 8820 15384 8832
rect 15151 8792 15384 8820
rect 15151 8789 15163 8792
rect 15105 8783 15163 8789
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15764 8820 15792 8848
rect 16301 8823 16359 8829
rect 16301 8820 16313 8823
rect 15764 8792 16313 8820
rect 16301 8789 16313 8792
rect 16347 8789 16359 8823
rect 16301 8783 16359 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 3050 8576 3056 8628
rect 3108 8616 3114 8628
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 3108 8588 3341 8616
rect 3108 8576 3114 8588
rect 3329 8585 3341 8588
rect 3375 8585 3387 8619
rect 6086 8616 6092 8628
rect 6047 8588 6092 8616
rect 3329 8579 3387 8585
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 7742 8616 7748 8628
rect 6196 8588 7748 8616
rect 4249 8551 4307 8557
rect 4249 8517 4261 8551
rect 4295 8548 4307 8551
rect 6196 8548 6224 8588
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 9769 8619 9827 8625
rect 9769 8616 9781 8619
rect 8352 8588 9781 8616
rect 8352 8576 8358 8588
rect 9769 8585 9781 8588
rect 9815 8616 9827 8619
rect 13538 8616 13544 8628
rect 9815 8588 13544 8616
rect 9815 8585 9827 8588
rect 9769 8579 9827 8585
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 13906 8616 13912 8628
rect 13771 8588 13912 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 15286 8616 15292 8628
rect 15247 8588 15292 8616
rect 15286 8576 15292 8588
rect 15344 8576 15350 8628
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 17129 8619 17187 8625
rect 17129 8616 17141 8619
rect 16908 8588 17141 8616
rect 16908 8576 16914 8588
rect 17129 8585 17141 8588
rect 17175 8585 17187 8619
rect 17129 8579 17187 8585
rect 7837 8551 7895 8557
rect 7837 8548 7849 8551
rect 4295 8520 6224 8548
rect 6932 8520 7849 8548
rect 4295 8517 4307 8520
rect 4249 8511 4307 8517
rect 2958 8440 2964 8492
rect 3016 8480 3022 8492
rect 3053 8483 3111 8489
rect 3053 8480 3065 8483
rect 3016 8452 3065 8480
rect 3016 8440 3022 8452
rect 3053 8449 3065 8452
rect 3099 8480 3111 8483
rect 5350 8480 5356 8492
rect 3099 8452 5356 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 5350 8440 5356 8452
rect 5408 8480 5414 8492
rect 5534 8480 5540 8492
rect 5408 8452 5540 8480
rect 5408 8440 5414 8452
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 5994 8480 6000 8492
rect 5859 8452 6000 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6178 8440 6184 8492
rect 6236 8480 6242 8492
rect 6932 8489 6960 8520
rect 7837 8517 7849 8520
rect 7883 8517 7895 8551
rect 7837 8511 7895 8517
rect 8202 8508 8208 8560
rect 8260 8548 8266 8560
rect 9401 8551 9459 8557
rect 9401 8548 9413 8551
rect 8260 8520 9413 8548
rect 8260 8508 8266 8520
rect 9401 8517 9413 8520
rect 9447 8548 9459 8551
rect 12161 8551 12219 8557
rect 12161 8548 12173 8551
rect 9447 8520 12173 8548
rect 9447 8517 9459 8520
rect 9401 8511 9459 8517
rect 12161 8517 12173 8520
rect 12207 8517 12219 8551
rect 12161 8511 12219 8517
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6236 8452 6929 8480
rect 6236 8440 6242 8452
rect 6917 8449 6929 8452
rect 6963 8449 6975 8483
rect 7282 8480 7288 8492
rect 7243 8452 7288 8480
rect 6917 8443 6975 8449
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 8386 8480 8392 8492
rect 8347 8452 8392 8480
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8480 8539 8483
rect 8570 8480 8576 8492
rect 8527 8452 8576 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 10870 8480 10876 8492
rect 10831 8452 10876 8480
rect 10870 8440 10876 8452
rect 10928 8440 10934 8492
rect 11514 8480 11520 8492
rect 11475 8452 11520 8480
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 4065 8415 4123 8421
rect 4065 8412 4077 8415
rect 3988 8384 4077 8412
rect 3988 8288 4016 8384
rect 4065 8381 4077 8384
rect 4111 8381 4123 8415
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 4065 8375 4123 8381
rect 5000 8384 5181 8412
rect 5000 8288 5028 8384
rect 5169 8381 5181 8384
rect 5215 8412 5227 8415
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 5215 8384 6561 8412
rect 5215 8381 5227 8384
rect 5169 8375 5227 8381
rect 6549 8381 6561 8384
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 6564 8344 6592 8375
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6696 8384 6837 8412
rect 6696 8372 6702 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 7116 8344 7144 8375
rect 8110 8372 8116 8424
rect 8168 8412 8174 8424
rect 9674 8412 9680 8424
rect 8168 8384 9680 8412
rect 8168 8372 8174 8384
rect 9674 8372 9680 8384
rect 9732 8412 9738 8424
rect 10045 8415 10103 8421
rect 10045 8412 10057 8415
rect 9732 8384 10057 8412
rect 9732 8372 9738 8384
rect 10045 8381 10057 8384
rect 10091 8381 10103 8415
rect 12176 8412 12204 8511
rect 12710 8508 12716 8560
rect 12768 8548 12774 8560
rect 12768 8520 14596 8548
rect 12768 8508 12774 8520
rect 14568 8489 14596 8520
rect 17034 8508 17040 8560
rect 17092 8548 17098 8560
rect 18187 8551 18245 8557
rect 18187 8548 18199 8551
rect 17092 8520 18199 8548
rect 17092 8508 17098 8520
rect 18187 8517 18199 8520
rect 18233 8517 18245 8551
rect 18187 8511 18245 8517
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 14553 8443 14611 8449
rect 16316 8452 16865 8480
rect 16316 8424 16344 8452
rect 16853 8449 16865 8452
rect 16899 8480 16911 8483
rect 19334 8480 19340 8492
rect 16899 8452 19340 8480
rect 16899 8449 16911 8452
rect 16853 8443 16911 8449
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 15746 8412 15752 8424
rect 12176 8384 12388 8412
rect 15707 8384 15752 8412
rect 10045 8375 10103 8381
rect 6564 8316 7144 8344
rect 8386 8304 8392 8356
rect 8444 8344 8450 8356
rect 8802 8347 8860 8353
rect 8802 8344 8814 8347
rect 8444 8316 8814 8344
rect 8444 8304 8450 8316
rect 8802 8313 8814 8316
rect 8848 8313 8860 8347
rect 8802 8307 8860 8313
rect 10134 8304 10140 8356
rect 10192 8344 10198 8356
rect 10594 8344 10600 8356
rect 10192 8316 10600 8344
rect 10192 8304 10198 8316
rect 10594 8304 10600 8316
rect 10652 8304 10658 8356
rect 10689 8347 10747 8353
rect 10689 8313 10701 8347
rect 10735 8344 10747 8347
rect 10962 8344 10968 8356
rect 10735 8316 10968 8344
rect 10735 8313 10747 8316
rect 10689 8307 10747 8313
rect 10962 8304 10968 8316
rect 11020 8344 11026 8356
rect 12250 8344 12256 8356
rect 11020 8316 12256 8344
rect 11020 8304 11026 8316
rect 12250 8304 12256 8316
rect 12308 8304 12314 8356
rect 842 8236 848 8288
rect 900 8276 906 8288
rect 1486 8276 1492 8288
rect 900 8248 1492 8276
rect 900 8236 906 8248
rect 1486 8236 1492 8248
rect 1544 8276 1550 8288
rect 1581 8279 1639 8285
rect 1581 8276 1593 8279
rect 1544 8248 1593 8276
rect 1544 8236 1550 8248
rect 1581 8245 1593 8248
rect 1627 8245 1639 8279
rect 3970 8276 3976 8288
rect 3931 8248 3976 8276
rect 1581 8239 1639 8245
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 4522 8276 4528 8288
rect 4483 8248 4528 8276
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 4982 8276 4988 8288
rect 4943 8248 4988 8276
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 12360 8276 12388 8384
rect 15746 8372 15752 8384
rect 15804 8372 15810 8424
rect 16298 8412 16304 8424
rect 16211 8384 16304 8412
rect 16298 8372 16304 8384
rect 16356 8372 16362 8424
rect 17862 8412 17868 8424
rect 17823 8384 17868 8412
rect 17862 8372 17868 8384
rect 17920 8412 17926 8424
rect 18084 8415 18142 8421
rect 18084 8412 18096 8415
rect 17920 8384 18096 8412
rect 17920 8372 17926 8384
rect 18084 8381 18096 8384
rect 18130 8381 18142 8415
rect 18084 8375 18142 8381
rect 12710 8344 12716 8356
rect 12671 8316 12716 8344
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 12805 8347 12863 8353
rect 12805 8313 12817 8347
rect 12851 8313 12863 8347
rect 13354 8344 13360 8356
rect 13315 8316 13360 8344
rect 12805 8307 12863 8313
rect 12820 8276 12848 8307
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 14274 8344 14280 8356
rect 14235 8316 14280 8344
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8313 14427 8347
rect 14369 8307 14427 8313
rect 14001 8279 14059 8285
rect 14001 8276 14013 8279
rect 12360 8248 14013 8276
rect 14001 8245 14013 8248
rect 14047 8276 14059 8279
rect 14384 8276 14412 8307
rect 14047 8248 14412 8276
rect 14047 8245 14059 8248
rect 14001 8239 14059 8245
rect 15930 8236 15936 8288
rect 15988 8276 15994 8288
rect 16025 8279 16083 8285
rect 16025 8276 16037 8279
rect 15988 8248 16037 8276
rect 15988 8236 15994 8248
rect 16025 8245 16037 8248
rect 16071 8245 16083 8279
rect 18782 8276 18788 8288
rect 18743 8248 18788 8276
rect 16025 8239 16083 8245
rect 18782 8236 18788 8248
rect 18840 8236 18846 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 6178 8032 6184 8084
rect 6236 8072 6242 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 6236 8044 6837 8072
rect 6236 8032 6242 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 7926 8072 7932 8084
rect 7887 8044 7932 8072
rect 6825 8035 6883 8041
rect 7926 8032 7932 8044
rect 7984 8032 7990 8084
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 9033 8075 9091 8081
rect 9033 8072 9045 8075
rect 8628 8044 9045 8072
rect 8628 8032 8634 8044
rect 9033 8041 9045 8044
rect 9079 8041 9091 8075
rect 11238 8072 11244 8084
rect 11199 8044 11244 8072
rect 9033 8035 9091 8041
rect 11238 8032 11244 8044
rect 11296 8032 11302 8084
rect 13630 8072 13636 8084
rect 13591 8044 13636 8072
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 15378 8072 15384 8084
rect 15339 8044 15384 8072
rect 15378 8032 15384 8044
rect 15436 8032 15442 8084
rect 16298 8072 16304 8084
rect 16259 8044 16304 8072
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 17218 8072 17224 8084
rect 17179 8044 17224 8072
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 6273 8007 6331 8013
rect 6273 7973 6285 8007
rect 6319 8004 6331 8007
rect 8110 8004 8116 8016
rect 6319 7976 8116 8004
rect 6319 7973 6331 7976
rect 6273 7967 6331 7973
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 8202 7964 8208 8016
rect 8260 8004 8266 8016
rect 8260 7976 8305 8004
rect 8260 7964 8266 7976
rect 10042 7964 10048 8016
rect 10100 8004 10106 8016
rect 10366 8007 10424 8013
rect 10366 8004 10378 8007
rect 10100 7976 10378 8004
rect 10100 7964 10106 7976
rect 10366 7973 10378 7976
rect 10412 7973 10424 8007
rect 10366 7967 10424 7973
rect 12250 7964 12256 8016
rect 12308 8004 12314 8016
rect 12805 8007 12863 8013
rect 12805 8004 12817 8007
rect 12308 7976 12817 8004
rect 12308 7964 12314 7976
rect 12805 7973 12817 7976
rect 12851 7973 12863 8007
rect 13354 8004 13360 8016
rect 13315 7976 13360 8004
rect 12805 7967 12863 7973
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 13814 7964 13820 8016
rect 13872 8004 13878 8016
rect 13872 7976 15608 8004
rect 13872 7964 13878 7976
rect 4522 7936 4528 7948
rect 4483 7908 4528 7936
rect 4522 7896 4528 7908
rect 4580 7936 4586 7948
rect 5442 7936 5448 7948
rect 4580 7908 5448 7936
rect 4580 7896 4586 7908
rect 5442 7896 5448 7908
rect 5500 7936 5506 7948
rect 5537 7939 5595 7945
rect 5537 7936 5549 7939
rect 5500 7908 5549 7936
rect 5500 7896 5506 7908
rect 5537 7905 5549 7908
rect 5583 7905 5595 7939
rect 5537 7899 5595 7905
rect 5813 7939 5871 7945
rect 5813 7905 5825 7939
rect 5859 7905 5871 7939
rect 5813 7899 5871 7905
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 5828 7868 5856 7899
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 6696 7908 7205 7936
rect 6696 7896 6702 7908
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 14182 7936 14188 7948
rect 14143 7908 14188 7936
rect 7193 7899 7251 7905
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 15580 7945 15608 7976
rect 15565 7939 15623 7945
rect 15565 7905 15577 7939
rect 15611 7936 15623 7939
rect 15654 7936 15660 7948
rect 15611 7908 15660 7936
rect 15611 7905 15623 7908
rect 15565 7899 15623 7905
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 15838 7936 15844 7948
rect 15751 7908 15844 7936
rect 15838 7896 15844 7908
rect 15896 7936 15902 7948
rect 16316 7936 16344 8032
rect 15896 7908 16344 7936
rect 15896 7896 15902 7908
rect 8110 7868 8116 7880
rect 5040 7840 5856 7868
rect 8071 7840 8116 7868
rect 5040 7828 5046 7840
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 8754 7868 8760 7880
rect 8715 7840 8760 7868
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 10042 7868 10048 7880
rect 10003 7840 10048 7868
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 12713 7871 12771 7877
rect 12713 7868 12725 7871
rect 11940 7840 12725 7868
rect 11940 7828 11946 7840
rect 12713 7837 12725 7840
rect 12759 7868 12771 7871
rect 14323 7871 14381 7877
rect 14323 7868 14335 7871
rect 12759 7840 14335 7868
rect 12759 7837 12771 7840
rect 12713 7831 12771 7837
rect 14323 7837 14335 7840
rect 14369 7837 14381 7871
rect 14323 7831 14381 7837
rect 5534 7760 5540 7812
rect 5592 7800 5598 7812
rect 5629 7803 5687 7809
rect 5629 7800 5641 7803
rect 5592 7772 5641 7800
rect 5592 7760 5598 7772
rect 5629 7769 5641 7772
rect 5675 7769 5687 7803
rect 5629 7763 5687 7769
rect 4709 7735 4767 7741
rect 4709 7701 4721 7735
rect 4755 7732 4767 7735
rect 6454 7732 6460 7744
rect 4755 7704 6460 7732
rect 4755 7701 4767 7704
rect 4709 7695 4767 7701
rect 6454 7692 6460 7704
rect 6512 7692 6518 7744
rect 10962 7732 10968 7744
rect 10923 7704 10968 7732
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 12529 7735 12587 7741
rect 12529 7701 12541 7735
rect 12575 7732 12587 7735
rect 12710 7732 12716 7744
rect 12575 7704 12716 7732
rect 12575 7701 12587 7704
rect 12529 7695 12587 7701
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 14274 7692 14280 7744
rect 14332 7732 14338 7744
rect 14642 7732 14648 7744
rect 14332 7704 14648 7732
rect 14332 7692 14338 7704
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 6089 7531 6147 7537
rect 6089 7528 6101 7531
rect 5500 7500 6101 7528
rect 5500 7488 5506 7500
rect 6089 7497 6101 7500
rect 6135 7497 6147 7531
rect 7006 7528 7012 7540
rect 6967 7500 7012 7528
rect 6089 7491 6147 7497
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 8202 7528 8208 7540
rect 7975 7500 8208 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 8297 7531 8355 7537
rect 8297 7497 8309 7531
rect 8343 7528 8355 7531
rect 8386 7528 8392 7540
rect 8343 7500 8392 7528
rect 8343 7497 8355 7500
rect 8297 7491 8355 7497
rect 1448 7327 1506 7333
rect 1448 7293 1460 7327
rect 1494 7324 1506 7327
rect 1854 7324 1860 7336
rect 1494 7296 1860 7324
rect 1494 7293 1506 7296
rect 1448 7287 1506 7293
rect 1854 7284 1860 7296
rect 1912 7284 1918 7336
rect 5074 7284 5080 7336
rect 5132 7324 5138 7336
rect 5169 7327 5227 7333
rect 5169 7324 5181 7327
rect 5132 7296 5181 7324
rect 5132 7284 5138 7296
rect 5169 7293 5181 7296
rect 5215 7293 5227 7327
rect 5169 7287 5227 7293
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6788 7296 6837 7324
rect 6788 7284 6794 7296
rect 6825 7293 6837 7296
rect 6871 7324 6883 7327
rect 7285 7327 7343 7333
rect 7285 7324 7297 7327
rect 6871 7296 7297 7324
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 7285 7293 7297 7296
rect 7331 7293 7343 7327
rect 7285 7287 7343 7293
rect 1535 7259 1593 7265
rect 1535 7225 1547 7259
rect 1581 7256 1593 7259
rect 5442 7256 5448 7268
rect 1581 7228 5448 7256
rect 1581 7225 1593 7228
rect 1535 7219 1593 7225
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 5718 7216 5724 7268
rect 5776 7256 5782 7268
rect 5813 7259 5871 7265
rect 5813 7256 5825 7259
rect 5776 7228 5825 7256
rect 5776 7216 5782 7228
rect 5813 7225 5825 7228
rect 5859 7256 5871 7259
rect 5994 7256 6000 7268
rect 5859 7228 6000 7256
rect 5859 7225 5871 7228
rect 5813 7219 5871 7225
rect 5994 7216 6000 7228
rect 6052 7256 6058 7268
rect 6457 7259 6515 7265
rect 6457 7256 6469 7259
rect 6052 7228 6469 7256
rect 6052 7216 6058 7228
rect 6457 7225 6469 7228
rect 6503 7225 6515 7259
rect 8312 7256 8340 7491
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 8846 7488 8852 7540
rect 8904 7528 8910 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 8904 7500 9597 7528
rect 8904 7488 8910 7500
rect 9585 7497 9597 7500
rect 9631 7528 9643 7531
rect 10318 7528 10324 7540
rect 9631 7500 10324 7528
rect 9631 7497 9643 7500
rect 9585 7491 9643 7497
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 11882 7528 11888 7540
rect 11843 7500 11888 7528
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12250 7528 12256 7540
rect 12211 7500 12256 7528
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 12575 7531 12633 7537
rect 12575 7528 12587 7531
rect 12492 7500 12587 7528
rect 12492 7488 12498 7500
rect 12575 7497 12587 7500
rect 12621 7497 12633 7531
rect 12575 7491 12633 7497
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 13587 7531 13645 7537
rect 13587 7528 13599 7531
rect 12768 7500 13599 7528
rect 12768 7488 12774 7500
rect 13587 7497 13599 7500
rect 13633 7497 13645 7531
rect 13587 7491 13645 7497
rect 15381 7531 15439 7537
rect 15381 7497 15393 7531
rect 15427 7528 15439 7531
rect 15838 7528 15844 7540
rect 15427 7500 15844 7528
rect 15427 7497 15439 7500
rect 15381 7491 15439 7497
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 9950 7460 9956 7472
rect 9911 7432 9956 7460
rect 9950 7420 9956 7432
rect 10008 7420 10014 7472
rect 12989 7463 13047 7469
rect 12989 7429 13001 7463
rect 13035 7460 13047 7463
rect 13170 7460 13176 7472
rect 13035 7432 13176 7460
rect 13035 7429 13047 7432
rect 12989 7423 13047 7429
rect 8754 7352 8760 7404
rect 8812 7392 8818 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 8812 7364 10517 7392
rect 8812 7352 8818 7364
rect 10505 7361 10517 7364
rect 10551 7392 10563 7395
rect 10870 7392 10876 7404
rect 10551 7364 10876 7392
rect 10551 7361 10563 7364
rect 10505 7355 10563 7361
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 8389 7327 8447 7333
rect 8389 7293 8401 7327
rect 8435 7324 8447 7327
rect 9766 7324 9772 7336
rect 8435 7296 9772 7324
rect 8435 7293 8447 7296
rect 8389 7287 8447 7293
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 12504 7327 12562 7333
rect 12504 7293 12516 7327
rect 12550 7324 12562 7327
rect 13004 7324 13032 7423
rect 13170 7420 13176 7432
rect 13228 7420 13234 7472
rect 14274 7392 14280 7404
rect 14235 7364 14280 7392
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 13484 7327 13542 7333
rect 13484 7324 13496 7327
rect 12550 7296 13032 7324
rect 13280 7296 13496 7324
rect 12550 7293 12562 7296
rect 12504 7287 12562 7293
rect 8710 7259 8768 7265
rect 8710 7256 8722 7259
rect 8312 7228 8722 7256
rect 6457 7219 6515 7225
rect 8710 7225 8722 7228
rect 8756 7225 8768 7259
rect 8710 7219 8768 7225
rect 9858 7216 9864 7268
rect 9916 7256 9922 7268
rect 10229 7259 10287 7265
rect 10229 7256 10241 7259
rect 9916 7228 10241 7256
rect 9916 7216 9922 7228
rect 10229 7225 10241 7228
rect 10275 7225 10287 7259
rect 10229 7219 10287 7225
rect 4522 7188 4528 7200
rect 4483 7160 4528 7188
rect 4522 7148 4528 7160
rect 4580 7148 4586 7200
rect 4982 7188 4988 7200
rect 4943 7160 4988 7188
rect 4982 7148 4988 7160
rect 5040 7148 5046 7200
rect 9306 7188 9312 7200
rect 9267 7160 9312 7188
rect 9306 7148 9312 7160
rect 9364 7148 9370 7200
rect 10244 7188 10272 7219
rect 10318 7216 10324 7268
rect 10376 7256 10382 7268
rect 10376 7228 10421 7256
rect 10376 7216 10382 7228
rect 12894 7216 12900 7268
rect 12952 7256 12958 7268
rect 13280 7265 13308 7296
rect 13484 7293 13496 7296
rect 13530 7324 13542 7327
rect 15746 7324 15752 7336
rect 13530 7296 15752 7324
rect 13530 7293 13542 7296
rect 13484 7287 13542 7293
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 13265 7259 13323 7265
rect 13265 7256 13277 7259
rect 12952 7228 13277 7256
rect 12952 7216 12958 7228
rect 13265 7225 13277 7228
rect 13311 7225 13323 7259
rect 13265 7219 13323 7225
rect 11149 7191 11207 7197
rect 11149 7188 11161 7191
rect 10244 7160 11161 7188
rect 11149 7157 11161 7160
rect 11195 7157 11207 7191
rect 15654 7188 15660 7200
rect 15615 7160 15660 7188
rect 11149 7151 11207 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 6089 6987 6147 6993
rect 6089 6984 6101 6987
rect 4028 6956 6101 6984
rect 4028 6944 4034 6956
rect 6089 6953 6101 6956
rect 6135 6953 6147 6987
rect 6089 6947 6147 6953
rect 9125 6987 9183 6993
rect 9125 6953 9137 6987
rect 9171 6984 9183 6987
rect 9766 6984 9772 6996
rect 9171 6956 9772 6984
rect 9171 6953 9183 6956
rect 9125 6947 9183 6953
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 10134 6984 10140 6996
rect 10095 6956 10140 6984
rect 10134 6944 10140 6956
rect 10192 6944 10198 6996
rect 13863 6987 13921 6993
rect 13863 6953 13875 6987
rect 13909 6984 13921 6987
rect 14642 6984 14648 6996
rect 13909 6956 14648 6984
rect 13909 6953 13921 6956
rect 13863 6947 13921 6953
rect 14642 6944 14648 6956
rect 14700 6944 14706 6996
rect 5442 6876 5448 6928
rect 5500 6916 5506 6928
rect 7837 6919 7895 6925
rect 7837 6916 7849 6919
rect 5500 6888 7849 6916
rect 5500 6876 5506 6888
rect 7837 6885 7849 6888
rect 7883 6916 7895 6919
rect 8110 6916 8116 6928
rect 7883 6888 8116 6916
rect 7883 6885 7895 6888
rect 7837 6879 7895 6885
rect 8110 6876 8116 6888
rect 8168 6876 8174 6928
rect 8757 6919 8815 6925
rect 8757 6885 8769 6919
rect 8803 6916 8815 6919
rect 10042 6916 10048 6928
rect 8803 6888 10048 6916
rect 8803 6885 8815 6888
rect 8757 6879 8815 6885
rect 10042 6876 10048 6888
rect 10100 6916 10106 6928
rect 10597 6919 10655 6925
rect 10597 6916 10609 6919
rect 10100 6888 10609 6916
rect 10100 6876 10106 6888
rect 10597 6885 10609 6888
rect 10643 6885 10655 6919
rect 10597 6879 10655 6885
rect 10962 6876 10968 6928
rect 11020 6916 11026 6928
rect 11330 6916 11336 6928
rect 11020 6888 11336 6916
rect 11020 6876 11026 6888
rect 11330 6876 11336 6888
rect 11388 6876 11394 6928
rect 11885 6919 11943 6925
rect 11885 6885 11897 6919
rect 11931 6916 11943 6919
rect 13262 6916 13268 6928
rect 11931 6888 13268 6916
rect 11931 6885 11943 6888
rect 11885 6879 11943 6885
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 5350 6808 5356 6860
rect 5408 6848 5414 6860
rect 5629 6851 5687 6857
rect 5629 6848 5641 6851
rect 5408 6820 5641 6848
rect 5408 6808 5414 6820
rect 5629 6817 5641 6820
rect 5675 6817 5687 6851
rect 5629 6811 5687 6817
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 5905 6851 5963 6857
rect 5776 6820 5821 6848
rect 5776 6808 5782 6820
rect 5905 6817 5917 6851
rect 5951 6817 5963 6851
rect 5905 6811 5963 6817
rect 4982 6740 4988 6792
rect 5040 6780 5046 6792
rect 5534 6780 5540 6792
rect 5040 6752 5540 6780
rect 5040 6740 5046 6752
rect 5534 6740 5540 6752
rect 5592 6780 5598 6792
rect 5920 6780 5948 6811
rect 7742 6808 7748 6860
rect 7800 6848 7806 6860
rect 12795 6857 12823 6888
rect 13262 6876 13268 6888
rect 13320 6876 13326 6928
rect 13814 6857 13820 6860
rect 8021 6851 8079 6857
rect 8021 6848 8033 6851
rect 7800 6820 8033 6848
rect 7800 6808 7806 6820
rect 8021 6817 8033 6820
rect 8067 6817 8079 6851
rect 8021 6811 8079 6817
rect 8481 6851 8539 6857
rect 8481 6817 8493 6851
rect 8527 6817 8539 6851
rect 8481 6811 8539 6817
rect 12780 6851 12838 6857
rect 12780 6817 12792 6851
rect 12826 6817 12838 6851
rect 12780 6811 12838 6817
rect 13792 6851 13820 6857
rect 13792 6817 13804 6851
rect 13872 6848 13878 6860
rect 17862 6848 17868 6860
rect 13872 6820 17868 6848
rect 13792 6811 13820 6817
rect 5592 6752 5948 6780
rect 5592 6740 5598 6752
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 8496 6780 8524 6811
rect 13814 6808 13820 6811
rect 13872 6808 13878 6820
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 7984 6752 8524 6780
rect 7984 6740 7990 6752
rect 10870 6740 10876 6792
rect 10928 6780 10934 6792
rect 11241 6783 11299 6789
rect 11241 6780 11253 6783
rect 10928 6752 11253 6780
rect 10928 6740 10934 6752
rect 11241 6749 11253 6752
rect 11287 6780 11299 6783
rect 11698 6780 11704 6792
rect 11287 6752 11704 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 1535 6715 1593 6721
rect 1535 6681 1547 6715
rect 1581 6712 1593 6715
rect 9858 6712 9864 6724
rect 1581 6684 9864 6712
rect 1581 6681 1593 6684
rect 1535 6675 1593 6681
rect 9858 6672 9864 6684
rect 9916 6672 9922 6724
rect 5074 6644 5080 6656
rect 5035 6616 5080 6644
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 12851 6647 12909 6653
rect 12851 6613 12863 6647
rect 12897 6644 12909 6647
rect 13078 6644 13084 6656
rect 12897 6616 13084 6644
rect 12897 6613 12909 6616
rect 12851 6607 12909 6613
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 106 6400 112 6452
rect 164 6440 170 6452
rect 1394 6440 1400 6452
rect 164 6412 1400 6440
rect 164 6400 170 6412
rect 1394 6400 1400 6412
rect 1452 6440 1458 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1452 6412 1593 6440
rect 1452 6400 1458 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 5994 6440 6000 6452
rect 5955 6412 6000 6440
rect 1581 6403 1639 6409
rect 5994 6400 6000 6412
rect 6052 6400 6058 6452
rect 7926 6400 7932 6452
rect 7984 6440 7990 6452
rect 8021 6443 8079 6449
rect 8021 6440 8033 6443
rect 7984 6412 8033 6440
rect 7984 6400 7990 6412
rect 8021 6409 8033 6412
rect 8067 6409 8079 6443
rect 8386 6440 8392 6452
rect 8347 6412 8392 6440
rect 8021 6403 8079 6409
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 11330 6440 11336 6452
rect 11291 6412 11336 6440
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 11698 6440 11704 6452
rect 11659 6412 11704 6440
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 12805 6443 12863 6449
rect 12805 6409 12817 6443
rect 12851 6440 12863 6443
rect 13170 6440 13176 6452
rect 12851 6412 13176 6440
rect 12851 6409 12863 6412
rect 12805 6403 12863 6409
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 13872 6412 13917 6440
rect 13872 6400 13878 6412
rect 5350 6332 5356 6384
rect 5408 6372 5414 6384
rect 6365 6375 6423 6381
rect 6365 6372 6377 6375
rect 5408 6344 6377 6372
rect 5408 6332 5414 6344
rect 6365 6341 6377 6344
rect 6411 6341 6423 6375
rect 6365 6335 6423 6341
rect 13265 6375 13323 6381
rect 13265 6341 13277 6375
rect 13311 6372 13323 6375
rect 14642 6372 14648 6384
rect 13311 6344 14648 6372
rect 13311 6341 13323 6344
rect 13265 6335 13323 6341
rect 14642 6332 14648 6344
rect 14700 6332 14706 6384
rect 7742 6304 7748 6316
rect 7703 6276 7748 6304
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 8662 6304 8668 6316
rect 8619 6276 8668 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 9508 6276 10241 6304
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 9508 6245 9536 6276
rect 10229 6273 10241 6276
rect 10275 6304 10287 6307
rect 10502 6304 10508 6316
rect 10275 6276 10508 6304
rect 10275 6273 10287 6276
rect 10229 6267 10287 6273
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 10870 6304 10876 6316
rect 10831 6276 10876 6304
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 9493 6239 9551 6245
rect 9493 6236 9505 6239
rect 8812 6208 9505 6236
rect 8812 6196 8818 6208
rect 9493 6205 9505 6208
rect 9539 6205 9551 6239
rect 13078 6236 13084 6248
rect 13039 6208 13084 6236
rect 9493 6199 9551 6205
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 8386 6128 8392 6180
rect 8444 6168 8450 6180
rect 8894 6171 8952 6177
rect 8894 6168 8906 6171
rect 8444 6140 8906 6168
rect 8444 6128 8450 6140
rect 8894 6137 8906 6140
rect 8940 6137 8952 6171
rect 8894 6131 8952 6137
rect 9861 6171 9919 6177
rect 9861 6137 9873 6171
rect 9907 6168 9919 6171
rect 10413 6171 10471 6177
rect 10413 6168 10425 6171
rect 9907 6140 10425 6168
rect 9907 6137 9919 6140
rect 9861 6131 9919 6137
rect 10413 6137 10425 6140
rect 10459 6137 10471 6171
rect 10413 6131 10471 6137
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 5629 6103 5687 6109
rect 5629 6100 5641 6103
rect 5592 6072 5641 6100
rect 5592 6060 5598 6072
rect 5629 6069 5641 6072
rect 5675 6069 5687 6103
rect 10428 6100 10456 6131
rect 10502 6128 10508 6180
rect 10560 6168 10566 6180
rect 11514 6168 11520 6180
rect 10560 6140 11520 6168
rect 10560 6128 10566 6140
rect 11514 6128 11520 6140
rect 11572 6128 11578 6180
rect 10962 6100 10968 6112
rect 10428 6072 10968 6100
rect 5629 6063 5687 6069
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8720 5868 8953 5896
rect 8720 5856 8726 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 10042 5896 10048 5908
rect 9955 5868 10048 5896
rect 8941 5859 8999 5865
rect 10042 5856 10048 5868
rect 10100 5896 10106 5908
rect 10100 5868 10916 5896
rect 10100 5856 10106 5868
rect 10888 5840 10916 5868
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 12851 5899 12909 5905
rect 12851 5896 12863 5899
rect 11020 5868 12863 5896
rect 11020 5856 11026 5868
rect 12851 5865 12863 5868
rect 12897 5865 12909 5899
rect 12851 5859 12909 5865
rect 13078 5856 13084 5908
rect 13136 5896 13142 5908
rect 13173 5899 13231 5905
rect 13173 5896 13185 5899
rect 13136 5868 13185 5896
rect 13136 5856 13142 5868
rect 13173 5865 13185 5868
rect 13219 5865 13231 5899
rect 13173 5859 13231 5865
rect 10321 5831 10379 5837
rect 10321 5797 10333 5831
rect 10367 5828 10379 5831
rect 10686 5828 10692 5840
rect 10367 5800 10692 5828
rect 10367 5797 10379 5800
rect 10321 5791 10379 5797
rect 10686 5788 10692 5800
rect 10744 5788 10750 5840
rect 10870 5828 10876 5840
rect 10831 5800 10876 5828
rect 10870 5788 10876 5800
rect 10928 5788 10934 5840
rect 8478 5760 8484 5772
rect 8439 5732 8484 5760
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 11790 5720 11796 5772
rect 11848 5760 11854 5772
rect 12710 5760 12716 5772
rect 12768 5769 12774 5772
rect 12768 5763 12806 5769
rect 11848 5732 12716 5760
rect 11848 5720 11854 5732
rect 12710 5720 12716 5732
rect 12794 5729 12806 5763
rect 12768 5723 12806 5729
rect 12768 5720 12774 5723
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 10229 5695 10287 5701
rect 10229 5692 10241 5695
rect 9548 5664 10241 5692
rect 9548 5652 9554 5664
rect 10229 5661 10241 5664
rect 10275 5692 10287 5695
rect 11701 5695 11759 5701
rect 11701 5692 11713 5695
rect 10275 5664 11713 5692
rect 10275 5661 10287 5664
rect 10229 5655 10287 5661
rect 11701 5661 11713 5664
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 7926 5584 7932 5636
rect 7984 5624 7990 5636
rect 8665 5627 8723 5633
rect 8665 5624 8677 5627
rect 7984 5596 8677 5624
rect 7984 5584 7990 5596
rect 8665 5593 8677 5596
rect 8711 5593 8723 5627
rect 8665 5587 8723 5593
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 8297 5355 8355 5361
rect 8297 5321 8309 5355
rect 8343 5352 8355 5355
rect 8478 5352 8484 5364
rect 8343 5324 8484 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 9490 5352 9496 5364
rect 9451 5324 9496 5352
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 12710 5352 12716 5364
rect 12671 5324 12716 5352
rect 12710 5312 12716 5324
rect 12768 5312 12774 5364
rect 7190 5244 7196 5296
rect 7248 5284 7254 5296
rect 8662 5284 8668 5296
rect 7248 5256 8668 5284
rect 7248 5244 7254 5256
rect 8662 5244 8668 5256
rect 8720 5244 8726 5296
rect 10042 5216 10048 5228
rect 10003 5188 10048 5216
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10321 5219 10379 5225
rect 10321 5216 10333 5219
rect 10192 5188 10333 5216
rect 10192 5176 10198 5188
rect 10321 5185 10333 5188
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 7929 5083 7987 5089
rect 7929 5049 7941 5083
rect 7975 5080 7987 5083
rect 8478 5080 8484 5092
rect 7975 5052 8484 5080
rect 7975 5049 7987 5052
rect 7929 5043 7987 5049
rect 8478 5040 8484 5052
rect 8536 5040 8542 5092
rect 8573 5083 8631 5089
rect 8573 5049 8585 5083
rect 8619 5080 8631 5083
rect 8754 5080 8760 5092
rect 8619 5052 8760 5080
rect 8619 5049 8631 5052
rect 8573 5043 8631 5049
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 9122 5080 9128 5092
rect 9083 5052 9128 5080
rect 9122 5040 9128 5052
rect 9180 5040 9186 5092
rect 10137 5083 10195 5089
rect 10137 5049 10149 5083
rect 10183 5049 10195 5083
rect 10137 5043 10195 5049
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 9732 4984 9781 5012
rect 9732 4972 9738 4984
rect 9769 4981 9781 4984
rect 9815 5012 9827 5015
rect 10152 5012 10180 5043
rect 9815 4984 10180 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 11054 5012 11060 5024
rect 10744 4984 11060 5012
rect 10744 4972 10750 4984
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 8711 4811 8769 4817
rect 8711 4808 8723 4811
rect 8536 4780 8723 4808
rect 8536 4768 8542 4780
rect 8711 4777 8723 4780
rect 8757 4777 8769 4811
rect 8711 4771 8769 4777
rect 9306 4700 9312 4752
rect 9364 4740 9370 4752
rect 9766 4740 9772 4752
rect 9364 4712 9772 4740
rect 9364 4700 9370 4712
rect 9766 4700 9772 4712
rect 9824 4740 9830 4752
rect 10045 4743 10103 4749
rect 10045 4740 10057 4743
rect 9824 4712 10057 4740
rect 9824 4700 9830 4712
rect 10045 4709 10057 4712
rect 10091 4709 10103 4743
rect 10045 4703 10103 4709
rect 11054 4700 11060 4752
rect 11112 4740 11118 4752
rect 11425 4743 11483 4749
rect 11425 4740 11437 4743
rect 11112 4712 11437 4740
rect 11112 4700 11118 4712
rect 11425 4709 11437 4712
rect 11471 4709 11483 4743
rect 11425 4703 11483 4709
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 8662 4672 8668 4684
rect 8619 4644 8668 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 8662 4632 8668 4644
rect 8720 4632 8726 4684
rect 11514 4672 11520 4684
rect 11475 4644 11520 4672
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 8481 4607 8539 4613
rect 8481 4573 8493 4607
rect 8527 4604 8539 4607
rect 8754 4604 8760 4616
rect 8527 4576 8760 4604
rect 8527 4573 8539 4576
rect 8481 4567 8539 4573
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 9950 4604 9956 4616
rect 9911 4576 9956 4604
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4573 10287 4607
rect 10229 4567 10287 4573
rect 9398 4496 9404 4548
rect 9456 4536 9462 4548
rect 10134 4536 10140 4548
rect 9456 4508 10140 4536
rect 9456 4496 9462 4508
rect 10134 4496 10140 4508
rect 10192 4536 10198 4548
rect 10244 4536 10272 4567
rect 10192 4508 10272 4536
rect 10192 4496 10198 4508
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 10870 4468 10876 4480
rect 10008 4440 10876 4468
rect 10008 4428 10014 4440
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 8662 4264 8668 4276
rect 8623 4236 8668 4264
rect 8662 4224 8668 4236
rect 8720 4224 8726 4276
rect 9122 4224 9128 4276
rect 9180 4264 9186 4276
rect 9217 4267 9275 4273
rect 9217 4264 9229 4267
rect 9180 4236 9229 4264
rect 9180 4224 9186 4236
rect 9217 4233 9229 4236
rect 9263 4264 9275 4267
rect 9950 4264 9956 4276
rect 9263 4236 9956 4264
rect 9263 4233 9275 4236
rect 9217 4227 9275 4233
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 10134 4224 10140 4276
rect 10192 4264 10198 4276
rect 10229 4267 10287 4273
rect 10229 4264 10241 4267
rect 10192 4236 10241 4264
rect 10192 4224 10198 4236
rect 10229 4233 10241 4236
rect 10275 4264 10287 4267
rect 11054 4264 11060 4276
rect 10275 4236 11060 4264
rect 10275 4233 10287 4236
rect 10229 4227 10287 4233
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 11514 4264 11520 4276
rect 11475 4236 11520 4264
rect 11514 4224 11520 4236
rect 11572 4224 11578 4276
rect 9766 4128 9772 4140
rect 9727 4100 9772 4128
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4128 10471 4131
rect 10686 4128 10692 4140
rect 10459 4100 10692 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 10686 4088 10692 4100
rect 10744 4088 10750 4140
rect 10870 4128 10876 4140
rect 10831 4100 10876 4128
rect 10870 4088 10876 4100
rect 10928 4088 10934 4140
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 9398 4060 9404 4072
rect 9355 4032 9404 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 9398 4020 9404 4032
rect 9456 4020 9462 4072
rect 20232 4063 20290 4069
rect 20232 4029 20244 4063
rect 20278 4060 20290 4063
rect 20278 4032 20760 4060
rect 20278 4029 20290 4032
rect 20232 4023 20290 4029
rect 10505 3995 10563 4001
rect 10505 3961 10517 3995
rect 10551 3961 10563 3995
rect 10505 3955 10563 3961
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 9447 3927 9505 3933
rect 9447 3924 9459 3927
rect 8812 3896 9459 3924
rect 8812 3884 8818 3896
rect 9447 3893 9459 3896
rect 9493 3893 9505 3927
rect 9447 3887 9505 3893
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10520 3924 10548 3955
rect 10192 3896 10548 3924
rect 10192 3884 10198 3896
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 20732 3933 20760 4032
rect 20303 3927 20361 3933
rect 20303 3924 20315 3927
rect 10836 3896 20315 3924
rect 10836 3884 10842 3896
rect 20303 3893 20315 3896
rect 20349 3893 20361 3927
rect 20303 3887 20361 3893
rect 20717 3927 20775 3933
rect 20717 3893 20729 3927
rect 20763 3924 20775 3927
rect 21726 3924 21732 3936
rect 20763 3896 21732 3924
rect 20763 3893 20775 3896
rect 20717 3887 20775 3893
rect 21726 3884 21732 3896
rect 21784 3884 21790 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 9398 3720 9404 3732
rect 9359 3692 9404 3720
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 10778 3720 10784 3732
rect 10739 3692 10784 3720
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 9674 3652 9680 3664
rect 9635 3624 9680 3652
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 9766 3584 9772 3596
rect 9727 3556 9772 3584
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 8754 3176 8760 3188
rect 8715 3148 8760 3176
rect 8754 3136 8760 3148
rect 8812 3136 8818 3188
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 11330 3136 11336 3188
rect 11388 3176 11394 3188
rect 11425 3179 11483 3185
rect 11425 3176 11437 3179
rect 11388 3148 11437 3176
rect 11388 3136 11394 3148
rect 11425 3145 11437 3148
rect 11471 3145 11483 3179
rect 11425 3139 11483 3145
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 8849 2975 8907 2981
rect 8849 2972 8861 2975
rect 8812 2944 8861 2972
rect 8812 2932 8818 2944
rect 8849 2941 8861 2944
rect 8895 2941 8907 2975
rect 8849 2935 8907 2941
rect 11032 2975 11090 2981
rect 11032 2941 11044 2975
rect 11078 2972 11090 2975
rect 11330 2972 11336 2984
rect 11078 2944 11336 2972
rect 11078 2941 11090 2944
rect 11032 2935 11090 2941
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 5626 2864 5632 2916
rect 5684 2904 5690 2916
rect 12618 2904 12624 2916
rect 5684 2876 12624 2904
rect 5684 2864 5690 2876
rect 12618 2864 12624 2876
rect 12676 2864 12682 2916
rect 9033 2839 9091 2845
rect 9033 2805 9045 2839
rect 9079 2836 9091 2839
rect 9306 2836 9312 2848
rect 9079 2808 9312 2836
rect 9079 2805 9091 2808
rect 9033 2799 9091 2805
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 10962 2796 10968 2848
rect 11020 2836 11026 2848
rect 11103 2839 11161 2845
rect 11103 2836 11115 2839
rect 11020 2808 11115 2836
rect 11020 2796 11026 2808
rect 11103 2805 11115 2808
rect 11149 2805 11161 2839
rect 11103 2799 11161 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 4338 2592 4344 2644
rect 4396 2632 4402 2644
rect 4479 2635 4537 2641
rect 4479 2632 4491 2635
rect 4396 2604 4491 2632
rect 4396 2592 4402 2604
rect 4479 2601 4491 2604
rect 4525 2601 4537 2635
rect 4479 2595 4537 2601
rect 5491 2635 5549 2641
rect 5491 2601 5503 2635
rect 5537 2632 5549 2635
rect 5626 2632 5632 2644
rect 5537 2604 5632 2632
rect 5537 2601 5549 2604
rect 5491 2595 5549 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 10962 2632 10968 2644
rect 10923 2604 10968 2632
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 12759 2635 12817 2641
rect 12759 2601 12771 2635
rect 12805 2632 12817 2635
rect 13446 2632 13452 2644
rect 12805 2604 13452 2632
rect 12805 2601 12817 2604
rect 12759 2595 12817 2601
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 19383 2635 19441 2641
rect 19383 2601 19395 2635
rect 19429 2632 19441 2635
rect 19518 2632 19524 2644
rect 19429 2604 19524 2632
rect 19429 2601 19441 2604
rect 19383 2595 19441 2601
rect 19518 2592 19524 2604
rect 19576 2592 19582 2644
rect 4408 2499 4466 2505
rect 4408 2465 4420 2499
rect 4454 2496 4466 2499
rect 4614 2496 4620 2508
rect 4454 2468 4620 2496
rect 4454 2465 4466 2468
rect 4408 2459 4466 2465
rect 4614 2456 4620 2468
rect 4672 2496 4678 2508
rect 4801 2499 4859 2505
rect 4801 2496 4813 2499
rect 4672 2468 4813 2496
rect 4672 2456 4678 2468
rect 4801 2465 4813 2468
rect 4847 2465 4859 2499
rect 4801 2459 4859 2465
rect 5420 2499 5478 2505
rect 5420 2465 5432 2499
rect 5466 2496 5478 2499
rect 10321 2499 10379 2505
rect 5466 2468 5948 2496
rect 5466 2465 5478 2468
rect 5420 2459 5478 2465
rect 5920 2301 5948 2468
rect 10321 2465 10333 2499
rect 10367 2496 10379 2499
rect 10980 2496 11008 2592
rect 10367 2468 11008 2496
rect 12688 2499 12746 2505
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 12688 2465 12700 2499
rect 12734 2496 12746 2499
rect 13170 2496 13176 2508
rect 12734 2468 13176 2496
rect 12734 2465 12746 2468
rect 12688 2459 12746 2465
rect 13170 2456 13176 2468
rect 13228 2456 13234 2508
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14369 2499 14427 2505
rect 14369 2496 14381 2499
rect 13872 2468 14381 2496
rect 13872 2456 13878 2468
rect 14369 2465 14381 2468
rect 14415 2465 14427 2499
rect 15746 2496 15752 2508
rect 15659 2468 15752 2496
rect 14369 2459 14427 2465
rect 15746 2456 15752 2468
rect 15804 2496 15810 2508
rect 16850 2496 16856 2508
rect 15804 2468 16436 2496
rect 16811 2468 16856 2496
rect 15804 2456 15810 2468
rect 16408 2437 16436 2468
rect 16850 2456 16856 2468
rect 16908 2496 16914 2508
rect 17405 2499 17463 2505
rect 17405 2496 17417 2499
rect 16908 2468 17417 2496
rect 16908 2456 16914 2468
rect 17405 2465 17417 2468
rect 17451 2465 17463 2499
rect 17405 2459 17463 2465
rect 19312 2499 19370 2505
rect 19312 2465 19324 2499
rect 19358 2496 19370 2499
rect 19358 2468 19840 2496
rect 19358 2465 19370 2468
rect 19312 2459 19370 2465
rect 16393 2431 16451 2437
rect 16393 2397 16405 2431
rect 16439 2428 16451 2431
rect 19426 2428 19432 2440
rect 16439 2400 19432 2428
rect 16439 2397 16451 2400
rect 16393 2391 16451 2397
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 19812 2437 19840 2468
rect 20070 2456 20076 2508
rect 20128 2496 20134 2508
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 20128 2468 22753 2496
rect 20128 2456 20134 2468
rect 22741 2465 22753 2468
rect 22787 2496 22799 2499
rect 23293 2499 23351 2505
rect 23293 2496 23305 2499
rect 22787 2468 23305 2496
rect 22787 2465 22799 2468
rect 22741 2459 22799 2465
rect 23293 2465 23305 2468
rect 23339 2465 23351 2499
rect 23293 2459 23351 2465
rect 24210 2456 24216 2508
rect 24268 2496 24274 2508
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 24268 2468 24593 2496
rect 24268 2456 24274 2468
rect 24581 2465 24593 2468
rect 24627 2496 24639 2499
rect 25133 2499 25191 2505
rect 25133 2496 25145 2499
rect 24627 2468 25145 2496
rect 24627 2465 24639 2468
rect 24581 2459 24639 2465
rect 25133 2465 25145 2468
rect 25179 2465 25191 2499
rect 25133 2459 25191 2465
rect 19797 2431 19855 2437
rect 19797 2397 19809 2431
rect 19843 2428 19855 2431
rect 26050 2428 26056 2440
rect 19843 2400 26056 2428
rect 19843 2397 19855 2400
rect 19797 2391 19855 2397
rect 26050 2388 26056 2400
rect 26108 2388 26114 2440
rect 14001 2363 14059 2369
rect 14001 2329 14013 2363
rect 14047 2360 14059 2363
rect 15470 2360 15476 2372
rect 14047 2332 15476 2360
rect 14047 2329 14059 2332
rect 14001 2323 14059 2329
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 15933 2363 15991 2369
rect 15933 2329 15945 2363
rect 15979 2360 15991 2363
rect 16758 2360 16764 2372
rect 15979 2332 16764 2360
rect 15979 2329 15991 2332
rect 15933 2323 15991 2329
rect 16758 2320 16764 2332
rect 16816 2320 16822 2372
rect 22925 2363 22983 2369
rect 22925 2329 22937 2363
rect 22971 2360 22983 2363
rect 24854 2360 24860 2372
rect 22971 2332 24860 2360
rect 22971 2329 22983 2332
rect 22925 2323 22983 2329
rect 24854 2320 24860 2332
rect 24912 2320 24918 2372
rect 5905 2295 5963 2301
rect 5905 2261 5917 2295
rect 5951 2292 5963 2295
rect 5994 2292 6000 2304
rect 5951 2264 6000 2292
rect 5951 2261 5963 2264
rect 5905 2255 5963 2261
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 10505 2295 10563 2301
rect 10505 2261 10517 2295
rect 10551 2292 10563 2295
rect 10778 2292 10784 2304
rect 10551 2264 10784 2292
rect 10551 2261 10563 2264
rect 10505 2255 10563 2261
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 13170 2292 13176 2304
rect 13131 2264 13176 2292
rect 13170 2252 13176 2264
rect 13228 2252 13234 2304
rect 17037 2295 17095 2301
rect 17037 2261 17049 2295
rect 17083 2292 17095 2295
rect 18046 2292 18052 2304
rect 17083 2264 18052 2292
rect 17083 2261 17095 2264
rect 17037 2255 17095 2261
rect 18046 2252 18052 2264
rect 18104 2252 18110 2304
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 24765 2295 24823 2301
rect 24765 2292 24777 2295
rect 18748 2264 24777 2292
rect 18748 2252 18754 2264
rect 24765 2261 24777 2264
rect 24811 2261 24823 2295
rect 24765 2255 24823 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 3050 76 3056 128
rect 3108 116 3114 128
rect 3786 116 3792 128
rect 3108 88 3792 116
rect 3108 76 3114 88
rect 3786 76 3792 88
rect 3844 76 3850 128
rect 11054 76 11060 128
rect 11112 116 11118 128
rect 11974 116 11980 128
rect 11112 88 11980 116
rect 11112 76 11118 88
rect 11974 76 11980 88
rect 12032 76 12038 128
rect 12526 76 12532 128
rect 12584 116 12590 128
rect 13262 116 13268 128
rect 12584 88 13268 116
rect 12584 76 12590 88
rect 13262 76 13268 88
rect 13320 76 13326 128
rect 22186 76 22192 128
rect 22244 116 22250 128
rect 23382 116 23388 128
rect 22244 88 23388 116
rect 22244 76 22250 88
rect 23382 76 23388 88
rect 23440 76 23446 128
rect 26234 76 26240 128
rect 26292 116 26298 128
rect 27246 116 27252 128
rect 26292 88 27252 116
rect 26292 76 26298 88
rect 27246 76 27252 88
rect 27304 76 27310 128
<< via1 >>
rect 13452 27480 13504 27532
rect 14740 27480 14792 27532
rect 15292 27480 15344 27532
rect 26424 27480 26476 27532
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 11428 25347 11480 25356
rect 11428 25313 11437 25347
rect 11437 25313 11471 25347
rect 11471 25313 11480 25347
rect 11428 25304 11480 25313
rect 13544 25304 13596 25356
rect 14556 25304 14608 25356
rect 15384 25304 15436 25356
rect 11336 25236 11388 25288
rect 12992 25168 13044 25220
rect 10784 25100 10836 25152
rect 12624 25100 12676 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10784 24939 10836 24948
rect 10784 24905 10793 24939
rect 10793 24905 10827 24939
rect 10827 24905 10836 24939
rect 10784 24896 10836 24905
rect 11060 24939 11112 24948
rect 11060 24905 11069 24939
rect 11069 24905 11103 24939
rect 11103 24905 11112 24939
rect 11060 24896 11112 24905
rect 14556 24939 14608 24948
rect 14556 24905 14565 24939
rect 14565 24905 14599 24939
rect 14599 24905 14608 24939
rect 14556 24896 14608 24905
rect 11704 24828 11756 24880
rect 14096 24828 14148 24880
rect 14464 24828 14516 24880
rect 10784 24692 10836 24744
rect 11428 24692 11480 24744
rect 12348 24692 12400 24744
rect 13084 24760 13136 24812
rect 13544 24803 13596 24812
rect 13544 24769 13553 24803
rect 13553 24769 13587 24803
rect 13587 24769 13596 24803
rect 13544 24760 13596 24769
rect 15292 24896 15344 24948
rect 11244 24624 11296 24676
rect 9220 24556 9272 24608
rect 9312 24599 9364 24608
rect 9312 24565 9321 24599
rect 9321 24565 9355 24599
rect 9355 24565 9364 24599
rect 9312 24556 9364 24565
rect 12072 24556 12124 24608
rect 12716 24599 12768 24608
rect 12716 24565 12725 24599
rect 12725 24565 12759 24599
rect 12759 24565 12768 24599
rect 12716 24556 12768 24565
rect 14280 24556 14332 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 5448 24352 5500 24404
rect 6460 24352 6512 24404
rect 9220 24352 9272 24404
rect 9680 24352 9732 24404
rect 12440 24352 12492 24404
rect 23388 24352 23440 24404
rect 12624 24327 12676 24336
rect 12624 24293 12633 24327
rect 12633 24293 12667 24327
rect 12667 24293 12676 24327
rect 12624 24284 12676 24293
rect 12808 24284 12860 24336
rect 1216 24216 1268 24268
rect 5356 24216 5408 24268
rect 8944 24216 8996 24268
rect 10324 24216 10376 24268
rect 14096 24259 14148 24268
rect 14096 24225 14105 24259
rect 14105 24225 14139 24259
rect 14139 24225 14148 24259
rect 14096 24216 14148 24225
rect 10876 24148 10928 24200
rect 12900 24191 12952 24200
rect 12900 24157 12909 24191
rect 12909 24157 12943 24191
rect 12943 24157 12952 24191
rect 12900 24148 12952 24157
rect 12532 24080 12584 24132
rect 8392 24012 8444 24064
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1216 23808 1268 23860
rect 8944 23851 8996 23860
rect 8944 23817 8953 23851
rect 8953 23817 8987 23851
rect 8987 23817 8996 23851
rect 8944 23808 8996 23817
rect 10140 23808 10192 23860
rect 10324 23851 10376 23860
rect 10324 23817 10333 23851
rect 10333 23817 10367 23851
rect 10367 23817 10376 23851
rect 10324 23808 10376 23817
rect 11980 23808 12032 23860
rect 9036 23740 9088 23792
rect 12900 23740 12952 23792
rect 10876 23715 10928 23724
rect 10876 23681 10885 23715
rect 10885 23681 10919 23715
rect 10919 23681 10928 23715
rect 10876 23672 10928 23681
rect 12532 23715 12584 23724
rect 12532 23681 12541 23715
rect 12541 23681 12575 23715
rect 12575 23681 12584 23715
rect 12532 23672 12584 23681
rect 14004 23740 14056 23792
rect 16396 23808 16448 23860
rect 17408 23808 17460 23860
rect 20444 23808 20496 23860
rect 24216 23808 24268 23860
rect 22376 23740 22428 23792
rect 14280 23672 14332 23724
rect 14372 23715 14424 23724
rect 14372 23681 14381 23715
rect 14381 23681 14415 23715
rect 14415 23681 14424 23715
rect 14372 23672 14424 23681
rect 14556 23672 14608 23724
rect 1124 23604 1176 23656
rect 2688 23604 2740 23656
rect 3700 23604 3752 23656
rect 4436 23604 4488 23656
rect 7012 23647 7064 23656
rect 7012 23613 7021 23647
rect 7021 23613 7055 23647
rect 7055 23613 7064 23647
rect 7012 23604 7064 23613
rect 9404 23647 9456 23656
rect 9404 23613 9413 23647
rect 9413 23613 9447 23647
rect 9447 23613 9456 23647
rect 9404 23604 9456 23613
rect 9680 23647 9732 23656
rect 9680 23613 9689 23647
rect 9689 23613 9723 23647
rect 9723 23613 9732 23647
rect 9680 23604 9732 23613
rect 18604 23672 18656 23724
rect 17316 23604 17368 23656
rect 18512 23647 18564 23656
rect 18512 23613 18521 23647
rect 18521 23613 18555 23647
rect 18555 23613 18564 23647
rect 18512 23604 18564 23613
rect 1676 23468 1728 23520
rect 3424 23468 3476 23520
rect 3700 23468 3752 23520
rect 7104 23468 7156 23520
rect 7932 23468 7984 23520
rect 12532 23536 12584 23588
rect 13176 23579 13228 23588
rect 11428 23468 11480 23520
rect 12164 23468 12216 23520
rect 13176 23545 13185 23579
rect 13185 23545 13219 23579
rect 13219 23545 13228 23579
rect 13176 23536 13228 23545
rect 14188 23579 14240 23588
rect 14188 23545 14197 23579
rect 14197 23545 14231 23579
rect 14231 23545 14240 23579
rect 14188 23536 14240 23545
rect 19984 23536 20036 23588
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 7012 23264 7064 23316
rect 7104 23264 7156 23316
rect 11244 23264 11296 23316
rect 14096 23307 14148 23316
rect 14096 23273 14105 23307
rect 14105 23273 14139 23307
rect 14139 23273 14148 23307
rect 14096 23264 14148 23273
rect 14372 23307 14424 23316
rect 14372 23273 14381 23307
rect 14381 23273 14415 23307
rect 14415 23273 14424 23307
rect 14372 23264 14424 23273
rect 18604 23264 18656 23316
rect 6368 23239 6420 23248
rect 6368 23205 6377 23239
rect 6377 23205 6411 23239
rect 6411 23205 6420 23239
rect 6368 23196 6420 23205
rect 11336 23239 11388 23248
rect 11336 23205 11345 23239
rect 11345 23205 11379 23239
rect 11379 23205 11388 23239
rect 11336 23196 11388 23205
rect 11428 23239 11480 23248
rect 11428 23205 11437 23239
rect 11437 23205 11471 23239
rect 11471 23205 11480 23239
rect 12900 23239 12952 23248
rect 11428 23196 11480 23205
rect 12900 23205 12909 23239
rect 12909 23205 12943 23239
rect 12943 23205 12952 23239
rect 12900 23196 12952 23205
rect 13268 23196 13320 23248
rect 4988 23128 5040 23180
rect 8484 23128 8536 23180
rect 9772 23171 9824 23180
rect 9772 23137 9781 23171
rect 9781 23137 9815 23171
rect 9815 23137 9824 23171
rect 9772 23128 9824 23137
rect 9956 23128 10008 23180
rect 16120 23128 16172 23180
rect 6276 23103 6328 23112
rect 6276 23069 6285 23103
rect 6285 23069 6319 23103
rect 6319 23069 6328 23103
rect 6276 23060 6328 23069
rect 7196 23060 7248 23112
rect 11796 23060 11848 23112
rect 13176 23103 13228 23112
rect 13176 23069 13185 23103
rect 13185 23069 13219 23103
rect 13219 23069 13228 23103
rect 13176 23060 13228 23069
rect 10324 22924 10376 22976
rect 10784 22967 10836 22976
rect 10784 22933 10793 22967
rect 10793 22933 10827 22967
rect 10827 22933 10836 22967
rect 10784 22924 10836 22933
rect 12808 22924 12860 22976
rect 13268 22924 13320 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 3424 22720 3476 22772
rect 6276 22720 6328 22772
rect 6368 22720 6420 22772
rect 8484 22763 8536 22772
rect 8484 22729 8493 22763
rect 8493 22729 8527 22763
rect 8527 22729 8536 22763
rect 8484 22720 8536 22729
rect 11336 22763 11388 22772
rect 11336 22729 11345 22763
rect 11345 22729 11379 22763
rect 11379 22729 11388 22763
rect 11336 22720 11388 22729
rect 11428 22720 11480 22772
rect 12624 22763 12676 22772
rect 12624 22729 12633 22763
rect 12633 22729 12667 22763
rect 12667 22729 12676 22763
rect 12624 22720 12676 22729
rect 13268 22720 13320 22772
rect 16120 22763 16172 22772
rect 9772 22695 9824 22704
rect 9772 22661 9781 22695
rect 9781 22661 9815 22695
rect 9815 22661 9824 22695
rect 9772 22652 9824 22661
rect 11152 22652 11204 22704
rect 14096 22652 14148 22704
rect 16120 22729 16129 22763
rect 16129 22729 16163 22763
rect 16163 22729 16172 22763
rect 16120 22720 16172 22729
rect 19432 22720 19484 22772
rect 7104 22584 7156 22636
rect 7196 22627 7248 22636
rect 7196 22593 7205 22627
rect 7205 22593 7239 22627
rect 7239 22593 7248 22627
rect 10324 22627 10376 22636
rect 7196 22584 7248 22593
rect 10324 22593 10333 22627
rect 10333 22593 10367 22627
rect 10367 22593 10376 22627
rect 10324 22584 10376 22593
rect 14372 22584 14424 22636
rect 8668 22559 8720 22568
rect 8668 22525 8677 22559
rect 8677 22525 8711 22559
rect 8711 22525 8720 22559
rect 8668 22516 8720 22525
rect 7012 22491 7064 22500
rect 7012 22457 7021 22491
rect 7021 22457 7055 22491
rect 7055 22457 7064 22491
rect 7012 22448 7064 22457
rect 9404 22491 9456 22500
rect 9404 22457 9413 22491
rect 9413 22457 9447 22491
rect 9447 22457 9456 22491
rect 9404 22448 9456 22457
rect 11980 22516 12032 22568
rect 10784 22448 10836 22500
rect 10968 22491 11020 22500
rect 10968 22457 10977 22491
rect 10977 22457 11011 22491
rect 11011 22457 11020 22491
rect 10968 22448 11020 22457
rect 13728 22491 13780 22500
rect 13728 22457 13737 22491
rect 13737 22457 13771 22491
rect 13771 22457 13780 22491
rect 13728 22448 13780 22457
rect 4988 22380 5040 22432
rect 6000 22380 6052 22432
rect 9956 22380 10008 22432
rect 14004 22380 14056 22432
rect 15476 22516 15528 22568
rect 14924 22423 14976 22432
rect 14924 22389 14933 22423
rect 14933 22389 14967 22423
rect 14967 22389 14976 22423
rect 14924 22380 14976 22389
rect 15384 22423 15436 22432
rect 15384 22389 15393 22423
rect 15393 22389 15427 22423
rect 15427 22389 15436 22423
rect 15384 22380 15436 22389
rect 19156 22423 19208 22432
rect 19156 22389 19165 22423
rect 19165 22389 19199 22423
rect 19199 22389 19208 22423
rect 19156 22380 19208 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 7012 22176 7064 22228
rect 6368 22108 6420 22160
rect 6920 22108 6972 22160
rect 9772 22108 9824 22160
rect 11428 22176 11480 22228
rect 11888 22219 11940 22228
rect 11888 22185 11897 22219
rect 11897 22185 11931 22219
rect 11931 22185 11940 22219
rect 11888 22176 11940 22185
rect 12900 22219 12952 22228
rect 12900 22185 12909 22219
rect 12909 22185 12943 22219
rect 12943 22185 12952 22219
rect 12900 22176 12952 22185
rect 13728 22176 13780 22228
rect 19156 22176 19208 22228
rect 10968 22151 11020 22160
rect 10968 22117 10977 22151
rect 10977 22117 11011 22151
rect 11011 22117 11020 22151
rect 10968 22108 11020 22117
rect 11520 22108 11572 22160
rect 20 22040 72 22092
rect 2044 22083 2096 22092
rect 2044 22049 2088 22083
rect 2088 22049 2096 22083
rect 2044 22040 2096 22049
rect 5356 22040 5408 22092
rect 6184 22040 6236 22092
rect 11612 22040 11664 22092
rect 12072 22040 12124 22092
rect 12256 22083 12308 22092
rect 12256 22049 12265 22083
rect 12265 22049 12299 22083
rect 12299 22049 12308 22083
rect 12256 22040 12308 22049
rect 13176 22108 13228 22160
rect 13636 22108 13688 22160
rect 14096 22151 14148 22160
rect 14096 22117 14105 22151
rect 14105 22117 14139 22151
rect 14139 22117 14148 22151
rect 14096 22108 14148 22117
rect 17408 22108 17460 22160
rect 13268 22083 13320 22092
rect 13268 22049 13277 22083
rect 13277 22049 13311 22083
rect 13311 22049 13320 22083
rect 13268 22040 13320 22049
rect 15844 22083 15896 22092
rect 6000 21972 6052 22024
rect 7288 21972 7340 22024
rect 8944 21972 8996 22024
rect 10692 21972 10744 22024
rect 5540 21904 5592 21956
rect 8668 21947 8720 21956
rect 8668 21913 8677 21947
rect 8677 21913 8711 21947
rect 8711 21913 8720 21947
rect 8668 21904 8720 21913
rect 12256 21904 12308 21956
rect 14924 21972 14976 22024
rect 15844 22049 15853 22083
rect 15853 22049 15887 22083
rect 15887 22049 15896 22083
rect 15844 22040 15896 22049
rect 18328 22083 18380 22092
rect 18328 22049 18337 22083
rect 18337 22049 18371 22083
rect 18371 22049 18380 22083
rect 18328 22040 18380 22049
rect 16028 22015 16080 22024
rect 16028 21981 16037 22015
rect 16037 21981 16071 22015
rect 16071 21981 16080 22015
rect 16028 21972 16080 21981
rect 17684 22015 17736 22024
rect 17684 21981 17693 22015
rect 17693 21981 17727 22015
rect 17727 21981 17736 22015
rect 17684 21972 17736 21981
rect 15660 21904 15712 21956
rect 2596 21836 2648 21888
rect 4344 21879 4396 21888
rect 4344 21845 4353 21879
rect 4353 21845 4387 21879
rect 4387 21845 4396 21879
rect 4344 21836 4396 21845
rect 6092 21836 6144 21888
rect 6736 21836 6788 21888
rect 16488 21879 16540 21888
rect 16488 21845 16497 21879
rect 16497 21845 16531 21879
rect 16531 21845 16540 21879
rect 16488 21836 16540 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2044 21675 2096 21684
rect 2044 21641 2053 21675
rect 2053 21641 2087 21675
rect 2087 21641 2096 21675
rect 2044 21632 2096 21641
rect 6000 21632 6052 21684
rect 7012 21632 7064 21684
rect 8024 21632 8076 21684
rect 9772 21675 9824 21684
rect 9772 21641 9781 21675
rect 9781 21641 9815 21675
rect 9815 21641 9824 21675
rect 9772 21632 9824 21641
rect 10784 21632 10836 21684
rect 13176 21632 13228 21684
rect 13636 21632 13688 21684
rect 15476 21632 15528 21684
rect 20168 21675 20220 21684
rect 5356 21607 5408 21616
rect 2688 21496 2740 21548
rect 5356 21573 5365 21607
rect 5365 21573 5399 21607
rect 5399 21573 5408 21607
rect 5356 21564 5408 21573
rect 9680 21564 9732 21616
rect 11612 21564 11664 21616
rect 14280 21564 14332 21616
rect 4344 21539 4396 21548
rect 4344 21505 4353 21539
rect 4353 21505 4387 21539
rect 4387 21505 4396 21539
rect 4344 21496 4396 21505
rect 6092 21496 6144 21548
rect 8852 21496 8904 21548
rect 8944 21539 8996 21548
rect 8944 21505 8953 21539
rect 8953 21505 8987 21539
rect 8987 21505 8996 21539
rect 8944 21496 8996 21505
rect 9956 21496 10008 21548
rect 12256 21496 12308 21548
rect 13268 21539 13320 21548
rect 13268 21505 13277 21539
rect 13277 21505 13311 21539
rect 13311 21505 13320 21539
rect 13268 21496 13320 21505
rect 14096 21496 14148 21548
rect 4988 21403 5040 21412
rect 3976 21292 4028 21344
rect 4988 21369 4997 21403
rect 4997 21369 5031 21403
rect 5031 21369 5040 21403
rect 4988 21360 5040 21369
rect 6644 21403 6696 21412
rect 6644 21369 6653 21403
rect 6653 21369 6687 21403
rect 6687 21369 6696 21403
rect 6644 21360 6696 21369
rect 7748 21360 7800 21412
rect 10048 21428 10100 21480
rect 14924 21471 14976 21480
rect 14924 21437 14933 21471
rect 14933 21437 14967 21471
rect 14967 21437 14976 21471
rect 14924 21428 14976 21437
rect 20168 21641 20177 21675
rect 20177 21641 20211 21675
rect 20211 21641 20220 21675
rect 20168 21632 20220 21641
rect 8484 21360 8536 21412
rect 5080 21292 5132 21344
rect 6184 21292 6236 21344
rect 8024 21292 8076 21344
rect 13360 21403 13412 21412
rect 13360 21369 13369 21403
rect 13369 21369 13403 21403
rect 13403 21369 13412 21403
rect 16488 21428 16540 21480
rect 20168 21428 20220 21480
rect 25412 21632 25464 21684
rect 15568 21403 15620 21412
rect 13360 21360 13412 21369
rect 10140 21335 10192 21344
rect 10140 21301 10149 21335
rect 10149 21301 10183 21335
rect 10183 21301 10192 21335
rect 10140 21292 10192 21301
rect 11612 21292 11664 21344
rect 14280 21292 14332 21344
rect 15568 21369 15577 21403
rect 15577 21369 15611 21403
rect 15611 21369 15620 21403
rect 15568 21360 15620 21369
rect 15844 21360 15896 21412
rect 17592 21360 17644 21412
rect 18144 21403 18196 21412
rect 18144 21369 18153 21403
rect 18153 21369 18187 21403
rect 18187 21369 18196 21403
rect 18144 21360 18196 21369
rect 16488 21335 16540 21344
rect 16488 21301 16497 21335
rect 16497 21301 16531 21335
rect 16531 21301 16540 21335
rect 16488 21292 16540 21301
rect 16948 21292 17000 21344
rect 17408 21335 17460 21344
rect 17408 21301 17417 21335
rect 17417 21301 17451 21335
rect 17451 21301 17460 21335
rect 17408 21292 17460 21301
rect 17776 21335 17828 21344
rect 17776 21301 17785 21335
rect 17785 21301 17819 21335
rect 17819 21301 17828 21335
rect 18328 21360 18380 21412
rect 20076 21360 20128 21412
rect 17776 21292 17828 21301
rect 19524 21292 19576 21344
rect 20536 21292 20588 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1584 21131 1636 21140
rect 1584 21097 1593 21131
rect 1593 21097 1627 21131
rect 1627 21097 1636 21131
rect 1584 21088 1636 21097
rect 6920 21131 6972 21140
rect 6920 21097 6929 21131
rect 6929 21097 6963 21131
rect 6963 21097 6972 21131
rect 6920 21088 6972 21097
rect 8852 21131 8904 21140
rect 8852 21097 8861 21131
rect 8861 21097 8895 21131
rect 8895 21097 8904 21131
rect 8852 21088 8904 21097
rect 10692 21131 10744 21140
rect 10692 21097 10701 21131
rect 10701 21097 10735 21131
rect 10735 21097 10744 21131
rect 10692 21088 10744 21097
rect 11336 21131 11388 21140
rect 11336 21097 11345 21131
rect 11345 21097 11379 21131
rect 11379 21097 11388 21131
rect 11336 21088 11388 21097
rect 12164 21088 12216 21140
rect 13728 21088 13780 21140
rect 14924 21131 14976 21140
rect 14924 21097 14933 21131
rect 14933 21097 14967 21131
rect 14967 21097 14976 21131
rect 14924 21088 14976 21097
rect 15660 21088 15712 21140
rect 16028 21131 16080 21140
rect 16028 21097 16037 21131
rect 16037 21097 16071 21131
rect 16071 21097 16080 21131
rect 16028 21088 16080 21097
rect 4252 21063 4304 21072
rect 4252 21029 4261 21063
rect 4261 21029 4295 21063
rect 4295 21029 4304 21063
rect 4252 21020 4304 21029
rect 6092 21020 6144 21072
rect 6644 21020 6696 21072
rect 7932 21063 7984 21072
rect 7932 21029 7941 21063
rect 7941 21029 7975 21063
rect 7975 21029 7984 21063
rect 7932 21020 7984 21029
rect 8024 21063 8076 21072
rect 8024 21029 8033 21063
rect 8033 21029 8067 21063
rect 8067 21029 8076 21063
rect 8024 21020 8076 21029
rect 13176 21020 13228 21072
rect 1768 20952 1820 21004
rect 9680 20952 9732 21004
rect 11888 20952 11940 21004
rect 12900 20952 12952 21004
rect 15384 20952 15436 21004
rect 16396 21088 16448 21140
rect 17776 21088 17828 21140
rect 19524 21088 19576 21140
rect 17684 21063 17736 21072
rect 17684 21029 17693 21063
rect 17693 21029 17727 21063
rect 17727 21029 17736 21063
rect 17684 21020 17736 21029
rect 18972 21020 19024 21072
rect 3792 20884 3844 20936
rect 4436 20927 4488 20936
rect 4436 20893 4445 20927
rect 4445 20893 4479 20927
rect 4479 20893 4488 20927
rect 4436 20884 4488 20893
rect 6000 20927 6052 20936
rect 6000 20893 6009 20927
rect 6009 20893 6043 20927
rect 6043 20893 6052 20927
rect 6000 20884 6052 20893
rect 7656 20884 7708 20936
rect 11796 20884 11848 20936
rect 14096 20884 14148 20936
rect 18144 20884 18196 20936
rect 6184 20816 6236 20868
rect 11612 20816 11664 20868
rect 19248 20884 19300 20936
rect 20536 20884 20588 20936
rect 20352 20816 20404 20868
rect 4804 20748 4856 20800
rect 10048 20748 10100 20800
rect 18144 20791 18196 20800
rect 18144 20757 18153 20791
rect 18153 20757 18187 20791
rect 18187 20757 18196 20791
rect 18144 20748 18196 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2596 20587 2648 20596
rect 2596 20553 2605 20587
rect 2605 20553 2639 20587
rect 2639 20553 2648 20587
rect 4252 20587 4304 20596
rect 2596 20544 2648 20553
rect 4252 20553 4261 20587
rect 4261 20553 4295 20587
rect 4295 20553 4304 20587
rect 4252 20544 4304 20553
rect 6092 20587 6144 20596
rect 6092 20553 6101 20587
rect 6101 20553 6135 20587
rect 6135 20553 6144 20587
rect 6092 20544 6144 20553
rect 6920 20544 6972 20596
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 11428 20544 11480 20596
rect 11888 20587 11940 20596
rect 11888 20553 11897 20587
rect 11897 20553 11931 20587
rect 11931 20553 11940 20587
rect 11888 20544 11940 20553
rect 13636 20544 13688 20596
rect 14096 20587 14148 20596
rect 14096 20553 14105 20587
rect 14105 20553 14139 20587
rect 14139 20553 14148 20587
rect 14096 20544 14148 20553
rect 4344 20476 4396 20528
rect 4436 20408 4488 20460
rect 4804 20451 4856 20460
rect 4804 20417 4813 20451
rect 4813 20417 4847 20451
rect 4847 20417 4856 20451
rect 4804 20408 4856 20417
rect 17868 20476 17920 20528
rect 20812 20476 20864 20528
rect 25136 20519 25188 20528
rect 25136 20485 25145 20519
rect 25145 20485 25179 20519
rect 25179 20485 25188 20519
rect 25136 20476 25188 20485
rect 6736 20408 6788 20460
rect 7656 20451 7708 20460
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 9404 20408 9456 20460
rect 10692 20408 10744 20460
rect 12900 20451 12952 20460
rect 12900 20417 12909 20451
rect 12909 20417 12943 20451
rect 12943 20417 12952 20451
rect 12900 20408 12952 20417
rect 15568 20408 15620 20460
rect 17684 20408 17736 20460
rect 18880 20408 18932 20460
rect 19524 20408 19576 20460
rect 8852 20340 8904 20392
rect 15108 20383 15160 20392
rect 1768 20204 1820 20256
rect 2964 20247 3016 20256
rect 2964 20213 2973 20247
rect 2973 20213 3007 20247
rect 3007 20213 3016 20247
rect 2964 20204 3016 20213
rect 3148 20204 3200 20256
rect 4252 20204 4304 20256
rect 7012 20272 7064 20324
rect 15108 20349 15117 20383
rect 15117 20349 15151 20383
rect 15151 20349 15160 20383
rect 15108 20340 15160 20349
rect 6368 20204 6420 20256
rect 8484 20204 8536 20256
rect 9680 20204 9732 20256
rect 10140 20272 10192 20324
rect 11336 20272 11388 20324
rect 13176 20272 13228 20324
rect 15384 20272 15436 20324
rect 16396 20272 16448 20324
rect 18144 20315 18196 20324
rect 18144 20281 18153 20315
rect 18153 20281 18187 20315
rect 18187 20281 18196 20315
rect 18144 20272 18196 20281
rect 15476 20204 15528 20256
rect 17776 20247 17828 20256
rect 17776 20213 17785 20247
rect 17785 20213 17819 20247
rect 17819 20213 17828 20247
rect 18328 20272 18380 20324
rect 19340 20272 19392 20324
rect 20352 20315 20404 20324
rect 20352 20281 20361 20315
rect 20361 20281 20395 20315
rect 20395 20281 20404 20315
rect 20352 20272 20404 20281
rect 17776 20204 17828 20213
rect 18972 20204 19024 20256
rect 19524 20204 19576 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 3792 20043 3844 20052
rect 3792 20009 3801 20043
rect 3801 20009 3835 20043
rect 3835 20009 3844 20043
rect 3792 20000 3844 20009
rect 6000 20000 6052 20052
rect 8024 20000 8076 20052
rect 10692 20043 10744 20052
rect 10692 20009 10701 20043
rect 10701 20009 10735 20043
rect 10735 20009 10744 20043
rect 10692 20000 10744 20009
rect 13360 20000 13412 20052
rect 14188 20000 14240 20052
rect 14832 20000 14884 20052
rect 16396 20043 16448 20052
rect 16396 20009 16405 20043
rect 16405 20009 16439 20043
rect 16439 20009 16448 20043
rect 16396 20000 16448 20009
rect 16948 20043 17000 20052
rect 16948 20009 16957 20043
rect 16957 20009 16991 20043
rect 16991 20009 17000 20043
rect 16948 20000 17000 20009
rect 18144 20000 18196 20052
rect 3148 19975 3200 19984
rect 3148 19941 3157 19975
rect 3157 19941 3191 19975
rect 3191 19941 3200 19975
rect 3148 19932 3200 19941
rect 4068 19932 4120 19984
rect 4988 19932 5040 19984
rect 6736 19932 6788 19984
rect 2964 19907 3016 19916
rect 2964 19873 2973 19907
rect 2973 19873 3007 19907
rect 3007 19873 3016 19907
rect 2964 19864 3016 19873
rect 6184 19864 6236 19916
rect 6368 19907 6420 19916
rect 6368 19873 6377 19907
rect 6377 19873 6411 19907
rect 6411 19873 6420 19907
rect 6368 19864 6420 19873
rect 7748 19864 7800 19916
rect 9680 19932 9732 19984
rect 11060 19932 11112 19984
rect 12164 19932 12216 19984
rect 13176 19932 13228 19984
rect 13912 19932 13964 19984
rect 18328 19975 18380 19984
rect 18328 19941 18337 19975
rect 18337 19941 18371 19975
rect 18371 19941 18380 19975
rect 18328 19932 18380 19941
rect 18880 19975 18932 19984
rect 18880 19941 18889 19975
rect 18889 19941 18923 19975
rect 18923 19941 18932 19975
rect 18880 19932 18932 19941
rect 19248 19975 19300 19984
rect 19248 19941 19257 19975
rect 19257 19941 19291 19975
rect 19291 19941 19300 19975
rect 19248 19932 19300 19941
rect 9404 19864 9456 19916
rect 12716 19907 12768 19916
rect 12716 19873 12725 19907
rect 12725 19873 12759 19907
rect 12759 19873 12768 19907
rect 12716 19864 12768 19873
rect 16120 19864 16172 19916
rect 16488 19864 16540 19916
rect 19708 19907 19760 19916
rect 19708 19873 19717 19907
rect 19717 19873 19751 19907
rect 19751 19873 19760 19907
rect 19708 19864 19760 19873
rect 3884 19796 3936 19848
rect 4436 19796 4488 19848
rect 7380 19796 7432 19848
rect 11336 19796 11388 19848
rect 11520 19839 11572 19848
rect 11520 19805 11529 19839
rect 11529 19805 11563 19839
rect 11563 19805 11572 19839
rect 11520 19796 11572 19805
rect 17868 19796 17920 19848
rect 20 19660 72 19712
rect 4988 19660 5040 19712
rect 8760 19703 8812 19712
rect 8760 19669 8769 19703
rect 8769 19669 8803 19703
rect 8803 19669 8812 19703
rect 8760 19660 8812 19669
rect 9956 19660 10008 19712
rect 19432 19660 19484 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 6184 19499 6236 19508
rect 6184 19465 6193 19499
rect 6193 19465 6227 19499
rect 6227 19465 6236 19499
rect 6184 19456 6236 19465
rect 11060 19499 11112 19508
rect 4344 19320 4396 19372
rect 7472 19388 7524 19440
rect 8208 19388 8260 19440
rect 11060 19465 11069 19499
rect 11069 19465 11103 19499
rect 11103 19465 11112 19499
rect 11060 19456 11112 19465
rect 11336 19499 11388 19508
rect 11336 19465 11345 19499
rect 11345 19465 11379 19499
rect 11379 19465 11388 19499
rect 11336 19456 11388 19465
rect 14096 19456 14148 19508
rect 17592 19456 17644 19508
rect 17868 19499 17920 19508
rect 17868 19465 17877 19499
rect 17877 19465 17911 19499
rect 17911 19465 17920 19499
rect 17868 19456 17920 19465
rect 19340 19499 19392 19508
rect 19340 19465 19349 19499
rect 19349 19465 19383 19499
rect 19383 19465 19392 19499
rect 19340 19456 19392 19465
rect 19432 19456 19484 19508
rect 11152 19388 11204 19440
rect 7380 19320 7432 19372
rect 7656 19320 7708 19372
rect 8668 19320 8720 19372
rect 8852 19320 8904 19372
rect 6368 19252 6420 19304
rect 13912 19320 13964 19372
rect 15384 19363 15436 19372
rect 15384 19329 15393 19363
rect 15393 19329 15427 19363
rect 15427 19329 15436 19363
rect 15384 19320 15436 19329
rect 18788 19363 18840 19372
rect 18788 19329 18797 19363
rect 18797 19329 18831 19363
rect 18831 19329 18840 19363
rect 18788 19320 18840 19329
rect 3240 19184 3292 19236
rect 2964 19116 3016 19168
rect 4344 19116 4396 19168
rect 4528 19159 4580 19168
rect 4528 19125 4537 19159
rect 4537 19125 4571 19159
rect 4571 19125 4580 19159
rect 4528 19116 4580 19125
rect 6920 19227 6972 19236
rect 6920 19193 6929 19227
rect 6929 19193 6963 19227
rect 6963 19193 6972 19227
rect 6920 19184 6972 19193
rect 7012 19227 7064 19236
rect 7012 19193 7021 19227
rect 7021 19193 7055 19227
rect 7055 19193 7064 19227
rect 7012 19184 7064 19193
rect 6736 19116 6788 19168
rect 7748 19116 7800 19168
rect 8760 19184 8812 19236
rect 9588 19184 9640 19236
rect 9956 19184 10008 19236
rect 11060 19252 11112 19304
rect 14188 19295 14240 19304
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 9404 19116 9456 19168
rect 10048 19159 10100 19168
rect 10048 19125 10057 19159
rect 10057 19125 10091 19159
rect 10091 19125 10100 19159
rect 10048 19116 10100 19125
rect 12808 19159 12860 19168
rect 12808 19125 12817 19159
rect 12817 19125 12851 19159
rect 12851 19125 12860 19159
rect 12808 19116 12860 19125
rect 13820 19184 13872 19236
rect 14372 19116 14424 19168
rect 14648 19227 14700 19236
rect 14648 19193 14657 19227
rect 14657 19193 14691 19227
rect 14691 19193 14700 19227
rect 14648 19184 14700 19193
rect 20076 19320 20128 19372
rect 15568 19295 15620 19304
rect 15568 19261 15577 19295
rect 15577 19261 15611 19295
rect 15611 19261 15620 19295
rect 15568 19252 15620 19261
rect 16304 19184 16356 19236
rect 18328 19227 18380 19236
rect 16580 19116 16632 19168
rect 18328 19193 18337 19227
rect 18337 19193 18371 19227
rect 18371 19193 18380 19227
rect 18328 19184 18380 19193
rect 19708 19295 19760 19304
rect 19708 19261 19717 19295
rect 19717 19261 19751 19295
rect 19751 19261 19760 19295
rect 19708 19252 19760 19261
rect 20076 19184 20128 19236
rect 19524 19116 19576 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 3884 18955 3936 18964
rect 3884 18921 3893 18955
rect 3893 18921 3927 18955
rect 3927 18921 3936 18955
rect 3884 18912 3936 18921
rect 7380 18912 7432 18964
rect 8668 18912 8720 18964
rect 12716 18955 12768 18964
rect 12716 18921 12725 18955
rect 12725 18921 12759 18955
rect 12759 18921 12768 18955
rect 12716 18912 12768 18921
rect 12808 18912 12860 18964
rect 13912 18912 13964 18964
rect 14648 18912 14700 18964
rect 16120 18955 16172 18964
rect 16120 18921 16129 18955
rect 16129 18921 16163 18955
rect 16163 18921 16172 18955
rect 16120 18912 16172 18921
rect 16580 18955 16632 18964
rect 16580 18921 16589 18955
rect 16589 18921 16623 18955
rect 16623 18921 16632 18955
rect 16580 18912 16632 18921
rect 18236 18912 18288 18964
rect 18328 18912 18380 18964
rect 20076 18955 20128 18964
rect 20076 18921 20085 18955
rect 20085 18921 20119 18955
rect 20119 18921 20128 18955
rect 20076 18912 20128 18921
rect 3240 18887 3292 18896
rect 3240 18853 3249 18887
rect 3249 18853 3283 18887
rect 3283 18853 3292 18887
rect 3240 18844 3292 18853
rect 4068 18887 4120 18896
rect 4068 18853 4077 18887
rect 4077 18853 4111 18887
rect 4111 18853 4120 18887
rect 4068 18844 4120 18853
rect 4528 18844 4580 18896
rect 7012 18844 7064 18896
rect 7564 18887 7616 18896
rect 7564 18853 7573 18887
rect 7573 18853 7607 18887
rect 7607 18853 7616 18887
rect 7564 18844 7616 18853
rect 10140 18844 10192 18896
rect 11796 18844 11848 18896
rect 13084 18844 13136 18896
rect 15568 18887 15620 18896
rect 15568 18853 15577 18887
rect 15577 18853 15611 18887
rect 15611 18853 15620 18887
rect 15568 18844 15620 18853
rect 17868 18844 17920 18896
rect 1308 18776 1360 18828
rect 3056 18776 3108 18828
rect 3976 18776 4028 18828
rect 4804 18776 4856 18828
rect 7288 18776 7340 18828
rect 13820 18819 13872 18828
rect 13820 18785 13829 18819
rect 13829 18785 13863 18819
rect 13863 18785 13872 18819
rect 14096 18819 14148 18828
rect 13820 18776 13872 18785
rect 14096 18785 14105 18819
rect 14105 18785 14139 18819
rect 14139 18785 14148 18819
rect 14096 18776 14148 18785
rect 19248 18776 19300 18828
rect 4436 18640 4488 18692
rect 6644 18708 6696 18760
rect 7196 18640 7248 18692
rect 9588 18640 9640 18692
rect 1676 18572 1728 18624
rect 3516 18615 3568 18624
rect 3516 18581 3525 18615
rect 3525 18581 3559 18615
rect 3559 18581 3568 18615
rect 3516 18572 3568 18581
rect 5264 18615 5316 18624
rect 5264 18581 5273 18615
rect 5273 18581 5307 18615
rect 5307 18581 5316 18615
rect 5264 18572 5316 18581
rect 7472 18572 7524 18624
rect 11244 18572 11296 18624
rect 12808 18708 12860 18760
rect 16212 18751 16264 18760
rect 16212 18717 16221 18751
rect 16221 18717 16255 18751
rect 16255 18717 16264 18751
rect 16212 18708 16264 18717
rect 18052 18751 18104 18760
rect 18052 18717 18061 18751
rect 18061 18717 18095 18751
rect 18095 18717 18104 18751
rect 18052 18708 18104 18717
rect 18420 18751 18472 18760
rect 18420 18717 18429 18751
rect 18429 18717 18463 18751
rect 18463 18717 18472 18751
rect 18420 18708 18472 18717
rect 19432 18708 19484 18760
rect 14464 18640 14516 18692
rect 18512 18640 18564 18692
rect 19340 18640 19392 18692
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 4344 18411 4396 18420
rect 4344 18377 4353 18411
rect 4353 18377 4387 18411
rect 4387 18377 4396 18411
rect 4344 18368 4396 18377
rect 6644 18411 6696 18420
rect 6644 18377 6653 18411
rect 6653 18377 6687 18411
rect 6687 18377 6696 18411
rect 6644 18368 6696 18377
rect 7564 18368 7616 18420
rect 14740 18368 14792 18420
rect 17868 18411 17920 18420
rect 5264 18300 5316 18352
rect 6460 18300 6512 18352
rect 9220 18300 9272 18352
rect 11888 18300 11940 18352
rect 13544 18300 13596 18352
rect 13728 18300 13780 18352
rect 14464 18300 14516 18352
rect 15384 18300 15436 18352
rect 17868 18377 17877 18411
rect 17877 18377 17911 18411
rect 17911 18377 17920 18411
rect 17868 18368 17920 18377
rect 19248 18300 19300 18352
rect 1308 18232 1360 18284
rect 7288 18232 7340 18284
rect 9312 18275 9364 18284
rect 9312 18241 9321 18275
rect 9321 18241 9355 18275
rect 9355 18241 9364 18275
rect 9312 18232 9364 18241
rect 9588 18275 9640 18284
rect 9588 18241 9597 18275
rect 9597 18241 9631 18275
rect 9631 18241 9640 18275
rect 9588 18232 9640 18241
rect 12624 18232 12676 18284
rect 12808 18275 12860 18284
rect 12808 18241 12817 18275
rect 12817 18241 12851 18275
rect 12851 18241 12860 18275
rect 12808 18232 12860 18241
rect 14648 18232 14700 18284
rect 18420 18275 18472 18284
rect 18420 18241 18429 18275
rect 18429 18241 18463 18275
rect 18463 18241 18472 18275
rect 18420 18232 18472 18241
rect 20352 18275 20404 18284
rect 20352 18241 20361 18275
rect 20361 18241 20395 18275
rect 20395 18241 20404 18275
rect 20352 18232 20404 18241
rect 1860 18028 1912 18080
rect 2504 18164 2556 18216
rect 3516 18164 3568 18216
rect 3884 18164 3936 18216
rect 2136 18028 2188 18080
rect 3056 18071 3108 18080
rect 3056 18037 3065 18071
rect 3065 18037 3099 18071
rect 3099 18037 3108 18071
rect 3056 18028 3108 18037
rect 3424 18028 3476 18080
rect 4804 18028 4856 18080
rect 5080 18071 5132 18080
rect 5080 18037 5089 18071
rect 5089 18037 5123 18071
rect 5123 18037 5132 18071
rect 5540 18164 5592 18216
rect 7472 18207 7524 18216
rect 5264 18096 5316 18148
rect 7472 18173 7481 18207
rect 7481 18173 7515 18207
rect 7515 18173 7524 18207
rect 7472 18164 7524 18173
rect 11428 18207 11480 18216
rect 6736 18096 6788 18148
rect 7380 18096 7432 18148
rect 5080 18028 5132 18037
rect 5540 18028 5592 18080
rect 7748 18028 7800 18080
rect 11428 18173 11437 18207
rect 11437 18173 11471 18207
rect 11471 18173 11480 18207
rect 11428 18164 11480 18173
rect 13820 18164 13872 18216
rect 16212 18164 16264 18216
rect 11520 18139 11572 18148
rect 11520 18105 11529 18139
rect 11529 18105 11563 18139
rect 11563 18105 11572 18139
rect 11520 18096 11572 18105
rect 10140 18028 10192 18080
rect 11796 18071 11848 18080
rect 11796 18037 11805 18071
rect 11805 18037 11839 18071
rect 11839 18037 11848 18071
rect 11796 18028 11848 18037
rect 12256 18071 12308 18080
rect 12256 18037 12265 18071
rect 12265 18037 12299 18071
rect 12299 18037 12308 18071
rect 15200 18096 15252 18148
rect 17132 18096 17184 18148
rect 18236 18139 18288 18148
rect 18236 18105 18245 18139
rect 18245 18105 18279 18139
rect 18279 18105 18288 18139
rect 18236 18096 18288 18105
rect 19340 18096 19392 18148
rect 14096 18071 14148 18080
rect 12256 18028 12308 18037
rect 14096 18037 14105 18071
rect 14105 18037 14139 18071
rect 14139 18037 14148 18071
rect 14096 18028 14148 18037
rect 15384 18028 15436 18080
rect 15660 18071 15712 18080
rect 15660 18037 15669 18071
rect 15669 18037 15703 18071
rect 15703 18037 15712 18071
rect 15660 18028 15712 18037
rect 19524 18028 19576 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1676 17867 1728 17876
rect 1676 17833 1685 17867
rect 1685 17833 1719 17867
rect 1719 17833 1728 17867
rect 1676 17824 1728 17833
rect 5264 17867 5316 17876
rect 5264 17833 5273 17867
rect 5273 17833 5307 17867
rect 5307 17833 5316 17867
rect 5264 17824 5316 17833
rect 6460 17867 6512 17876
rect 6460 17833 6469 17867
rect 6469 17833 6503 17867
rect 6503 17833 6512 17867
rect 6460 17824 6512 17833
rect 6920 17867 6972 17876
rect 6920 17833 6929 17867
rect 6929 17833 6963 17867
rect 6963 17833 6972 17867
rect 6920 17824 6972 17833
rect 7748 17867 7800 17876
rect 7748 17833 7757 17867
rect 7757 17833 7791 17867
rect 7791 17833 7800 17867
rect 7748 17824 7800 17833
rect 10140 17824 10192 17876
rect 1768 17756 1820 17808
rect 2412 17688 2464 17740
rect 3332 17688 3384 17740
rect 6000 17756 6052 17808
rect 9312 17799 9364 17808
rect 9312 17765 9321 17799
rect 9321 17765 9355 17799
rect 9355 17765 9364 17799
rect 9312 17756 9364 17765
rect 13912 17824 13964 17876
rect 15476 17824 15528 17876
rect 5172 17688 5224 17740
rect 9496 17688 9548 17740
rect 11520 17756 11572 17808
rect 12808 17756 12860 17808
rect 13452 17756 13504 17808
rect 13544 17756 13596 17808
rect 13820 17756 13872 17808
rect 14556 17799 14608 17808
rect 14556 17765 14565 17799
rect 14565 17765 14599 17799
rect 14599 17765 14608 17799
rect 14556 17756 14608 17765
rect 17500 17824 17552 17876
rect 18052 17824 18104 17876
rect 19524 17824 19576 17876
rect 16304 17756 16356 17808
rect 18420 17756 18472 17808
rect 10140 17731 10192 17740
rect 10140 17697 10149 17731
rect 10149 17697 10183 17731
rect 10183 17697 10192 17731
rect 10140 17688 10192 17697
rect 17592 17731 17644 17740
rect 17592 17697 17601 17731
rect 17601 17697 17635 17731
rect 17635 17697 17644 17731
rect 17592 17688 17644 17697
rect 17776 17688 17828 17740
rect 19156 17731 19208 17740
rect 19156 17697 19165 17731
rect 19165 17697 19199 17731
rect 19199 17697 19208 17731
rect 19156 17688 19208 17697
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 6644 17620 6696 17672
rect 11336 17620 11388 17672
rect 11888 17663 11940 17672
rect 11888 17629 11897 17663
rect 11897 17629 11931 17663
rect 11931 17629 11940 17663
rect 11888 17620 11940 17629
rect 2504 17595 2556 17604
rect 2504 17561 2513 17595
rect 2513 17561 2547 17595
rect 2547 17561 2556 17595
rect 2504 17552 2556 17561
rect 3516 17552 3568 17604
rect 11612 17552 11664 17604
rect 12532 17595 12584 17604
rect 12532 17561 12541 17595
rect 12541 17561 12575 17595
rect 12575 17561 12584 17595
rect 15200 17620 15252 17672
rect 12532 17552 12584 17561
rect 2872 17484 2924 17536
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 3424 17527 3476 17536
rect 3424 17493 3433 17527
rect 3433 17493 3467 17527
rect 3467 17493 3476 17527
rect 3424 17484 3476 17493
rect 4068 17484 4120 17536
rect 6736 17484 6788 17536
rect 7932 17484 7984 17536
rect 9036 17484 9088 17536
rect 10692 17527 10744 17536
rect 10692 17493 10701 17527
rect 10701 17493 10735 17527
rect 10735 17493 10744 17527
rect 10692 17484 10744 17493
rect 12624 17484 12676 17536
rect 13360 17484 13412 17536
rect 17132 17484 17184 17536
rect 18604 17527 18656 17536
rect 18604 17493 18613 17527
rect 18613 17493 18647 17527
rect 18647 17493 18656 17527
rect 18604 17484 18656 17493
rect 18972 17527 19024 17536
rect 18972 17493 18981 17527
rect 18981 17493 19015 17527
rect 19015 17493 19024 17527
rect 18972 17484 19024 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 3056 17280 3108 17332
rect 3332 17323 3384 17332
rect 3332 17289 3341 17323
rect 3341 17289 3375 17323
rect 3375 17289 3384 17323
rect 3332 17280 3384 17289
rect 4620 17280 4672 17332
rect 4804 17323 4856 17332
rect 4804 17289 4813 17323
rect 4813 17289 4847 17323
rect 4847 17289 4856 17323
rect 4804 17280 4856 17289
rect 5540 17280 5592 17332
rect 6644 17323 6696 17332
rect 6644 17289 6653 17323
rect 6653 17289 6687 17323
rect 6687 17289 6696 17323
rect 6644 17280 6696 17289
rect 6920 17280 6972 17332
rect 7380 17280 7432 17332
rect 10140 17280 10192 17332
rect 11520 17323 11572 17332
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 12808 17280 12860 17332
rect 15660 17323 15712 17332
rect 15660 17289 15669 17323
rect 15669 17289 15703 17323
rect 15703 17289 15712 17323
rect 15660 17280 15712 17289
rect 16304 17280 16356 17332
rect 19984 17280 20036 17332
rect 6000 17212 6052 17264
rect 11428 17212 11480 17264
rect 13452 17255 13504 17264
rect 13452 17221 13461 17255
rect 13461 17221 13495 17255
rect 13495 17221 13504 17255
rect 13452 17212 13504 17221
rect 27620 17212 27672 17264
rect 4068 17076 4120 17128
rect 6552 17144 6604 17196
rect 6276 17076 6328 17128
rect 6920 17076 6972 17128
rect 9404 17144 9456 17196
rect 10692 17144 10744 17196
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 12808 17187 12860 17196
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 16212 17144 16264 17196
rect 18972 17144 19024 17196
rect 7932 17076 7984 17128
rect 8116 17076 8168 17128
rect 8944 17119 8996 17128
rect 8944 17085 8953 17119
rect 8953 17085 8987 17119
rect 8987 17085 8996 17119
rect 8944 17076 8996 17085
rect 9220 17119 9272 17128
rect 9220 17085 9229 17119
rect 9229 17085 9263 17119
rect 9263 17085 9272 17119
rect 9220 17076 9272 17085
rect 10140 17076 10192 17128
rect 14556 17119 14608 17128
rect 3424 17008 3476 17060
rect 5172 17051 5224 17060
rect 5172 17017 5181 17051
rect 5181 17017 5215 17051
rect 5215 17017 5224 17051
rect 14556 17085 14565 17119
rect 14565 17085 14599 17119
rect 14599 17085 14608 17119
rect 14556 17076 14608 17085
rect 5172 17008 5224 17017
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 2412 16983 2464 16992
rect 2412 16949 2421 16983
rect 2421 16949 2455 16983
rect 2455 16949 2464 16983
rect 2412 16940 2464 16949
rect 3608 16940 3660 16992
rect 7748 16983 7800 16992
rect 7748 16949 7757 16983
rect 7757 16949 7791 16983
rect 7791 16949 7800 16983
rect 10140 16983 10192 16992
rect 7748 16940 7800 16949
rect 10140 16949 10149 16983
rect 10149 16949 10183 16983
rect 10183 16949 10192 16983
rect 10140 16940 10192 16949
rect 12256 17051 12308 17060
rect 12256 17017 12265 17051
rect 12265 17017 12299 17051
rect 12299 17017 12308 17051
rect 12624 17051 12676 17060
rect 12256 17008 12308 17017
rect 12624 17017 12633 17051
rect 12633 17017 12667 17051
rect 12667 17017 12676 17051
rect 12624 17008 12676 17017
rect 16028 17076 16080 17128
rect 18880 17119 18932 17128
rect 18880 17085 18889 17119
rect 18889 17085 18923 17119
rect 18923 17085 18932 17119
rect 18880 17076 18932 17085
rect 24216 17076 24268 17128
rect 12532 16940 12584 16992
rect 14556 16940 14608 16992
rect 15476 16940 15528 16992
rect 16764 17008 16816 17060
rect 18604 17008 18656 17060
rect 17040 16983 17092 16992
rect 17040 16949 17049 16983
rect 17049 16949 17083 16983
rect 17083 16949 17092 16983
rect 17040 16940 17092 16949
rect 17592 16983 17644 16992
rect 17592 16949 17601 16983
rect 17601 16949 17635 16983
rect 17635 16949 17644 16983
rect 17592 16940 17644 16949
rect 17684 16940 17736 16992
rect 19156 16983 19208 16992
rect 19156 16949 19165 16983
rect 19165 16949 19199 16983
rect 19199 16949 19208 16983
rect 19156 16940 19208 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 3148 16736 3200 16788
rect 2872 16668 2924 16720
rect 4068 16736 4120 16788
rect 8024 16736 8076 16788
rect 9220 16736 9272 16788
rect 9496 16779 9548 16788
rect 9496 16745 9505 16779
rect 9505 16745 9539 16779
rect 9539 16745 9548 16779
rect 9496 16736 9548 16745
rect 10140 16779 10192 16788
rect 10140 16745 10149 16779
rect 10149 16745 10183 16779
rect 10183 16745 10192 16779
rect 10140 16736 10192 16745
rect 11336 16779 11388 16788
rect 9036 16711 9088 16720
rect 1952 16643 2004 16652
rect 1952 16609 1961 16643
rect 1961 16609 1995 16643
rect 1995 16609 2004 16643
rect 1952 16600 2004 16609
rect 2780 16600 2832 16652
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4068 16600 4120 16609
rect 4712 16643 4764 16652
rect 4712 16609 4721 16643
rect 4721 16609 4755 16643
rect 4755 16609 4764 16643
rect 4712 16600 4764 16609
rect 4896 16643 4948 16652
rect 4896 16609 4905 16643
rect 4905 16609 4939 16643
rect 4939 16609 4948 16643
rect 4896 16600 4948 16609
rect 9036 16677 9045 16711
rect 9045 16677 9079 16711
rect 9079 16677 9088 16711
rect 9036 16668 9088 16677
rect 11336 16745 11345 16779
rect 11345 16745 11379 16779
rect 11379 16745 11388 16779
rect 11336 16736 11388 16745
rect 11796 16668 11848 16720
rect 12808 16736 12860 16788
rect 16764 16779 16816 16788
rect 16764 16745 16773 16779
rect 16773 16745 16807 16779
rect 16807 16745 16816 16779
rect 16764 16736 16816 16745
rect 18604 16736 18656 16788
rect 19524 16736 19576 16788
rect 12624 16668 12676 16720
rect 16948 16668 17000 16720
rect 18696 16668 18748 16720
rect 18880 16711 18932 16720
rect 18880 16677 18889 16711
rect 18889 16677 18923 16711
rect 18923 16677 18932 16711
rect 18880 16668 18932 16677
rect 7380 16643 7432 16652
rect 2228 16532 2280 16584
rect 2412 16532 2464 16584
rect 5356 16532 5408 16584
rect 1768 16464 1820 16516
rect 7380 16609 7389 16643
rect 7389 16609 7423 16643
rect 7423 16609 7432 16643
rect 7380 16600 7432 16609
rect 8576 16643 8628 16652
rect 8576 16609 8585 16643
rect 8585 16609 8619 16643
rect 8619 16609 8628 16643
rect 8576 16600 8628 16609
rect 13452 16643 13504 16652
rect 13452 16609 13461 16643
rect 13461 16609 13495 16643
rect 13495 16609 13504 16643
rect 13452 16600 13504 16609
rect 15292 16600 15344 16652
rect 17500 16600 17552 16652
rect 24676 16600 24728 16652
rect 7472 16575 7524 16584
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 9496 16532 9548 16584
rect 11612 16575 11664 16584
rect 11612 16541 11621 16575
rect 11621 16541 11655 16575
rect 11655 16541 11664 16575
rect 11612 16532 11664 16541
rect 18420 16532 18472 16584
rect 1952 16396 2004 16448
rect 3332 16396 3384 16448
rect 7748 16464 7800 16516
rect 9956 16464 10008 16516
rect 17224 16464 17276 16516
rect 8024 16439 8076 16448
rect 8024 16405 8033 16439
rect 8033 16405 8067 16439
rect 8067 16405 8076 16439
rect 8024 16396 8076 16405
rect 14832 16396 14884 16448
rect 15844 16439 15896 16448
rect 15844 16405 15853 16439
rect 15853 16405 15887 16439
rect 15887 16405 15896 16439
rect 15844 16396 15896 16405
rect 16028 16396 16080 16448
rect 17776 16396 17828 16448
rect 18052 16439 18104 16448
rect 18052 16405 18061 16439
rect 18061 16405 18095 16439
rect 18095 16405 18104 16439
rect 18052 16396 18104 16405
rect 21364 16439 21416 16448
rect 21364 16405 21373 16439
rect 21373 16405 21407 16439
rect 21407 16405 21416 16439
rect 21364 16396 21416 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2780 16192 2832 16244
rect 6552 16192 6604 16244
rect 11244 16192 11296 16244
rect 11796 16235 11848 16244
rect 11796 16201 11805 16235
rect 11805 16201 11839 16235
rect 11839 16201 11848 16235
rect 13452 16235 13504 16244
rect 11796 16192 11848 16201
rect 13452 16201 13461 16235
rect 13461 16201 13495 16235
rect 13495 16201 13504 16235
rect 13452 16192 13504 16201
rect 15292 16235 15344 16244
rect 15292 16201 15301 16235
rect 15301 16201 15335 16235
rect 15335 16201 15344 16235
rect 15292 16192 15344 16201
rect 16948 16192 17000 16244
rect 17040 16192 17092 16244
rect 18328 16192 18380 16244
rect 18696 16192 18748 16244
rect 24676 16235 24728 16244
rect 24676 16201 24685 16235
rect 24685 16201 24719 16235
rect 24719 16201 24728 16235
rect 24676 16192 24728 16201
rect 4068 16124 4120 16176
rect 7380 16124 7432 16176
rect 10140 16124 10192 16176
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 4068 16031 4120 16040
rect 4068 15997 4077 16031
rect 4077 15997 4111 16031
rect 4111 15997 4120 16031
rect 4068 15988 4120 15997
rect 4712 16031 4764 16040
rect 4712 15997 4721 16031
rect 4721 15997 4755 16031
rect 4755 15997 4764 16031
rect 4712 15988 4764 15997
rect 4896 16031 4948 16040
rect 4896 15997 4905 16031
rect 4905 15997 4939 16031
rect 4939 15997 4948 16031
rect 4896 15988 4948 15997
rect 9496 16099 9548 16108
rect 9496 16065 9505 16099
rect 9505 16065 9539 16099
rect 9539 16065 9548 16099
rect 9496 16056 9548 16065
rect 6000 15988 6052 16040
rect 7288 15988 7340 16040
rect 7932 15988 7984 16040
rect 8944 16031 8996 16040
rect 1952 15920 2004 15972
rect 2412 15920 2464 15972
rect 3792 15963 3844 15972
rect 3792 15929 3801 15963
rect 3801 15929 3835 15963
rect 3835 15929 3844 15963
rect 3792 15920 3844 15929
rect 7748 15920 7800 15972
rect 8944 15997 8953 16031
rect 8953 15997 8987 16031
rect 8987 15997 8996 16031
rect 8944 15988 8996 15997
rect 9128 15988 9180 16040
rect 9864 15988 9916 16040
rect 17500 16167 17552 16176
rect 17500 16133 17509 16167
rect 17509 16133 17543 16167
rect 17543 16133 17552 16167
rect 17500 16124 17552 16133
rect 11060 16099 11112 16108
rect 11060 16065 11069 16099
rect 11069 16065 11103 16099
rect 11103 16065 11112 16099
rect 11060 16056 11112 16065
rect 18052 16056 18104 16108
rect 18236 16099 18288 16108
rect 18236 16065 18245 16099
rect 18245 16065 18279 16099
rect 18279 16065 18288 16099
rect 18236 16056 18288 16065
rect 18880 16099 18932 16108
rect 18880 16065 18889 16099
rect 18889 16065 18923 16099
rect 18923 16065 18932 16099
rect 18880 16056 18932 16065
rect 18972 16056 19024 16108
rect 19984 16056 20036 16108
rect 21364 16099 21416 16108
rect 21364 16065 21373 16099
rect 21373 16065 21407 16099
rect 21407 16065 21416 16099
rect 21364 16056 21416 16065
rect 10784 15988 10836 16040
rect 14556 16031 14608 16040
rect 12440 15963 12492 15972
rect 12440 15929 12449 15963
rect 12449 15929 12483 15963
rect 12483 15929 12492 15963
rect 12440 15920 12492 15929
rect 3884 15852 3936 15904
rect 7564 15852 7616 15904
rect 8024 15852 8076 15904
rect 10140 15895 10192 15904
rect 10140 15861 10149 15895
rect 10149 15861 10183 15895
rect 10183 15861 10192 15895
rect 10140 15852 10192 15861
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 14832 16031 14884 16040
rect 14832 15997 14841 16031
rect 14841 15997 14875 16031
rect 14875 15997 14884 16031
rect 14832 15988 14884 15997
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 15016 15963 15068 15972
rect 15016 15929 15025 15963
rect 15025 15929 15059 15963
rect 15059 15929 15068 15963
rect 15016 15920 15068 15929
rect 12900 15852 12952 15904
rect 15476 15852 15528 15904
rect 16212 15920 16264 15972
rect 18328 15963 18380 15972
rect 18328 15929 18337 15963
rect 18337 15929 18371 15963
rect 18371 15929 18380 15963
rect 18328 15920 18380 15929
rect 19616 15920 19668 15972
rect 18880 15852 18932 15904
rect 20076 15920 20128 15972
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 3148 15648 3200 15700
rect 3516 15648 3568 15700
rect 8576 15648 8628 15700
rect 11612 15691 11664 15700
rect 11612 15657 11621 15691
rect 11621 15657 11655 15691
rect 11655 15657 11664 15691
rect 11612 15648 11664 15657
rect 15016 15648 15068 15700
rect 16212 15691 16264 15700
rect 1768 15623 1820 15632
rect 1768 15589 1777 15623
rect 1777 15589 1811 15623
rect 1811 15589 1820 15623
rect 1768 15580 1820 15589
rect 1952 15580 2004 15632
rect 3976 15580 4028 15632
rect 4160 15580 4212 15632
rect 4344 15580 4396 15632
rect 4804 15512 4856 15564
rect 7932 15580 7984 15632
rect 6276 15555 6328 15564
rect 2412 15444 2464 15496
rect 4344 15444 4396 15496
rect 2320 15419 2372 15428
rect 2320 15385 2329 15419
rect 2329 15385 2363 15419
rect 2363 15385 2372 15419
rect 2320 15376 2372 15385
rect 3148 15419 3200 15428
rect 3148 15385 3157 15419
rect 3157 15385 3191 15419
rect 3191 15385 3200 15419
rect 3148 15376 3200 15385
rect 4252 15376 4304 15428
rect 1952 15308 2004 15360
rect 3884 15308 3936 15360
rect 4620 15444 4672 15496
rect 6276 15521 6285 15555
rect 6285 15521 6319 15555
rect 6319 15521 6328 15555
rect 6276 15512 6328 15521
rect 7656 15555 7708 15564
rect 6644 15444 6696 15496
rect 7656 15521 7665 15555
rect 7665 15521 7699 15555
rect 7699 15521 7708 15555
rect 7656 15512 7708 15521
rect 7932 15444 7984 15496
rect 6276 15376 6328 15428
rect 8944 15376 8996 15428
rect 9864 15580 9916 15632
rect 11980 15580 12032 15632
rect 12440 15580 12492 15632
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 10784 15512 10836 15564
rect 13544 15555 13596 15564
rect 13544 15521 13553 15555
rect 13553 15521 13587 15555
rect 13587 15521 13596 15555
rect 13544 15512 13596 15521
rect 16212 15657 16221 15691
rect 16221 15657 16255 15691
rect 16255 15657 16264 15691
rect 16212 15648 16264 15657
rect 17408 15580 17460 15632
rect 18880 15580 18932 15632
rect 19432 15555 19484 15564
rect 19432 15521 19441 15555
rect 19441 15521 19475 15555
rect 19475 15521 19484 15555
rect 19432 15512 19484 15521
rect 11796 15444 11848 15496
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 12624 15444 12676 15496
rect 17960 15487 18012 15496
rect 17960 15453 17969 15487
rect 17969 15453 18003 15487
rect 18003 15453 18012 15487
rect 17960 15444 18012 15453
rect 9772 15419 9824 15428
rect 9772 15385 9781 15419
rect 9781 15385 9815 15419
rect 9815 15385 9824 15419
rect 9772 15376 9824 15385
rect 18420 15376 18472 15428
rect 6000 15308 6052 15360
rect 9128 15308 9180 15360
rect 10784 15351 10836 15360
rect 10784 15317 10793 15351
rect 10793 15317 10827 15351
rect 10827 15317 10836 15351
rect 10784 15308 10836 15317
rect 11060 15351 11112 15360
rect 11060 15317 11069 15351
rect 11069 15317 11103 15351
rect 11103 15317 11112 15351
rect 11060 15308 11112 15317
rect 12900 15351 12952 15360
rect 12900 15317 12909 15351
rect 12909 15317 12943 15351
rect 12943 15317 12952 15351
rect 12900 15308 12952 15317
rect 13268 15351 13320 15360
rect 13268 15317 13277 15351
rect 13277 15317 13311 15351
rect 13311 15317 13320 15351
rect 13268 15308 13320 15317
rect 17408 15308 17460 15360
rect 17868 15308 17920 15360
rect 18144 15308 18196 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2044 15104 2096 15156
rect 3148 14968 3200 15020
rect 3608 14900 3660 14952
rect 4160 14900 4212 14952
rect 4804 14968 4856 15020
rect 4620 14900 4672 14952
rect 5540 14900 5592 14952
rect 6000 14900 6052 14952
rect 10048 15104 10100 15156
rect 11980 15147 12032 15156
rect 11980 15113 11989 15147
rect 11989 15113 12023 15147
rect 12023 15113 12032 15147
rect 11980 15104 12032 15113
rect 17408 15147 17460 15156
rect 17408 15113 17417 15147
rect 17417 15113 17451 15147
rect 17451 15113 17460 15147
rect 17408 15104 17460 15113
rect 17960 15104 18012 15156
rect 12348 15036 12400 15088
rect 17776 15036 17828 15088
rect 9404 14968 9456 15020
rect 11060 14968 11112 15020
rect 13268 14968 13320 15020
rect 18144 15011 18196 15020
rect 18144 14977 18153 15011
rect 18153 14977 18187 15011
rect 18187 14977 18196 15011
rect 18144 14968 18196 14977
rect 18420 15011 18472 15020
rect 18420 14977 18429 15011
rect 18429 14977 18463 15011
rect 18463 14977 18472 15011
rect 18420 14968 18472 14977
rect 7656 14900 7708 14952
rect 7932 14943 7984 14952
rect 7932 14909 7941 14943
rect 7941 14909 7975 14943
rect 7975 14909 7984 14943
rect 7932 14900 7984 14909
rect 8300 14900 8352 14952
rect 8760 14943 8812 14952
rect 3424 14832 3476 14884
rect 5356 14832 5408 14884
rect 1400 14807 1452 14816
rect 1400 14773 1409 14807
rect 1409 14773 1443 14807
rect 1443 14773 1452 14807
rect 1400 14764 1452 14773
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 2596 14807 2648 14816
rect 2596 14773 2605 14807
rect 2605 14773 2639 14807
rect 2639 14773 2648 14807
rect 2596 14764 2648 14773
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 4068 14807 4120 14816
rect 4068 14773 4077 14807
rect 4077 14773 4111 14807
rect 4111 14773 4120 14807
rect 4068 14764 4120 14773
rect 4528 14807 4580 14816
rect 4528 14773 4537 14807
rect 4537 14773 4571 14807
rect 4571 14773 4580 14807
rect 4528 14764 4580 14773
rect 6276 14807 6328 14816
rect 6276 14773 6285 14807
rect 6285 14773 6319 14807
rect 6319 14773 6328 14807
rect 6276 14764 6328 14773
rect 7012 14807 7064 14816
rect 7012 14773 7021 14807
rect 7021 14773 7055 14807
rect 7055 14773 7064 14807
rect 7012 14764 7064 14773
rect 8760 14909 8769 14943
rect 8769 14909 8803 14943
rect 8803 14909 8812 14943
rect 8760 14900 8812 14909
rect 9128 14943 9180 14952
rect 9128 14909 9137 14943
rect 9137 14909 9171 14943
rect 9171 14909 9180 14943
rect 9128 14900 9180 14909
rect 10692 14832 10744 14884
rect 9772 14764 9824 14816
rect 10876 14807 10928 14816
rect 10876 14773 10885 14807
rect 10885 14773 10919 14807
rect 10919 14773 10928 14807
rect 10876 14764 10928 14773
rect 12900 14832 12952 14884
rect 14832 14900 14884 14952
rect 16488 14900 16540 14952
rect 13544 14807 13596 14816
rect 13544 14773 13553 14807
rect 13553 14773 13587 14807
rect 13587 14773 13596 14807
rect 13544 14764 13596 14773
rect 14280 14807 14332 14816
rect 14280 14773 14289 14807
rect 14289 14773 14323 14807
rect 14323 14773 14332 14807
rect 14280 14764 14332 14773
rect 15476 14807 15528 14816
rect 15476 14773 15485 14807
rect 15485 14773 15519 14807
rect 15519 14773 15528 14807
rect 15476 14764 15528 14773
rect 18144 14832 18196 14884
rect 18328 14832 18380 14884
rect 19800 14968 19852 15020
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 21180 14943 21232 14952
rect 21180 14909 21189 14943
rect 21189 14909 21223 14943
rect 21223 14909 21232 14943
rect 21180 14900 21232 14909
rect 19524 14832 19576 14884
rect 19800 14875 19852 14884
rect 19800 14841 19809 14875
rect 19809 14841 19843 14875
rect 19843 14841 19852 14875
rect 19800 14832 19852 14841
rect 19432 14807 19484 14816
rect 19432 14773 19441 14807
rect 19441 14773 19475 14807
rect 19475 14773 19484 14807
rect 19432 14764 19484 14773
rect 20260 14764 20312 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1952 14560 2004 14612
rect 3608 14560 3660 14612
rect 4252 14560 4304 14612
rect 6184 14603 6236 14612
rect 6184 14569 6193 14603
rect 6193 14569 6227 14603
rect 6227 14569 6236 14603
rect 6184 14560 6236 14569
rect 9680 14560 9732 14612
rect 2596 14492 2648 14544
rect 4528 14492 4580 14544
rect 11796 14560 11848 14612
rect 14832 14560 14884 14612
rect 16488 14603 16540 14612
rect 16488 14569 16497 14603
rect 16497 14569 16531 14603
rect 16531 14569 16540 14603
rect 16488 14560 16540 14569
rect 18144 14560 18196 14612
rect 18420 14560 18472 14612
rect 20076 14560 20128 14612
rect 10876 14492 10928 14544
rect 12256 14492 12308 14544
rect 12624 14535 12676 14544
rect 12624 14501 12633 14535
rect 12633 14501 12667 14535
rect 12667 14501 12676 14535
rect 12624 14492 12676 14501
rect 13268 14492 13320 14544
rect 15476 14492 15528 14544
rect 17224 14535 17276 14544
rect 17224 14501 17233 14535
rect 17233 14501 17267 14535
rect 17267 14501 17276 14535
rect 17224 14492 17276 14501
rect 17408 14492 17460 14544
rect 17868 14535 17920 14544
rect 17868 14501 17877 14535
rect 17877 14501 17911 14535
rect 17911 14501 17920 14535
rect 17868 14492 17920 14501
rect 18052 14492 18104 14544
rect 18880 14535 18932 14544
rect 18880 14501 18889 14535
rect 18889 14501 18923 14535
rect 18923 14501 18932 14535
rect 18880 14492 18932 14501
rect 19248 14492 19300 14544
rect 19984 14492 20036 14544
rect 4160 14424 4212 14476
rect 4620 14424 4672 14476
rect 3148 14288 3200 14340
rect 3792 14288 3844 14340
rect 5540 14424 5592 14476
rect 6000 14424 6052 14476
rect 6828 14467 6880 14476
rect 6828 14433 6837 14467
rect 6837 14433 6871 14467
rect 6871 14433 6880 14467
rect 6828 14424 6880 14433
rect 9588 14424 9640 14476
rect 11796 14424 11848 14476
rect 14004 14424 14056 14476
rect 14740 14424 14792 14476
rect 20812 14467 20864 14476
rect 20812 14433 20821 14467
rect 20821 14433 20855 14467
rect 20855 14433 20864 14467
rect 20812 14424 20864 14433
rect 25044 14424 25096 14476
rect 6276 14356 6328 14408
rect 7932 14356 7984 14408
rect 8760 14356 8812 14408
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 18144 14356 18196 14408
rect 4252 14288 4304 14340
rect 5080 14288 5132 14340
rect 12624 14288 12676 14340
rect 18236 14288 18288 14340
rect 19248 14288 19300 14340
rect 24768 14331 24820 14340
rect 24768 14297 24777 14331
rect 24777 14297 24811 14331
rect 24811 14297 24820 14331
rect 24768 14288 24820 14297
rect 6092 14220 6144 14272
rect 6644 14263 6696 14272
rect 6644 14229 6653 14263
rect 6653 14229 6687 14263
rect 6687 14229 6696 14263
rect 6644 14220 6696 14229
rect 7472 14220 7524 14272
rect 8300 14220 8352 14272
rect 9312 14220 9364 14272
rect 10508 14263 10560 14272
rect 10508 14229 10517 14263
rect 10517 14229 10551 14263
rect 10551 14229 10560 14263
rect 10508 14220 10560 14229
rect 10784 14220 10836 14272
rect 12532 14220 12584 14272
rect 17408 14220 17460 14272
rect 19524 14220 19576 14272
rect 19800 14263 19852 14272
rect 19800 14229 19809 14263
rect 19809 14229 19843 14263
rect 19843 14229 19852 14263
rect 19800 14220 19852 14229
rect 20168 14220 20220 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1952 14016 2004 14068
rect 2228 14016 2280 14068
rect 3792 14016 3844 14068
rect 3976 14016 4028 14068
rect 4620 14016 4672 14068
rect 6276 14059 6328 14068
rect 1860 13880 1912 13932
rect 3056 13880 3108 13932
rect 6276 14025 6285 14059
rect 6285 14025 6319 14059
rect 6319 14025 6328 14059
rect 6276 14016 6328 14025
rect 8760 14016 8812 14068
rect 9680 14059 9732 14068
rect 9680 14025 9689 14059
rect 9689 14025 9723 14059
rect 9723 14025 9732 14059
rect 9680 14016 9732 14025
rect 10692 14016 10744 14068
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 14832 14016 14884 14068
rect 17408 14016 17460 14068
rect 18328 14016 18380 14068
rect 18880 14016 18932 14068
rect 19800 14016 19852 14068
rect 25044 14059 25096 14068
rect 25044 14025 25053 14059
rect 25053 14025 25087 14059
rect 25087 14025 25096 14059
rect 25044 14016 25096 14025
rect 5080 13948 5132 14000
rect 6000 13948 6052 14000
rect 8944 13948 8996 14000
rect 3976 13812 4028 13864
rect 5540 13855 5592 13864
rect 1676 13744 1728 13796
rect 1952 13744 2004 13796
rect 2320 13787 2372 13796
rect 2320 13753 2329 13787
rect 2329 13753 2363 13787
rect 2363 13753 2372 13787
rect 2320 13744 2372 13753
rect 2596 13719 2648 13728
rect 2596 13685 2605 13719
rect 2605 13685 2639 13719
rect 2639 13685 2648 13719
rect 2596 13676 2648 13685
rect 3516 13744 3568 13796
rect 3884 13787 3936 13796
rect 3884 13753 3893 13787
rect 3893 13753 3927 13787
rect 3927 13753 3936 13787
rect 3884 13744 3936 13753
rect 3424 13676 3476 13728
rect 5540 13821 5549 13855
rect 5549 13821 5583 13855
rect 5583 13821 5592 13855
rect 5540 13812 5592 13821
rect 6276 13812 6328 13864
rect 7564 13880 7616 13932
rect 9404 13923 9456 13932
rect 7472 13812 7524 13864
rect 7840 13812 7892 13864
rect 8300 13812 8352 13864
rect 6828 13744 6880 13796
rect 6184 13676 6236 13728
rect 7840 13676 7892 13728
rect 7932 13676 7984 13728
rect 8944 13812 8996 13864
rect 9404 13889 9413 13923
rect 9413 13889 9447 13923
rect 9447 13889 9456 13923
rect 9404 13880 9456 13889
rect 10140 13948 10192 14000
rect 10876 13948 10928 14000
rect 14004 13991 14056 14000
rect 14004 13957 14013 13991
rect 14013 13957 14047 13991
rect 14047 13957 14056 13991
rect 14004 13948 14056 13957
rect 20812 13948 20864 14000
rect 13268 13880 13320 13932
rect 14372 13880 14424 13932
rect 10508 13855 10560 13864
rect 10508 13821 10517 13855
rect 10517 13821 10551 13855
rect 10551 13821 10560 13855
rect 10508 13812 10560 13821
rect 15292 13880 15344 13932
rect 14832 13812 14884 13864
rect 18236 13880 18288 13932
rect 15936 13855 15988 13864
rect 15936 13821 15945 13855
rect 15945 13821 15979 13855
rect 15979 13821 15988 13855
rect 15936 13812 15988 13821
rect 16396 13812 16448 13864
rect 17776 13812 17828 13864
rect 20076 13855 20128 13864
rect 20076 13821 20085 13855
rect 20085 13821 20119 13855
rect 20119 13821 20128 13855
rect 20076 13812 20128 13821
rect 10968 13787 11020 13796
rect 10968 13753 10977 13787
rect 10977 13753 11011 13787
rect 11011 13753 11020 13787
rect 10968 13744 11020 13753
rect 12164 13744 12216 13796
rect 12532 13787 12584 13796
rect 12532 13753 12541 13787
rect 12541 13753 12575 13787
rect 12575 13753 12584 13787
rect 12532 13744 12584 13753
rect 12624 13787 12676 13796
rect 12624 13753 12633 13787
rect 12633 13753 12667 13787
rect 12667 13753 12676 13787
rect 12624 13744 12676 13753
rect 13544 13744 13596 13796
rect 18144 13787 18196 13796
rect 18144 13753 18153 13787
rect 18153 13753 18187 13787
rect 18187 13753 18196 13787
rect 18144 13744 18196 13753
rect 18328 13744 18380 13796
rect 14832 13676 14884 13728
rect 15476 13676 15528 13728
rect 15844 13676 15896 13728
rect 19432 13719 19484 13728
rect 19432 13685 19441 13719
rect 19441 13685 19475 13719
rect 19475 13685 19484 13719
rect 19432 13676 19484 13685
rect 26240 13744 26292 13796
rect 20076 13676 20128 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 3056 13472 3108 13524
rect 3424 13472 3476 13524
rect 7564 13515 7616 13524
rect 7564 13481 7573 13515
rect 7573 13481 7607 13515
rect 7607 13481 7616 13515
rect 7564 13472 7616 13481
rect 7748 13472 7800 13524
rect 8300 13472 8352 13524
rect 9680 13472 9732 13524
rect 12164 13472 12216 13524
rect 12624 13472 12676 13524
rect 12992 13472 13044 13524
rect 14372 13515 14424 13524
rect 1676 13447 1728 13456
rect 1676 13413 1685 13447
rect 1685 13413 1719 13447
rect 1719 13413 1728 13447
rect 1676 13404 1728 13413
rect 2228 13447 2280 13456
rect 2228 13413 2237 13447
rect 2237 13413 2271 13447
rect 2271 13413 2280 13447
rect 2228 13404 2280 13413
rect 4068 13447 4120 13456
rect 4068 13413 4077 13447
rect 4077 13413 4111 13447
rect 4111 13413 4120 13447
rect 4068 13404 4120 13413
rect 5080 13447 5132 13456
rect 5080 13413 5089 13447
rect 5089 13413 5123 13447
rect 5123 13413 5132 13447
rect 5080 13404 5132 13413
rect 3516 13336 3568 13388
rect 5540 13336 5592 13388
rect 6368 13336 6420 13388
rect 6460 13379 6512 13388
rect 6460 13345 6469 13379
rect 6469 13345 6503 13379
rect 6503 13345 6512 13379
rect 6460 13336 6512 13345
rect 7012 13336 7064 13388
rect 7932 13336 7984 13388
rect 9312 13404 9364 13456
rect 11612 13447 11664 13456
rect 11612 13413 11621 13447
rect 11621 13413 11655 13447
rect 11655 13413 11664 13447
rect 11612 13404 11664 13413
rect 14372 13481 14381 13515
rect 14381 13481 14415 13515
rect 14415 13481 14424 13515
rect 14372 13472 14424 13481
rect 15292 13472 15344 13524
rect 15936 13472 15988 13524
rect 17224 13515 17276 13524
rect 17224 13481 17233 13515
rect 17233 13481 17267 13515
rect 17267 13481 17276 13515
rect 17224 13472 17276 13481
rect 18052 13472 18104 13524
rect 19432 13472 19484 13524
rect 13544 13404 13596 13456
rect 16028 13447 16080 13456
rect 16028 13413 16037 13447
rect 16037 13413 16071 13447
rect 16071 13413 16080 13447
rect 16028 13404 16080 13413
rect 18236 13404 18288 13456
rect 18512 13447 18564 13456
rect 18512 13413 18521 13447
rect 18521 13413 18555 13447
rect 18555 13413 18564 13447
rect 18512 13404 18564 13413
rect 19248 13404 19300 13456
rect 10324 13336 10376 13388
rect 14096 13336 14148 13388
rect 15936 13336 15988 13388
rect 16396 13336 16448 13388
rect 17316 13379 17368 13388
rect 17316 13345 17325 13379
rect 17325 13345 17359 13379
rect 17359 13345 17368 13379
rect 17316 13336 17368 13345
rect 20812 13336 20864 13388
rect 23848 13336 23900 13388
rect 1400 13268 1452 13320
rect 4712 13268 4764 13320
rect 7472 13268 7524 13320
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 9036 13268 9088 13320
rect 9864 13311 9916 13320
rect 9864 13277 9873 13311
rect 9873 13277 9907 13311
rect 9907 13277 9916 13311
rect 9864 13268 9916 13277
rect 11888 13268 11940 13320
rect 13360 13311 13412 13320
rect 1492 13200 1544 13252
rect 4528 13200 4580 13252
rect 6184 13200 6236 13252
rect 3332 13132 3384 13184
rect 5080 13132 5132 13184
rect 7748 13132 7800 13184
rect 11796 13200 11848 13252
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 19432 13268 19484 13320
rect 16488 13200 16540 13252
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 10876 13175 10928 13184
rect 10876 13141 10885 13175
rect 10885 13141 10919 13175
rect 10919 13141 10928 13175
rect 10876 13132 10928 13141
rect 12532 13132 12584 13184
rect 18144 13175 18196 13184
rect 18144 13141 18153 13175
rect 18153 13141 18187 13175
rect 18187 13141 18196 13175
rect 18144 13132 18196 13141
rect 20168 13132 20220 13184
rect 24032 13132 24084 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1676 12928 1728 12980
rect 6368 12928 6420 12980
rect 10324 12971 10376 12980
rect 10324 12937 10333 12971
rect 10333 12937 10367 12971
rect 10367 12937 10376 12971
rect 10324 12928 10376 12937
rect 12900 12928 12952 12980
rect 12992 12928 13044 12980
rect 14280 12971 14332 12980
rect 14280 12937 14289 12971
rect 14289 12937 14323 12971
rect 14323 12937 14332 12971
rect 15936 12971 15988 12980
rect 14280 12928 14332 12937
rect 2228 12860 2280 12912
rect 6460 12860 6512 12912
rect 10784 12860 10836 12912
rect 20 12792 72 12844
rect 1492 12724 1544 12776
rect 4252 12792 4304 12844
rect 4436 12792 4488 12844
rect 10876 12792 10928 12844
rect 11796 12860 11848 12912
rect 14096 12860 14148 12912
rect 11612 12792 11664 12844
rect 13636 12792 13688 12844
rect 15936 12937 15945 12971
rect 15945 12937 15979 12971
rect 15979 12937 15988 12971
rect 15936 12928 15988 12937
rect 18512 12928 18564 12980
rect 19432 12971 19484 12980
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 20812 12928 20864 12980
rect 23848 12971 23900 12980
rect 23848 12937 23857 12971
rect 23857 12937 23891 12971
rect 23891 12937 23900 12971
rect 23848 12928 23900 12937
rect 17408 12860 17460 12912
rect 16488 12835 16540 12844
rect 16488 12801 16497 12835
rect 16497 12801 16531 12835
rect 16531 12801 16540 12835
rect 16488 12792 16540 12801
rect 18144 12835 18196 12844
rect 18144 12801 18153 12835
rect 18153 12801 18187 12835
rect 18187 12801 18196 12835
rect 18144 12792 18196 12801
rect 18972 12792 19024 12844
rect 19156 12792 19208 12844
rect 1860 12724 1912 12776
rect 4528 12767 4580 12776
rect 4528 12733 4537 12767
rect 4537 12733 4571 12767
rect 4571 12733 4580 12767
rect 4528 12724 4580 12733
rect 2136 12699 2188 12708
rect 2136 12665 2145 12699
rect 2145 12665 2179 12699
rect 2179 12665 2188 12699
rect 2136 12656 2188 12665
rect 3056 12699 3108 12708
rect 3056 12665 3065 12699
rect 3065 12665 3099 12699
rect 3099 12665 3108 12699
rect 3056 12656 3108 12665
rect 2872 12631 2924 12640
rect 2872 12597 2881 12631
rect 2881 12597 2915 12631
rect 2915 12597 2924 12631
rect 3884 12656 3936 12708
rect 2872 12588 2924 12597
rect 4252 12588 4304 12640
rect 4896 12724 4948 12776
rect 7196 12724 7248 12776
rect 8208 12767 8260 12776
rect 8208 12733 8217 12767
rect 8217 12733 8251 12767
rect 8251 12733 8260 12767
rect 8208 12724 8260 12733
rect 9036 12767 9088 12776
rect 7748 12656 7800 12708
rect 9036 12733 9045 12767
rect 9045 12733 9079 12767
rect 9079 12733 9088 12767
rect 9036 12724 9088 12733
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 6920 12588 6972 12640
rect 7932 12631 7984 12640
rect 7932 12597 7941 12631
rect 7941 12597 7975 12631
rect 7975 12597 7984 12631
rect 7932 12588 7984 12597
rect 8576 12588 8628 12640
rect 9128 12656 9180 12708
rect 17132 12767 17184 12776
rect 17132 12733 17141 12767
rect 17141 12733 17175 12767
rect 17175 12733 17184 12767
rect 17132 12724 17184 12733
rect 17960 12724 18012 12776
rect 12532 12699 12584 12708
rect 12532 12665 12541 12699
rect 12541 12665 12575 12699
rect 12575 12665 12584 12699
rect 12532 12656 12584 12665
rect 15016 12699 15068 12708
rect 10784 12631 10836 12640
rect 10784 12597 10793 12631
rect 10793 12597 10827 12631
rect 10827 12597 10836 12631
rect 10784 12588 10836 12597
rect 12256 12631 12308 12640
rect 12256 12597 12265 12631
rect 12265 12597 12299 12631
rect 12299 12597 12308 12631
rect 15016 12665 15025 12699
rect 15025 12665 15059 12699
rect 15059 12665 15068 12699
rect 15016 12656 15068 12665
rect 15660 12656 15712 12708
rect 18236 12699 18288 12708
rect 12256 12588 12308 12597
rect 13636 12588 13688 12640
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 17408 12631 17460 12640
rect 16212 12588 16264 12597
rect 17408 12597 17417 12631
rect 17417 12597 17451 12631
rect 17451 12597 17460 12631
rect 17408 12588 17460 12597
rect 17500 12588 17552 12640
rect 18236 12665 18245 12699
rect 18245 12665 18279 12699
rect 18279 12665 18288 12699
rect 18236 12656 18288 12665
rect 17960 12588 18012 12640
rect 20168 12631 20220 12640
rect 20168 12597 20177 12631
rect 20177 12597 20211 12631
rect 20211 12597 20220 12631
rect 20168 12588 20220 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1860 12427 1912 12436
rect 1860 12393 1869 12427
rect 1869 12393 1903 12427
rect 1903 12393 1912 12427
rect 1860 12384 1912 12393
rect 2872 12427 2924 12436
rect 2872 12393 2881 12427
rect 2881 12393 2915 12427
rect 2915 12393 2924 12427
rect 2872 12384 2924 12393
rect 3516 12427 3568 12436
rect 3516 12393 3525 12427
rect 3525 12393 3559 12427
rect 3559 12393 3568 12427
rect 3516 12384 3568 12393
rect 3792 12427 3844 12436
rect 3792 12393 3801 12427
rect 3801 12393 3835 12427
rect 3835 12393 3844 12427
rect 3792 12384 3844 12393
rect 4160 12427 4212 12436
rect 4160 12393 4169 12427
rect 4169 12393 4203 12427
rect 4203 12393 4212 12427
rect 4160 12384 4212 12393
rect 6000 12384 6052 12436
rect 8576 12384 8628 12436
rect 8944 12384 8996 12436
rect 9404 12427 9456 12436
rect 9404 12393 9413 12427
rect 9413 12393 9447 12427
rect 9447 12393 9456 12427
rect 9404 12384 9456 12393
rect 9772 12427 9824 12436
rect 9772 12393 9781 12427
rect 9781 12393 9815 12427
rect 9815 12393 9824 12427
rect 9772 12384 9824 12393
rect 11888 12427 11940 12436
rect 11888 12393 11897 12427
rect 11897 12393 11931 12427
rect 11931 12393 11940 12427
rect 11888 12384 11940 12393
rect 12072 12384 12124 12436
rect 13360 12384 13412 12436
rect 15016 12384 15068 12436
rect 15384 12384 15436 12436
rect 17500 12384 17552 12436
rect 17592 12384 17644 12436
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 2872 12291 2924 12300
rect 2872 12257 2881 12291
rect 2881 12257 2915 12291
rect 2915 12257 2924 12291
rect 2872 12248 2924 12257
rect 7380 12316 7432 12368
rect 4804 12291 4856 12300
rect 4804 12257 4813 12291
rect 4813 12257 4847 12291
rect 4847 12257 4856 12291
rect 4804 12248 4856 12257
rect 5080 12248 5132 12300
rect 5448 12180 5500 12232
rect 7656 12248 7708 12300
rect 8576 12291 8628 12300
rect 8576 12257 8585 12291
rect 8585 12257 8619 12291
rect 8619 12257 8628 12291
rect 8576 12248 8628 12257
rect 9864 12248 9916 12300
rect 8024 12180 8076 12232
rect 10048 12248 10100 12300
rect 10508 12291 10560 12300
rect 10508 12257 10517 12291
rect 10517 12257 10551 12291
rect 10551 12257 10560 12291
rect 10508 12248 10560 12257
rect 11520 12316 11572 12368
rect 15936 12316 15988 12368
rect 17776 12359 17828 12368
rect 17776 12325 17785 12359
rect 17785 12325 17819 12359
rect 17819 12325 17828 12359
rect 17776 12316 17828 12325
rect 17868 12359 17920 12368
rect 17868 12325 17877 12359
rect 17877 12325 17911 12359
rect 17911 12325 17920 12359
rect 17868 12316 17920 12325
rect 10968 12248 11020 12300
rect 13636 12291 13688 12300
rect 13636 12257 13645 12291
rect 13645 12257 13679 12291
rect 13679 12257 13688 12291
rect 13636 12248 13688 12257
rect 19248 12291 19300 12300
rect 19248 12257 19257 12291
rect 19257 12257 19291 12291
rect 19291 12257 19300 12291
rect 19248 12248 19300 12257
rect 19432 12248 19484 12300
rect 21456 12248 21508 12300
rect 23848 12248 23900 12300
rect 11428 12180 11480 12232
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 12256 12180 12308 12232
rect 4620 12112 4672 12164
rect 4712 12112 4764 12164
rect 8668 12155 8720 12164
rect 8668 12121 8677 12155
rect 8677 12121 8711 12155
rect 8711 12121 8720 12155
rect 8668 12112 8720 12121
rect 9864 12112 9916 12164
rect 10508 12112 10560 12164
rect 12624 12155 12676 12164
rect 12624 12121 12633 12155
rect 12633 12121 12667 12155
rect 12667 12121 12676 12155
rect 12624 12112 12676 12121
rect 16580 12112 16632 12164
rect 18512 12112 18564 12164
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 6000 12044 6052 12096
rect 6460 12044 6512 12096
rect 8208 12044 8260 12096
rect 10416 12044 10468 12096
rect 16948 12044 17000 12096
rect 17224 12087 17276 12096
rect 17224 12053 17233 12087
rect 17233 12053 17267 12087
rect 17267 12053 17276 12087
rect 17224 12044 17276 12053
rect 18420 12044 18472 12096
rect 18788 12087 18840 12096
rect 18788 12053 18797 12087
rect 18797 12053 18831 12087
rect 18831 12053 18840 12087
rect 18788 12044 18840 12053
rect 18880 12044 18932 12096
rect 24124 12044 24176 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 4896 11840 4948 11892
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 7932 11840 7984 11892
rect 9864 11883 9916 11892
rect 9864 11849 9873 11883
rect 9873 11849 9907 11883
rect 9907 11849 9916 11883
rect 9864 11840 9916 11849
rect 10784 11840 10836 11892
rect 13636 11883 13688 11892
rect 2136 11772 2188 11824
rect 3056 11704 3108 11756
rect 7656 11772 7708 11824
rect 7840 11772 7892 11824
rect 12348 11772 12400 11824
rect 13636 11849 13645 11883
rect 13645 11849 13679 11883
rect 13679 11849 13688 11883
rect 13636 11840 13688 11849
rect 15384 11883 15436 11892
rect 15384 11849 15393 11883
rect 15393 11849 15427 11883
rect 15427 11849 15436 11883
rect 15384 11840 15436 11849
rect 18788 11840 18840 11892
rect 23848 11883 23900 11892
rect 23848 11849 23857 11883
rect 23857 11849 23891 11883
rect 23891 11849 23900 11883
rect 23848 11840 23900 11849
rect 24768 11883 24820 11892
rect 24768 11849 24777 11883
rect 24777 11849 24811 11883
rect 24811 11849 24820 11883
rect 24768 11840 24820 11849
rect 7380 11747 7432 11756
rect 1216 11636 1268 11688
rect 2780 11636 2832 11688
rect 4160 11636 4212 11688
rect 4712 11679 4764 11688
rect 4712 11645 4721 11679
rect 4721 11645 4755 11679
rect 4755 11645 4764 11679
rect 4712 11636 4764 11645
rect 4896 11679 4948 11688
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 5448 11679 5500 11688
rect 5448 11645 5457 11679
rect 5457 11645 5491 11679
rect 5491 11645 5500 11679
rect 5448 11636 5500 11645
rect 5540 11636 5592 11688
rect 6000 11636 6052 11688
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 8208 11679 8260 11688
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 9036 11704 9088 11756
rect 10416 11747 10468 11756
rect 10416 11713 10425 11747
rect 10425 11713 10459 11747
rect 10459 11713 10468 11747
rect 10416 11704 10468 11713
rect 12256 11747 12308 11756
rect 12256 11713 12265 11747
rect 12265 11713 12299 11747
rect 12299 11713 12308 11747
rect 12256 11704 12308 11713
rect 13360 11704 13412 11756
rect 14832 11704 14884 11756
rect 15660 11704 15712 11756
rect 17224 11704 17276 11756
rect 18972 11772 19024 11824
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 9404 11679 9456 11688
rect 2596 11611 2648 11620
rect 2596 11577 2605 11611
rect 2605 11577 2639 11611
rect 2639 11577 2648 11611
rect 2596 11568 2648 11577
rect 3516 11568 3568 11620
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 3608 11500 3660 11509
rect 5080 11500 5132 11552
rect 5172 11500 5224 11552
rect 6092 11568 6144 11620
rect 7748 11568 7800 11620
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 15936 11679 15988 11688
rect 15936 11645 15945 11679
rect 15945 11645 15979 11679
rect 15979 11645 15988 11679
rect 15936 11636 15988 11645
rect 18972 11636 19024 11688
rect 16856 11568 16908 11620
rect 17316 11568 17368 11620
rect 17408 11568 17460 11620
rect 18236 11611 18288 11620
rect 7380 11500 7432 11552
rect 10784 11543 10836 11552
rect 10784 11509 10793 11543
rect 10793 11509 10827 11543
rect 10827 11509 10836 11543
rect 10784 11500 10836 11509
rect 11336 11543 11388 11552
rect 11336 11509 11345 11543
rect 11345 11509 11379 11543
rect 11379 11509 11388 11543
rect 11336 11500 11388 11509
rect 11520 11500 11572 11552
rect 13912 11543 13964 11552
rect 13912 11509 13921 11543
rect 13921 11509 13955 11543
rect 13955 11509 13964 11543
rect 13912 11500 13964 11509
rect 16212 11500 16264 11552
rect 17868 11500 17920 11552
rect 18236 11577 18245 11611
rect 18245 11577 18279 11611
rect 18279 11577 18288 11611
rect 18236 11568 18288 11577
rect 18512 11568 18564 11620
rect 24124 11636 24176 11688
rect 25504 11568 25556 11620
rect 21456 11543 21508 11552
rect 21456 11509 21465 11543
rect 21465 11509 21499 11543
rect 21499 11509 21508 11543
rect 21456 11500 21508 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1400 11296 1452 11348
rect 1860 11296 1912 11348
rect 2872 11339 2924 11348
rect 2872 11305 2881 11339
rect 2881 11305 2915 11339
rect 2915 11305 2924 11339
rect 2872 11296 2924 11305
rect 3608 11228 3660 11280
rect 4896 11296 4948 11348
rect 5172 11296 5224 11348
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 7656 11296 7708 11348
rect 10048 11296 10100 11348
rect 10968 11339 11020 11348
rect 10968 11305 10977 11339
rect 10977 11305 11011 11339
rect 11011 11305 11020 11339
rect 10968 11296 11020 11305
rect 11428 11339 11480 11348
rect 11428 11305 11437 11339
rect 11437 11305 11471 11339
rect 11471 11305 11480 11339
rect 11428 11296 11480 11305
rect 12348 11296 12400 11348
rect 16580 11339 16632 11348
rect 16580 11305 16589 11339
rect 16589 11305 16623 11339
rect 16623 11305 16632 11339
rect 16580 11296 16632 11305
rect 18236 11296 18288 11348
rect 19432 11296 19484 11348
rect 24768 11339 24820 11348
rect 24768 11305 24777 11339
rect 24777 11305 24811 11339
rect 24811 11305 24820 11339
rect 24768 11296 24820 11305
rect 1768 11203 1820 11212
rect 1768 11169 1777 11203
rect 1777 11169 1811 11203
rect 1811 11169 1820 11203
rect 1768 11160 1820 11169
rect 3424 11160 3476 11212
rect 4620 11228 4672 11280
rect 6644 11271 6696 11280
rect 6644 11237 6653 11271
rect 6653 11237 6687 11271
rect 6687 11237 6696 11271
rect 6644 11228 6696 11237
rect 7012 11271 7064 11280
rect 7012 11237 7021 11271
rect 7021 11237 7055 11271
rect 7055 11237 7064 11271
rect 7012 11228 7064 11237
rect 7564 11271 7616 11280
rect 7564 11237 7573 11271
rect 7573 11237 7607 11271
rect 7607 11237 7616 11271
rect 7564 11228 7616 11237
rect 7748 11228 7800 11280
rect 11336 11228 11388 11280
rect 5172 11160 5224 11212
rect 8116 11160 8168 11212
rect 8576 11203 8628 11212
rect 8576 11169 8620 11203
rect 8620 11169 8628 11203
rect 8576 11160 8628 11169
rect 9220 11160 9272 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 10416 11203 10468 11212
rect 10416 11169 10425 11203
rect 10425 11169 10459 11203
rect 10459 11169 10468 11203
rect 10416 11160 10468 11169
rect 14188 11228 14240 11280
rect 15936 11228 15988 11280
rect 16948 11228 17000 11280
rect 17776 11228 17828 11280
rect 19064 11228 19116 11280
rect 19800 11228 19852 11280
rect 14004 11160 14056 11212
rect 20260 11160 20312 11212
rect 21364 11203 21416 11212
rect 21364 11169 21373 11203
rect 21373 11169 21407 11203
rect 21407 11169 21416 11203
rect 21364 11160 21416 11169
rect 24032 11160 24084 11212
rect 24676 11160 24728 11212
rect 4712 11092 4764 11144
rect 6092 11092 6144 11144
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 11796 11092 11848 11144
rect 3700 11024 3752 11076
rect 11428 11024 11480 11076
rect 12624 11092 12676 11144
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 17132 11135 17184 11144
rect 17132 11101 17141 11135
rect 17141 11101 17175 11135
rect 17175 11101 17184 11135
rect 18696 11135 18748 11144
rect 17132 11092 17184 11101
rect 17316 11024 17368 11076
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 1676 10999 1728 11008
rect 1676 10965 1685 10999
rect 1685 10965 1719 10999
rect 1719 10965 1728 10999
rect 1676 10956 1728 10965
rect 5356 10956 5408 11008
rect 6000 10999 6052 11008
rect 6000 10965 6009 10999
rect 6009 10965 6043 10999
rect 6043 10965 6052 10999
rect 6000 10956 6052 10965
rect 8944 10956 8996 11008
rect 9128 10999 9180 11008
rect 9128 10965 9137 10999
rect 9137 10965 9171 10999
rect 9171 10965 9180 10999
rect 9128 10956 9180 10965
rect 12716 10956 12768 11008
rect 14832 10956 14884 11008
rect 16212 10999 16264 11008
rect 16212 10965 16221 10999
rect 16221 10965 16255 10999
rect 16255 10965 16264 10999
rect 16212 10956 16264 10965
rect 16856 10999 16908 11008
rect 16856 10965 16865 10999
rect 16865 10965 16899 10999
rect 16899 10965 16908 10999
rect 16856 10956 16908 10965
rect 17868 10956 17920 11008
rect 19156 10956 19208 11008
rect 22192 10956 22244 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1768 10752 1820 10804
rect 2412 10752 2464 10804
rect 1308 10616 1360 10668
rect 1492 10591 1544 10600
rect 1492 10557 1501 10591
rect 1501 10557 1535 10591
rect 1535 10557 1544 10591
rect 1492 10548 1544 10557
rect 1676 10548 1728 10600
rect 4252 10752 4304 10804
rect 5448 10752 5500 10804
rect 6920 10752 6972 10804
rect 8208 10795 8260 10804
rect 8208 10761 8217 10795
rect 8217 10761 8251 10795
rect 8251 10761 8260 10795
rect 8208 10752 8260 10761
rect 8576 10795 8628 10804
rect 8576 10761 8585 10795
rect 8585 10761 8619 10795
rect 8619 10761 8628 10795
rect 8576 10752 8628 10761
rect 11336 10752 11388 10804
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 15936 10795 15988 10804
rect 15936 10761 15945 10795
rect 15945 10761 15979 10795
rect 15979 10761 15988 10795
rect 15936 10752 15988 10761
rect 16948 10752 17000 10804
rect 18696 10752 18748 10804
rect 19800 10795 19852 10804
rect 19800 10761 19809 10795
rect 19809 10761 19843 10795
rect 19843 10761 19852 10795
rect 19800 10752 19852 10761
rect 21364 10795 21416 10804
rect 21364 10761 21373 10795
rect 21373 10761 21407 10795
rect 21407 10761 21416 10795
rect 21364 10752 21416 10761
rect 24676 10795 24728 10804
rect 24676 10761 24685 10795
rect 24685 10761 24719 10795
rect 24719 10761 24728 10795
rect 24676 10752 24728 10761
rect 4712 10727 4764 10736
rect 4712 10693 4721 10727
rect 4721 10693 4755 10727
rect 4755 10693 4764 10727
rect 4712 10684 4764 10693
rect 7564 10684 7616 10736
rect 7656 10684 7708 10736
rect 14188 10684 14240 10736
rect 19064 10727 19116 10736
rect 19064 10693 19073 10727
rect 19073 10693 19107 10727
rect 19107 10693 19116 10727
rect 19064 10684 19116 10693
rect 3700 10659 3752 10668
rect 3700 10625 3709 10659
rect 3709 10625 3743 10659
rect 3743 10625 3752 10659
rect 3700 10616 3752 10625
rect 3884 10616 3936 10668
rect 3424 10480 3476 10532
rect 3700 10480 3752 10532
rect 7012 10616 7064 10668
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 12716 10616 12768 10668
rect 6000 10548 6052 10600
rect 7104 10548 7156 10600
rect 5264 10523 5316 10532
rect 5264 10489 5273 10523
rect 5273 10489 5307 10523
rect 5307 10489 5316 10523
rect 5264 10480 5316 10489
rect 5356 10523 5408 10532
rect 5356 10489 5365 10523
rect 5365 10489 5399 10523
rect 5399 10489 5408 10523
rect 9128 10548 9180 10600
rect 10416 10548 10468 10600
rect 11336 10591 11388 10600
rect 11336 10557 11345 10591
rect 11345 10557 11379 10591
rect 11379 10557 11388 10591
rect 11336 10548 11388 10557
rect 13268 10548 13320 10600
rect 5356 10480 5408 10489
rect 3516 10412 3568 10464
rect 4620 10412 4672 10464
rect 9036 10480 9088 10532
rect 9680 10523 9732 10532
rect 9680 10489 9689 10523
rect 9689 10489 9723 10523
rect 9723 10489 9732 10523
rect 9680 10480 9732 10489
rect 14832 10616 14884 10668
rect 15660 10659 15712 10668
rect 15660 10625 15669 10659
rect 15669 10625 15703 10659
rect 15703 10625 15712 10659
rect 15660 10616 15712 10625
rect 7012 10412 7064 10464
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 11980 10412 12032 10464
rect 12808 10412 12860 10464
rect 16212 10480 16264 10532
rect 18420 10659 18472 10668
rect 18420 10625 18429 10659
rect 18429 10625 18463 10659
rect 18463 10625 18472 10659
rect 18420 10616 18472 10625
rect 19432 10548 19484 10600
rect 18236 10523 18288 10532
rect 18236 10489 18245 10523
rect 18245 10489 18279 10523
rect 18279 10489 18288 10523
rect 18236 10480 18288 10489
rect 14004 10455 14056 10464
rect 14004 10421 14013 10455
rect 14013 10421 14047 10455
rect 14047 10421 14056 10455
rect 14004 10412 14056 10421
rect 17960 10412 18012 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1492 10208 1544 10260
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 4436 10208 4488 10260
rect 5356 10208 5408 10260
rect 6092 10251 6144 10260
rect 6092 10217 6101 10251
rect 6101 10217 6135 10251
rect 6135 10217 6144 10251
rect 6092 10208 6144 10217
rect 7104 10251 7156 10260
rect 7104 10217 7113 10251
rect 7113 10217 7147 10251
rect 7147 10217 7156 10251
rect 7104 10208 7156 10217
rect 9036 10251 9088 10260
rect 9036 10217 9045 10251
rect 9045 10217 9079 10251
rect 9079 10217 9088 10251
rect 9036 10208 9088 10217
rect 9680 10208 9732 10260
rect 11336 10208 11388 10260
rect 11796 10251 11848 10260
rect 11796 10217 11805 10251
rect 11805 10217 11839 10251
rect 11839 10217 11848 10251
rect 11796 10208 11848 10217
rect 13912 10251 13964 10260
rect 13912 10217 13921 10251
rect 13921 10217 13955 10251
rect 13955 10217 13964 10251
rect 13912 10208 13964 10217
rect 15936 10251 15988 10260
rect 15936 10217 15945 10251
rect 15945 10217 15979 10251
rect 15979 10217 15988 10251
rect 15936 10208 15988 10217
rect 16856 10208 16908 10260
rect 17132 10251 17184 10260
rect 17132 10217 17141 10251
rect 17141 10217 17175 10251
rect 17175 10217 17184 10251
rect 17132 10208 17184 10217
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 17960 10208 18012 10260
rect 18328 10208 18380 10260
rect 19064 10208 19116 10260
rect 2228 10140 2280 10192
rect 1308 10072 1360 10124
rect 2872 10072 2924 10124
rect 4988 10140 5040 10192
rect 5264 10140 5316 10192
rect 8300 10140 8352 10192
rect 8392 10140 8444 10192
rect 10968 10140 11020 10192
rect 12348 10140 12400 10192
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 5080 10115 5132 10124
rect 5080 10081 5089 10115
rect 5089 10081 5123 10115
rect 5123 10081 5132 10115
rect 5080 10072 5132 10081
rect 4988 10004 5040 10056
rect 7104 10072 7156 10124
rect 8116 10115 8168 10124
rect 8116 10081 8125 10115
rect 8125 10081 8159 10115
rect 8159 10081 8168 10115
rect 8116 10072 8168 10081
rect 8208 10072 8260 10124
rect 13728 10072 13780 10124
rect 14280 10140 14332 10192
rect 18696 10140 18748 10192
rect 14004 10072 14056 10124
rect 10140 10004 10192 10056
rect 12072 10047 12124 10056
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 15384 10004 15436 10056
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 19248 10004 19300 10056
rect 3976 9936 4028 9988
rect 4160 9936 4212 9988
rect 5264 9936 5316 9988
rect 5540 9868 5592 9920
rect 6736 9868 6788 9920
rect 7656 9868 7708 9920
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 13360 9868 13412 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2412 9707 2464 9716
rect 2412 9673 2421 9707
rect 2421 9673 2455 9707
rect 2455 9673 2464 9707
rect 2412 9664 2464 9673
rect 8208 9664 8260 9716
rect 1308 9528 1360 9580
rect 1860 9571 1912 9580
rect 1860 9537 1869 9571
rect 1869 9537 1903 9571
rect 1903 9537 1912 9571
rect 1860 9528 1912 9537
rect 6736 9596 6788 9648
rect 8300 9596 8352 9648
rect 8944 9664 8996 9716
rect 12072 9664 12124 9716
rect 13728 9707 13780 9716
rect 13728 9673 13737 9707
rect 13737 9673 13771 9707
rect 13771 9673 13780 9707
rect 13728 9664 13780 9673
rect 13912 9664 13964 9716
rect 15936 9664 15988 9716
rect 18328 9664 18380 9716
rect 19248 9707 19300 9716
rect 19248 9673 19257 9707
rect 19257 9673 19291 9707
rect 19291 9673 19300 9707
rect 19248 9664 19300 9673
rect 9128 9639 9180 9648
rect 9128 9605 9137 9639
rect 9137 9605 9171 9639
rect 9171 9605 9180 9639
rect 9128 9596 9180 9605
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 2412 9460 2464 9512
rect 3700 9460 3752 9512
rect 7840 9528 7892 9580
rect 3976 9460 4028 9512
rect 4988 9460 5040 9512
rect 5264 9503 5316 9512
rect 5264 9469 5273 9503
rect 5273 9469 5307 9503
rect 5307 9469 5316 9503
rect 5264 9460 5316 9469
rect 6000 9460 6052 9512
rect 5540 9392 5592 9444
rect 6736 9392 6788 9444
rect 9680 9571 9732 9580
rect 9680 9537 9689 9571
rect 9689 9537 9723 9571
rect 9723 9537 9732 9571
rect 9680 9528 9732 9537
rect 13268 9528 13320 9580
rect 7748 9435 7800 9444
rect 7748 9401 7757 9435
rect 7757 9401 7791 9435
rect 7791 9401 7800 9435
rect 7748 9392 7800 9401
rect 8392 9392 8444 9444
rect 12348 9460 12400 9512
rect 15936 9503 15988 9512
rect 15936 9469 15945 9503
rect 15945 9469 15979 9503
rect 15979 9469 15988 9503
rect 15936 9460 15988 9469
rect 17224 9528 17276 9580
rect 18512 9571 18564 9580
rect 18512 9537 18521 9571
rect 18521 9537 18555 9571
rect 18555 9537 18564 9571
rect 18512 9528 18564 9537
rect 10048 9392 10100 9444
rect 4528 9324 4580 9376
rect 5080 9324 5132 9376
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 8852 9367 8904 9376
rect 8852 9333 8861 9367
rect 8861 9333 8895 9367
rect 8895 9333 8904 9367
rect 8852 9324 8904 9333
rect 10968 9367 11020 9376
rect 10968 9333 10977 9367
rect 10977 9333 11011 9367
rect 11011 9333 11020 9367
rect 10968 9324 11020 9333
rect 12440 9324 12492 9376
rect 12624 9435 12676 9444
rect 12624 9401 12633 9435
rect 12633 9401 12667 9435
rect 12667 9401 12676 9435
rect 12624 9392 12676 9401
rect 13360 9392 13412 9444
rect 14188 9435 14240 9444
rect 14188 9401 14197 9435
rect 14197 9401 14231 9435
rect 14231 9401 14240 9435
rect 17684 9460 17736 9512
rect 14188 9392 14240 9401
rect 18236 9435 18288 9444
rect 18236 9401 18245 9435
rect 18245 9401 18279 9435
rect 18279 9401 18288 9435
rect 18236 9392 18288 9401
rect 18328 9435 18380 9444
rect 18328 9401 18337 9435
rect 18337 9401 18371 9435
rect 18371 9401 18380 9435
rect 18328 9392 18380 9401
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2872 9163 2924 9172
rect 2872 9129 2881 9163
rect 2881 9129 2915 9163
rect 2915 9129 2924 9163
rect 2872 9120 2924 9129
rect 3332 9120 3384 9172
rect 3700 9163 3752 9172
rect 3700 9129 3709 9163
rect 3709 9129 3743 9163
rect 3743 9129 3752 9163
rect 3700 9120 3752 9129
rect 4068 9120 4120 9172
rect 1400 9095 1452 9104
rect 1400 9061 1409 9095
rect 1409 9061 1443 9095
rect 1443 9061 1452 9095
rect 1400 9052 1452 9061
rect 1492 9027 1544 9036
rect 1492 8993 1501 9027
rect 1501 8993 1535 9027
rect 1535 8993 1544 9027
rect 1492 8984 1544 8993
rect 2964 9027 3016 9036
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 2964 8984 3016 8993
rect 6644 9120 6696 9172
rect 7104 9163 7156 9172
rect 7104 9129 7113 9163
rect 7113 9129 7147 9163
rect 7147 9129 7156 9163
rect 7104 9120 7156 9129
rect 8116 9120 8168 9172
rect 11980 9163 12032 9172
rect 5540 9052 5592 9104
rect 6000 9052 6052 9104
rect 4528 8984 4580 9036
rect 6092 9027 6144 9036
rect 6092 8993 6101 9027
rect 6101 8993 6135 9027
rect 6135 8993 6144 9027
rect 6092 8984 6144 8993
rect 7932 9052 7984 9104
rect 8208 9052 8260 9104
rect 8300 9027 8352 9036
rect 8300 8993 8309 9027
rect 8309 8993 8343 9027
rect 8343 8993 8352 9027
rect 8300 8984 8352 8993
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 6184 8891 6236 8900
rect 5080 8780 5132 8832
rect 5264 8780 5316 8832
rect 6184 8857 6193 8891
rect 6193 8857 6227 8891
rect 6227 8857 6236 8891
rect 6184 8848 6236 8857
rect 11980 9129 11989 9163
rect 11989 9129 12023 9163
rect 12023 9129 12032 9163
rect 11980 9120 12032 9129
rect 12348 9120 12400 9172
rect 12624 9120 12676 9172
rect 14188 9120 14240 9172
rect 15936 9120 15988 9172
rect 18236 9120 18288 9172
rect 10048 9052 10100 9104
rect 11520 9052 11572 9104
rect 13912 9052 13964 9104
rect 14004 9052 14056 9104
rect 10140 8984 10192 9036
rect 11244 8984 11296 9036
rect 14556 8984 14608 9036
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 16856 9052 16908 9104
rect 17868 9095 17920 9104
rect 17868 9061 17877 9095
rect 17877 9061 17911 9095
rect 17911 9061 17920 9095
rect 17868 9052 17920 9061
rect 16304 8984 16356 9036
rect 18788 8984 18840 9036
rect 10692 8916 10744 8968
rect 13636 8916 13688 8968
rect 17224 8959 17276 8968
rect 14096 8848 14148 8900
rect 15752 8848 15804 8900
rect 17224 8925 17233 8959
rect 17233 8925 17267 8959
rect 17267 8925 17276 8959
rect 17224 8916 17276 8925
rect 17316 8916 17368 8968
rect 6000 8823 6052 8832
rect 6000 8789 6009 8823
rect 6009 8789 6043 8823
rect 6043 8789 6052 8823
rect 6000 8780 6052 8789
rect 10600 8823 10652 8832
rect 10600 8789 10609 8823
rect 10609 8789 10643 8823
rect 10643 8789 10652 8823
rect 10600 8780 10652 8789
rect 10968 8823 11020 8832
rect 10968 8789 10977 8823
rect 10977 8789 11011 8823
rect 11011 8789 11020 8823
rect 10968 8780 11020 8789
rect 15384 8780 15436 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 3056 8576 3108 8628
rect 6092 8619 6144 8628
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 7748 8576 7800 8628
rect 8300 8576 8352 8628
rect 13544 8576 13596 8628
rect 13912 8576 13964 8628
rect 15292 8619 15344 8628
rect 15292 8585 15301 8619
rect 15301 8585 15335 8619
rect 15335 8585 15344 8619
rect 15292 8576 15344 8585
rect 16856 8576 16908 8628
rect 2964 8440 3016 8492
rect 5356 8440 5408 8492
rect 5540 8440 5592 8492
rect 6000 8440 6052 8492
rect 6184 8440 6236 8492
rect 8208 8508 8260 8560
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 8576 8440 8628 8492
rect 10876 8483 10928 8492
rect 10876 8449 10885 8483
rect 10885 8449 10919 8483
rect 10919 8449 10928 8483
rect 10876 8440 10928 8449
rect 11520 8483 11572 8492
rect 11520 8449 11529 8483
rect 11529 8449 11563 8483
rect 11563 8449 11572 8483
rect 11520 8440 11572 8449
rect 6644 8372 6696 8424
rect 8116 8372 8168 8424
rect 9680 8372 9732 8424
rect 12716 8508 12768 8560
rect 17040 8508 17092 8560
rect 19340 8440 19392 8492
rect 15752 8415 15804 8424
rect 8392 8304 8444 8356
rect 10140 8304 10192 8356
rect 10600 8347 10652 8356
rect 10600 8313 10609 8347
rect 10609 8313 10643 8347
rect 10643 8313 10652 8347
rect 10600 8304 10652 8313
rect 10968 8304 11020 8356
rect 12256 8304 12308 8356
rect 848 8236 900 8288
rect 1492 8236 1544 8288
rect 3976 8279 4028 8288
rect 3976 8245 3985 8279
rect 3985 8245 4019 8279
rect 4019 8245 4028 8279
rect 3976 8236 4028 8245
rect 4528 8279 4580 8288
rect 4528 8245 4537 8279
rect 4537 8245 4571 8279
rect 4571 8245 4580 8279
rect 4528 8236 4580 8245
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 15752 8381 15761 8415
rect 15761 8381 15795 8415
rect 15795 8381 15804 8415
rect 15752 8372 15804 8381
rect 16304 8415 16356 8424
rect 16304 8381 16313 8415
rect 16313 8381 16347 8415
rect 16347 8381 16356 8415
rect 16304 8372 16356 8381
rect 17868 8415 17920 8424
rect 17868 8381 17877 8415
rect 17877 8381 17911 8415
rect 17911 8381 17920 8415
rect 17868 8372 17920 8381
rect 12716 8347 12768 8356
rect 12716 8313 12725 8347
rect 12725 8313 12759 8347
rect 12759 8313 12768 8347
rect 12716 8304 12768 8313
rect 13360 8347 13412 8356
rect 13360 8313 13369 8347
rect 13369 8313 13403 8347
rect 13403 8313 13412 8347
rect 13360 8304 13412 8313
rect 14280 8347 14332 8356
rect 14280 8313 14289 8347
rect 14289 8313 14323 8347
rect 14323 8313 14332 8347
rect 14280 8304 14332 8313
rect 15936 8236 15988 8288
rect 18788 8279 18840 8288
rect 18788 8245 18797 8279
rect 18797 8245 18831 8279
rect 18831 8245 18840 8279
rect 18788 8236 18840 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 6184 8032 6236 8084
rect 7932 8075 7984 8084
rect 7932 8041 7941 8075
rect 7941 8041 7975 8075
rect 7975 8041 7984 8075
rect 7932 8032 7984 8041
rect 8576 8032 8628 8084
rect 11244 8075 11296 8084
rect 11244 8041 11253 8075
rect 11253 8041 11287 8075
rect 11287 8041 11296 8075
rect 11244 8032 11296 8041
rect 13636 8075 13688 8084
rect 13636 8041 13645 8075
rect 13645 8041 13679 8075
rect 13679 8041 13688 8075
rect 13636 8032 13688 8041
rect 15384 8075 15436 8084
rect 15384 8041 15393 8075
rect 15393 8041 15427 8075
rect 15427 8041 15436 8075
rect 15384 8032 15436 8041
rect 16304 8075 16356 8084
rect 16304 8041 16313 8075
rect 16313 8041 16347 8075
rect 16347 8041 16356 8075
rect 16304 8032 16356 8041
rect 17224 8075 17276 8084
rect 17224 8041 17233 8075
rect 17233 8041 17267 8075
rect 17267 8041 17276 8075
rect 17224 8032 17276 8041
rect 8116 7964 8168 8016
rect 8208 8007 8260 8016
rect 8208 7973 8217 8007
rect 8217 7973 8251 8007
rect 8251 7973 8260 8007
rect 8208 7964 8260 7973
rect 10048 7964 10100 8016
rect 12256 7964 12308 8016
rect 13360 8007 13412 8016
rect 13360 7973 13369 8007
rect 13369 7973 13403 8007
rect 13403 7973 13412 8007
rect 13360 7964 13412 7973
rect 13820 7964 13872 8016
rect 4528 7939 4580 7948
rect 4528 7905 4537 7939
rect 4537 7905 4571 7939
rect 4571 7905 4580 7939
rect 4528 7896 4580 7905
rect 5448 7896 5500 7948
rect 4988 7828 5040 7880
rect 6644 7896 6696 7948
rect 14188 7939 14240 7948
rect 14188 7905 14197 7939
rect 14197 7905 14231 7939
rect 14231 7905 14240 7939
rect 14188 7896 14240 7905
rect 15660 7896 15712 7948
rect 15844 7939 15896 7948
rect 15844 7905 15853 7939
rect 15853 7905 15887 7939
rect 15887 7905 15896 7939
rect 15844 7896 15896 7905
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 8760 7871 8812 7880
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 10048 7871 10100 7880
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 11888 7828 11940 7880
rect 5540 7760 5592 7812
rect 6460 7692 6512 7744
rect 10968 7735 11020 7744
rect 10968 7701 10977 7735
rect 10977 7701 11011 7735
rect 11011 7701 11020 7735
rect 10968 7692 11020 7701
rect 12716 7692 12768 7744
rect 14280 7692 14332 7744
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 5448 7488 5500 7540
rect 7012 7531 7064 7540
rect 7012 7497 7021 7531
rect 7021 7497 7055 7531
rect 7055 7497 7064 7531
rect 7012 7488 7064 7497
rect 8208 7488 8260 7540
rect 1860 7327 1912 7336
rect 1860 7293 1869 7327
rect 1869 7293 1903 7327
rect 1903 7293 1912 7327
rect 1860 7284 1912 7293
rect 5080 7284 5132 7336
rect 6736 7284 6788 7336
rect 5448 7216 5500 7268
rect 5724 7216 5776 7268
rect 6000 7216 6052 7268
rect 8392 7488 8444 7540
rect 8852 7488 8904 7540
rect 10324 7488 10376 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 12256 7531 12308 7540
rect 12256 7497 12265 7531
rect 12265 7497 12299 7531
rect 12299 7497 12308 7531
rect 12256 7488 12308 7497
rect 12440 7488 12492 7540
rect 12716 7488 12768 7540
rect 15844 7488 15896 7540
rect 9956 7463 10008 7472
rect 9956 7429 9965 7463
rect 9965 7429 9999 7463
rect 9999 7429 10008 7463
rect 9956 7420 10008 7429
rect 8760 7352 8812 7404
rect 10876 7352 10928 7404
rect 9772 7284 9824 7336
rect 13176 7420 13228 7472
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 9864 7216 9916 7268
rect 4528 7191 4580 7200
rect 4528 7157 4537 7191
rect 4537 7157 4571 7191
rect 4571 7157 4580 7191
rect 4528 7148 4580 7157
rect 4988 7191 5040 7200
rect 4988 7157 4997 7191
rect 4997 7157 5031 7191
rect 5031 7157 5040 7191
rect 4988 7148 5040 7157
rect 9312 7191 9364 7200
rect 9312 7157 9321 7191
rect 9321 7157 9355 7191
rect 9355 7157 9364 7191
rect 9312 7148 9364 7157
rect 10324 7259 10376 7268
rect 10324 7225 10333 7259
rect 10333 7225 10367 7259
rect 10367 7225 10376 7259
rect 10324 7216 10376 7225
rect 12900 7216 12952 7268
rect 15752 7284 15804 7336
rect 15660 7191 15712 7200
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 3976 6944 4028 6996
rect 9772 6944 9824 6996
rect 10140 6987 10192 6996
rect 10140 6953 10149 6987
rect 10149 6953 10183 6987
rect 10183 6953 10192 6987
rect 10140 6944 10192 6953
rect 14648 6944 14700 6996
rect 5448 6876 5500 6928
rect 8116 6876 8168 6928
rect 10048 6876 10100 6928
rect 10968 6876 11020 6928
rect 11336 6919 11388 6928
rect 11336 6885 11345 6919
rect 11345 6885 11379 6919
rect 11379 6885 11388 6919
rect 11336 6876 11388 6885
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 5356 6808 5408 6860
rect 5724 6851 5776 6860
rect 5724 6817 5733 6851
rect 5733 6817 5767 6851
rect 5767 6817 5776 6851
rect 5724 6808 5776 6817
rect 4988 6740 5040 6792
rect 5540 6740 5592 6792
rect 7748 6808 7800 6860
rect 13268 6876 13320 6928
rect 13820 6851 13872 6860
rect 13820 6817 13838 6851
rect 13838 6817 13872 6851
rect 7932 6740 7984 6792
rect 13820 6808 13872 6817
rect 17868 6808 17920 6860
rect 10876 6740 10928 6792
rect 11704 6740 11756 6792
rect 9864 6672 9916 6724
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 13084 6604 13136 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 112 6400 164 6452
rect 1400 6400 1452 6452
rect 6000 6443 6052 6452
rect 6000 6409 6009 6443
rect 6009 6409 6043 6443
rect 6043 6409 6052 6443
rect 6000 6400 6052 6409
rect 7932 6400 7984 6452
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 11336 6443 11388 6452
rect 11336 6409 11345 6443
rect 11345 6409 11379 6443
rect 11379 6409 11388 6443
rect 11336 6400 11388 6409
rect 11704 6443 11756 6452
rect 11704 6409 11713 6443
rect 11713 6409 11747 6443
rect 11747 6409 11756 6443
rect 11704 6400 11756 6409
rect 13176 6400 13228 6452
rect 13820 6443 13872 6452
rect 13820 6409 13829 6443
rect 13829 6409 13863 6443
rect 13863 6409 13872 6443
rect 13820 6400 13872 6409
rect 5356 6332 5408 6384
rect 14648 6332 14700 6384
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 8668 6264 8720 6316
rect 8760 6196 8812 6248
rect 10508 6264 10560 6316
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 13084 6239 13136 6248
rect 13084 6205 13093 6239
rect 13093 6205 13127 6239
rect 13127 6205 13136 6239
rect 13084 6196 13136 6205
rect 8392 6128 8444 6180
rect 5540 6060 5592 6112
rect 10508 6171 10560 6180
rect 10508 6137 10517 6171
rect 10517 6137 10551 6171
rect 10551 6137 10560 6171
rect 10508 6128 10560 6137
rect 11520 6128 11572 6180
rect 10968 6060 11020 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 8668 5856 8720 5908
rect 10048 5899 10100 5908
rect 10048 5865 10057 5899
rect 10057 5865 10091 5899
rect 10091 5865 10100 5899
rect 10048 5856 10100 5865
rect 10968 5856 11020 5908
rect 13084 5856 13136 5908
rect 10692 5788 10744 5840
rect 10876 5831 10928 5840
rect 10876 5797 10885 5831
rect 10885 5797 10919 5831
rect 10919 5797 10928 5831
rect 10876 5788 10928 5797
rect 8484 5763 8536 5772
rect 8484 5729 8493 5763
rect 8493 5729 8527 5763
rect 8527 5729 8536 5763
rect 8484 5720 8536 5729
rect 11796 5720 11848 5772
rect 12716 5763 12768 5772
rect 12716 5729 12760 5763
rect 12760 5729 12768 5763
rect 12716 5720 12768 5729
rect 9496 5652 9548 5704
rect 7932 5584 7984 5636
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 8484 5312 8536 5364
rect 9496 5355 9548 5364
rect 9496 5321 9505 5355
rect 9505 5321 9539 5355
rect 9539 5321 9548 5355
rect 9496 5312 9548 5321
rect 12716 5355 12768 5364
rect 12716 5321 12725 5355
rect 12725 5321 12759 5355
rect 12759 5321 12768 5355
rect 12716 5312 12768 5321
rect 7196 5244 7248 5296
rect 8668 5244 8720 5296
rect 10048 5219 10100 5228
rect 10048 5185 10057 5219
rect 10057 5185 10091 5219
rect 10091 5185 10100 5219
rect 10048 5176 10100 5185
rect 10140 5176 10192 5228
rect 8484 5083 8536 5092
rect 8484 5049 8493 5083
rect 8493 5049 8527 5083
rect 8527 5049 8536 5083
rect 8484 5040 8536 5049
rect 8760 5040 8812 5092
rect 9128 5083 9180 5092
rect 9128 5049 9137 5083
rect 9137 5049 9171 5083
rect 9171 5049 9180 5083
rect 9128 5040 9180 5049
rect 9680 4972 9732 5024
rect 10692 4972 10744 5024
rect 11060 5015 11112 5024
rect 11060 4981 11069 5015
rect 11069 4981 11103 5015
rect 11103 4981 11112 5015
rect 11060 4972 11112 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 8484 4768 8536 4820
rect 9312 4700 9364 4752
rect 9772 4700 9824 4752
rect 11060 4700 11112 4752
rect 8668 4632 8720 4684
rect 11520 4675 11572 4684
rect 11520 4641 11529 4675
rect 11529 4641 11563 4675
rect 11563 4641 11572 4675
rect 11520 4632 11572 4641
rect 8760 4564 8812 4616
rect 9956 4607 10008 4616
rect 9956 4573 9965 4607
rect 9965 4573 9999 4607
rect 9999 4573 10008 4607
rect 9956 4564 10008 4573
rect 9404 4496 9456 4548
rect 10140 4496 10192 4548
rect 9956 4428 10008 4480
rect 10876 4428 10928 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 8668 4267 8720 4276
rect 8668 4233 8677 4267
rect 8677 4233 8711 4267
rect 8711 4233 8720 4267
rect 8668 4224 8720 4233
rect 9128 4224 9180 4276
rect 9956 4224 10008 4276
rect 10140 4224 10192 4276
rect 11060 4224 11112 4276
rect 11520 4267 11572 4276
rect 11520 4233 11529 4267
rect 11529 4233 11563 4267
rect 11563 4233 11572 4267
rect 11520 4224 11572 4233
rect 9772 4131 9824 4140
rect 9772 4097 9781 4131
rect 9781 4097 9815 4131
rect 9815 4097 9824 4131
rect 9772 4088 9824 4097
rect 10692 4088 10744 4140
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 9404 4020 9456 4072
rect 8760 3884 8812 3936
rect 10140 3884 10192 3936
rect 10784 3884 10836 3936
rect 21732 3884 21784 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 9404 3723 9456 3732
rect 9404 3689 9413 3723
rect 9413 3689 9447 3723
rect 9447 3689 9456 3723
rect 9404 3680 9456 3689
rect 10784 3723 10836 3732
rect 10784 3689 10793 3723
rect 10793 3689 10827 3723
rect 10827 3689 10836 3723
rect 10784 3680 10836 3689
rect 9680 3655 9732 3664
rect 9680 3621 9689 3655
rect 9689 3621 9723 3655
rect 9723 3621 9732 3655
rect 9680 3612 9732 3621
rect 9772 3587 9824 3596
rect 9772 3553 9781 3587
rect 9781 3553 9815 3587
rect 9815 3553 9824 3587
rect 9772 3544 9824 3553
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 8760 3179 8812 3188
rect 8760 3145 8769 3179
rect 8769 3145 8803 3179
rect 8803 3145 8812 3179
rect 8760 3136 8812 3145
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 11336 3136 11388 3188
rect 8760 2932 8812 2984
rect 11336 2932 11388 2984
rect 5632 2864 5684 2916
rect 12624 2864 12676 2916
rect 9312 2796 9364 2848
rect 10968 2796 11020 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 4344 2592 4396 2644
rect 5632 2592 5684 2644
rect 10968 2635 11020 2644
rect 10968 2601 10977 2635
rect 10977 2601 11011 2635
rect 11011 2601 11020 2635
rect 10968 2592 11020 2601
rect 13452 2592 13504 2644
rect 19524 2592 19576 2644
rect 4620 2456 4672 2508
rect 13176 2456 13228 2508
rect 13820 2499 13872 2508
rect 13820 2465 13829 2499
rect 13829 2465 13863 2499
rect 13863 2465 13872 2499
rect 13820 2456 13872 2465
rect 15752 2499 15804 2508
rect 15752 2465 15761 2499
rect 15761 2465 15795 2499
rect 15795 2465 15804 2499
rect 16856 2499 16908 2508
rect 15752 2456 15804 2465
rect 16856 2465 16865 2499
rect 16865 2465 16899 2499
rect 16899 2465 16908 2499
rect 16856 2456 16908 2465
rect 19432 2388 19484 2440
rect 20076 2456 20128 2508
rect 24216 2456 24268 2508
rect 26056 2388 26108 2440
rect 15476 2320 15528 2372
rect 16764 2320 16816 2372
rect 24860 2320 24912 2372
rect 6000 2252 6052 2304
rect 10784 2252 10836 2304
rect 13176 2295 13228 2304
rect 13176 2261 13185 2295
rect 13185 2261 13219 2295
rect 13219 2261 13228 2295
rect 13176 2252 13228 2261
rect 18052 2252 18104 2304
rect 18696 2252 18748 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 3056 76 3108 128
rect 3792 76 3844 128
rect 11060 76 11112 128
rect 11980 76 12032 128
rect 12532 76 12584 128
rect 13268 76 13320 128
rect 22192 76 22244 128
rect 23388 76 23440 128
rect 26240 76 26292 128
rect 27252 76 27304 128
<< metal2 >>
rect 478 27554 534 28000
rect 124 27526 534 27554
rect 18 24304 74 24313
rect 18 24239 74 24248
rect 32 22098 60 24239
rect 20 22092 72 22098
rect 20 22034 72 22040
rect 18 19816 74 19825
rect 18 19751 74 19760
rect 32 19718 60 19751
rect 20 19712 72 19718
rect 20 19654 72 19660
rect 124 13814 152 27526
rect 478 27520 534 27526
rect 1398 27554 1454 28000
rect 2410 27554 2466 28000
rect 3422 27554 3478 28000
rect 1398 27526 1808 27554
rect 1398 27520 1454 27526
rect 1122 26752 1178 26761
rect 1122 26687 1178 26696
rect 1136 23662 1164 26687
rect 1214 25256 1270 25265
rect 1214 25191 1270 25200
rect 1228 24274 1256 25191
rect 1216 24268 1268 24274
rect 1216 24210 1268 24216
rect 1228 23866 1256 24210
rect 1216 23860 1268 23866
rect 1216 23802 1268 23808
rect 1124 23656 1176 23662
rect 1124 23598 1176 23604
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1780 23474 1808 27526
rect 2410 27526 2728 27554
rect 2410 27520 2466 27526
rect 2700 23662 2728 27526
rect 3422 27526 3740 27554
rect 3422 27520 3478 27526
rect 3712 23662 3740 27526
rect 4434 27520 4490 28000
rect 5446 27554 5502 28000
rect 5368 27526 5502 27554
rect 4448 23662 4476 27520
rect 5368 24274 5396 27526
rect 5446 27520 5502 27526
rect 6458 27520 6514 28000
rect 7470 27520 7526 28000
rect 8390 27520 8446 28000
rect 9402 27554 9458 28000
rect 10414 27554 10470 28000
rect 11426 27554 11482 28000
rect 9048 27526 9458 27554
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6472 24410 6500 27520
rect 5448 24404 5500 24410
rect 5448 24346 5500 24352
rect 6460 24404 6512 24410
rect 6460 24346 6512 24352
rect 5356 24268 5408 24274
rect 5356 24210 5408 24216
rect 2688 23656 2740 23662
rect 2688 23598 2740 23604
rect 3700 23656 3752 23662
rect 3700 23598 3752 23604
rect 4436 23656 4488 23662
rect 4436 23598 4488 23604
rect 3424 23520 3476 23526
rect 1582 22264 1638 22273
rect 1582 22199 1638 22208
rect 1596 21146 1624 22199
rect 1584 21140 1636 21146
rect 1584 21082 1636 21088
rect 1688 20346 1716 23462
rect 1780 23446 1900 23474
rect 3424 23462 3476 23468
rect 3700 23520 3752 23526
rect 3700 23462 3752 23468
rect 1768 21004 1820 21010
rect 1768 20946 1820 20952
rect 1596 20318 1716 20346
rect 1308 18828 1360 18834
rect 1308 18770 1360 18776
rect 1320 18290 1348 18770
rect 1308 18284 1360 18290
rect 1308 18226 1360 18232
rect 1320 16017 1348 18226
rect 1596 17241 1624 20318
rect 1780 20262 1808 20946
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1688 17882 1716 18566
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1582 17232 1638 17241
rect 1582 17167 1638 17176
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 16697 1624 16934
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1688 16114 1716 17818
rect 1780 17814 1808 20198
rect 1872 19258 1900 23446
rect 3436 22778 3464 23462
rect 3424 22772 3476 22778
rect 3424 22714 3476 22720
rect 2044 22092 2096 22098
rect 2044 22034 2096 22040
rect 2056 21690 2084 22034
rect 2596 21888 2648 21894
rect 2596 21830 2648 21836
rect 2044 21684 2096 21690
rect 2044 21626 2096 21632
rect 2608 20602 2636 21830
rect 2688 21548 2740 21554
rect 2688 21490 2740 21496
rect 2596 20596 2648 20602
rect 2596 20538 2648 20544
rect 1872 19230 2084 19258
rect 1860 18080 1912 18086
rect 1860 18022 1912 18028
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1768 16516 1820 16522
rect 1768 16458 1820 16464
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1306 16008 1362 16017
rect 1306 15943 1362 15952
rect 1780 15638 1808 16458
rect 1768 15632 1820 15638
rect 1768 15574 1820 15580
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 32 13786 152 13814
rect 32 12850 60 13786
rect 1214 13696 1270 13705
rect 1214 13631 1270 13640
rect 20 12844 72 12850
rect 20 12786 72 12792
rect 1228 11694 1256 13631
rect 1412 13326 1440 14758
rect 1872 13938 1900 18022
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1964 16454 1992 16594
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 15978 1992 16390
rect 1952 15972 2004 15978
rect 1952 15914 2004 15920
rect 1964 15638 1992 15914
rect 1952 15632 2004 15638
rect 1952 15574 2004 15580
rect 1964 15366 1992 15574
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1964 14822 1992 15302
rect 2056 15162 2084 19230
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14618 1992 14758
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1964 13802 1992 14010
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1952 13796 2004 13802
rect 1952 13738 2004 13744
rect 1688 13462 1716 13738
rect 1676 13456 1728 13462
rect 1676 13398 1728 13404
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1492 13252 1544 13258
rect 1492 13194 1544 13200
rect 1504 12782 1532 13194
rect 1688 12986 1716 13398
rect 2148 13025 2176 18022
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2424 16998 2452 17682
rect 2516 17610 2544 18158
rect 2504 17604 2556 17610
rect 2504 17546 2556 17552
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2424 16590 2452 16934
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2240 14074 2268 16526
rect 2412 15972 2464 15978
rect 2412 15914 2464 15920
rect 2424 15502 2452 15914
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2320 15428 2372 15434
rect 2320 15370 2372 15376
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2226 13968 2282 13977
rect 2226 13903 2282 13912
rect 2240 13462 2268 13903
rect 2332 13802 2360 15370
rect 2424 13977 2452 15438
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 14550 2636 14758
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2410 13968 2466 13977
rect 2410 13903 2466 13912
rect 2320 13796 2372 13802
rect 2320 13738 2372 13744
rect 2608 13734 2636 14486
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2134 13016 2190 13025
rect 1676 12980 1728 12986
rect 2134 12951 2190 12960
rect 1676 12922 1728 12928
rect 2228 12912 2280 12918
rect 2228 12854 2280 12860
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1216 11688 1268 11694
rect 1216 11630 1268 11636
rect 1412 11354 1440 12242
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10130 1348 10610
rect 1504 10606 1532 12718
rect 1872 12442 1900 12718
rect 2136 12708 2188 12714
rect 2136 12650 2188 12656
rect 1860 12436 1912 12442
rect 1780 12396 1860 12424
rect 1780 11218 1808 12396
rect 1860 12378 1912 12384
rect 2148 11830 2176 12650
rect 2240 12102 2268 12854
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2136 11824 2188 11830
rect 2136 11766 2188 11772
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1688 10606 1716 10950
rect 1780 10810 1808 11154
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1504 10266 1532 10542
rect 1492 10260 1544 10266
rect 1412 10220 1492 10248
rect 1308 10124 1360 10130
rect 1308 10066 1360 10072
rect 1320 9586 1348 10066
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 848 8288 900 8294
rect 848 8230 900 8236
rect 110 6624 166 6633
rect 110 6559 166 6568
rect 124 6458 152 6559
rect 112 6452 164 6458
rect 112 6394 164 6400
rect 570 82 626 480
rect 860 82 888 8230
rect 1320 5681 1348 9522
rect 1412 9518 1440 10220
rect 1492 10202 1544 10208
rect 1872 9586 1900 11290
rect 2240 10198 2268 12038
rect 2608 11626 2636 13670
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2228 10192 2280 10198
rect 2228 10134 2280 10140
rect 2424 9722 2452 10746
rect 2700 10169 2728 21490
rect 2778 20768 2834 20777
rect 2778 20703 2834 20712
rect 2792 16658 2820 20703
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 2976 19922 3004 20198
rect 3160 19990 3188 20198
rect 3148 19984 3200 19990
rect 3148 19926 3200 19932
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 2976 19174 3004 19858
rect 3240 19236 3292 19242
rect 3240 19178 3292 19184
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 3252 18902 3280 19178
rect 3240 18896 3292 18902
rect 3240 18838 3292 18844
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 3068 18193 3096 18770
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3528 18222 3556 18566
rect 3516 18216 3568 18222
rect 3054 18184 3110 18193
rect 3516 18158 3568 18164
rect 3054 18119 3110 18128
rect 3068 18086 3096 18119
rect 3056 18080 3108 18086
rect 3056 18022 3108 18028
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2884 16726 2912 17478
rect 3068 17338 3096 18022
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3160 16794 3188 17478
rect 3344 17338 3372 17682
rect 3436 17542 3464 18022
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3436 17066 3464 17478
rect 3424 17060 3476 17066
rect 3424 17002 3476 17008
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 2780 16652 2832 16658
rect 2780 16594 2832 16600
rect 2792 16250 2820 16594
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 3160 15706 3188 16730
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 3160 15026 3188 15370
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3068 13530 3096 13874
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2884 12442 2912 12582
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2792 10266 2820 11630
rect 2884 11354 2912 12242
rect 3068 11762 3096 12650
rect 3056 11756 3108 11762
rect 3056 11698 3108 11704
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2686 10160 2742 10169
rect 2686 10095 2742 10104
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 2424 9518 2452 9658
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 1412 9110 1440 9454
rect 2042 9344 2098 9353
rect 2042 9279 2098 9288
rect 1400 9104 1452 9110
rect 1400 9046 1452 9052
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 1504 8294 1532 8978
rect 1492 8288 1544 8294
rect 1492 8230 1544 8236
rect 1858 7576 1914 7585
rect 1858 7511 1914 7520
rect 1872 7342 1900 7511
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1412 6458 1440 6802
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1306 5672 1362 5681
rect 1306 5607 1362 5616
rect 570 54 888 82
rect 1766 82 1822 480
rect 2056 82 2084 9279
rect 2884 9178 2912 10066
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2976 8498 3004 8978
rect 3068 8634 3096 11698
rect 3160 10266 3188 14282
rect 3344 13190 3372 16390
rect 3436 14890 3464 17002
rect 3528 15706 3556 17546
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3620 14958 3648 16934
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 3424 14884 3476 14890
rect 3424 14826 3476 14832
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14618 3648 14758
rect 3608 14612 3660 14618
rect 3528 14572 3608 14600
rect 3528 13802 3556 14572
rect 3608 14554 3660 14560
rect 3712 13814 3740 23462
rect 4988 23180 5040 23186
rect 4988 23122 5040 23128
rect 5000 22438 5028 23122
rect 4988 22432 5040 22438
rect 4988 22374 5040 22380
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 4356 21554 4384 21830
rect 4344 21548 4396 21554
rect 4344 21490 4396 21496
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 3792 20936 3844 20942
rect 3792 20878 3844 20884
rect 3804 20058 3832 20878
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3896 18970 3924 19790
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 3988 18834 4016 21286
rect 4252 21072 4304 21078
rect 4252 21014 4304 21020
rect 4264 20602 4292 21014
rect 4252 20596 4304 20602
rect 4252 20538 4304 20544
rect 4264 20262 4292 20538
rect 4356 20534 4384 21490
rect 5000 21418 5028 22374
rect 5356 22092 5408 22098
rect 5356 22034 5408 22040
rect 5368 21622 5396 22034
rect 5356 21616 5408 21622
rect 5356 21558 5408 21564
rect 4988 21412 5040 21418
rect 4988 21354 5040 21360
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 4344 20528 4396 20534
rect 4344 20470 4396 20476
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4068 19984 4120 19990
rect 4068 19926 4120 19932
rect 4080 18902 4108 19926
rect 4356 19378 4384 20470
rect 4448 20466 4476 20878
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4816 20466 4844 20742
rect 4436 20460 4488 20466
rect 4436 20402 4488 20408
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4448 19854 4476 20402
rect 4816 20369 4844 20402
rect 4802 20360 4858 20369
rect 4802 20295 4858 20304
rect 5000 19990 5028 21354
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 4988 19984 5040 19990
rect 4988 19926 5040 19932
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4988 19712 5040 19718
rect 5092 19700 5120 21286
rect 5040 19672 5120 19700
rect 4988 19654 5040 19660
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4344 19168 4396 19174
rect 4344 19110 4396 19116
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4068 18896 4120 18902
rect 4068 18838 4120 18844
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 4356 18426 4384 19110
rect 4540 18902 4568 19110
rect 4528 18896 4580 18902
rect 4528 18838 4580 18844
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4436 18692 4488 18698
rect 4436 18634 4488 18640
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3792 15972 3844 15978
rect 3792 15914 3844 15920
rect 3804 14346 3832 15914
rect 3896 15910 3924 18158
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4080 17134 4108 17478
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4080 16794 4108 17070
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4080 16182 4108 16594
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4080 16046 4108 16118
rect 4068 16040 4120 16046
rect 3988 16000 4068 16028
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3988 15638 4016 16000
rect 4068 15982 4120 15988
rect 3976 15632 4028 15638
rect 4160 15632 4212 15638
rect 3976 15574 4028 15580
rect 4080 15580 4160 15586
rect 4080 15574 4212 15580
rect 4344 15632 4396 15638
rect 4344 15574 4396 15580
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3792 14340 3844 14346
rect 3792 14282 3844 14288
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 3516 13796 3568 13802
rect 3516 13738 3568 13744
rect 3620 13786 3740 13814
rect 3424 13728 3476 13734
rect 3424 13670 3476 13676
rect 3436 13530 3464 13670
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3528 13394 3556 13738
rect 3620 13569 3648 13786
rect 3606 13560 3662 13569
rect 3606 13495 3662 13504
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3344 9178 3372 13126
rect 3528 12442 3556 13330
rect 3804 12442 3832 14010
rect 3896 13802 3924 15302
rect 3988 14074 4016 15574
rect 4080 15558 4200 15574
rect 4080 14822 4108 15558
rect 4356 15502 4384 15574
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 3884 13796 3936 13802
rect 3884 13738 3936 13744
rect 3896 13297 3924 13738
rect 3882 13288 3938 13297
rect 3882 13223 3938 13232
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3436 10538 3464 11154
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3436 10266 3464 10474
rect 3528 10470 3556 11562
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 11286 3648 11494
rect 3608 11280 3660 11286
rect 3608 11222 3660 11228
rect 3620 10520 3648 11222
rect 3700 11076 3752 11082
rect 3700 11018 3752 11024
rect 3712 10674 3740 11018
rect 3896 10674 3924 12650
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3988 10554 4016 13806
rect 4080 13462 4108 14758
rect 4172 14482 4200 14894
rect 4264 14618 4292 15370
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4252 14340 4304 14346
rect 4252 14282 4304 14288
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 4264 12850 4292 14282
rect 4448 13814 4476 18634
rect 4816 18086 4844 18770
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4816 17338 4844 18022
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 4632 15502 4660 17274
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4724 16046 4752 16594
rect 4908 16046 4936 16594
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4632 14958 4660 15438
rect 4816 15026 4844 15506
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4540 14550 4568 14758
rect 4528 14544 4580 14550
rect 4528 14486 4580 14492
rect 4632 14482 4660 14894
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4632 14074 4660 14418
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4816 13814 4844 14962
rect 5000 13814 5028 19654
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5276 18358 5304 18566
rect 5264 18352 5316 18358
rect 5264 18294 5316 18300
rect 5276 18154 5304 18294
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 5092 14346 5120 18022
rect 5276 17882 5304 18090
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5184 17066 5212 17682
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5368 14890 5396 16526
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 5080 14000 5132 14006
rect 5460 13977 5488 24346
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 7012 23656 7064 23662
rect 7012 23598 7064 23604
rect 7024 23322 7052 23598
rect 7104 23520 7156 23526
rect 7104 23462 7156 23468
rect 7116 23322 7144 23462
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 6368 23248 6420 23254
rect 6368 23190 6420 23196
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 6288 22778 6316 23054
rect 6380 22778 6408 23190
rect 6276 22772 6328 22778
rect 6276 22714 6328 22720
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 6012 22030 6040 22374
rect 6380 22166 6408 22714
rect 7116 22642 7144 23258
rect 7196 23112 7248 23118
rect 7196 23054 7248 23060
rect 7208 22642 7236 23054
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 7012 22500 7064 22506
rect 7012 22442 7064 22448
rect 7024 22234 7052 22442
rect 7012 22228 7064 22234
rect 7012 22170 7064 22176
rect 6368 22160 6420 22166
rect 6368 22102 6420 22108
rect 6920 22160 6972 22166
rect 6920 22102 6972 22108
rect 6184 22092 6236 22098
rect 6184 22034 6236 22040
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 5540 21956 5592 21962
rect 5540 21898 5592 21904
rect 5552 18222 5580 21898
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6012 21690 6040 21966
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 6104 21554 6132 21830
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 6196 21350 6224 22034
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6644 21412 6696 21418
rect 6644 21354 6696 21360
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6656 21078 6684 21354
rect 6092 21072 6144 21078
rect 6092 21014 6144 21020
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 6000 20936 6052 20942
rect 6000 20878 6052 20884
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 6012 20058 6040 20878
rect 6104 20602 6132 21014
rect 6184 20868 6236 20874
rect 6184 20810 6236 20816
rect 6092 20596 6144 20602
rect 6092 20538 6144 20544
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 6196 19922 6224 20810
rect 6748 20466 6776 21830
rect 6932 21146 6960 22102
rect 7024 21690 7052 22170
rect 7012 21684 7064 21690
rect 7012 21626 7064 21632
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 6932 20602 6960 21082
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6380 19922 6408 20198
rect 6748 19990 6776 20402
rect 6932 20312 6960 20538
rect 7012 20324 7064 20330
rect 6932 20284 7012 20312
rect 7012 20266 7064 20272
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6196 19514 6224 19858
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 6380 19310 6408 19858
rect 6368 19304 6420 19310
rect 6368 19246 6420 19252
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 7012 19236 7064 19242
rect 7012 19178 7064 19184
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6656 18426 6684 18702
rect 6644 18420 6696 18426
rect 6564 18380 6644 18408
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5552 17678 5580 18022
rect 6472 17882 6500 18294
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5552 17338 5580 17614
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 6012 17270 6040 17750
rect 6000 17264 6052 17270
rect 6000 17206 6052 17212
rect 6564 17202 6592 18380
rect 6644 18362 6696 18368
rect 6748 18154 6776 19110
rect 6736 18148 6788 18154
rect 6736 18090 6788 18096
rect 6932 17882 6960 19178
rect 7024 18902 7052 19178
rect 7012 18896 7064 18902
rect 7012 18838 7064 18844
rect 7208 18698 7236 22578
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7300 18834 7328 21966
rect 7484 20505 7512 27520
rect 8404 27492 8524 27520
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 7932 23520 7984 23526
rect 7932 23462 7984 23468
rect 7748 21412 7800 21418
rect 7748 21354 7800 21360
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7470 20496 7526 20505
rect 7668 20466 7696 20878
rect 7470 20431 7526 20440
rect 7656 20460 7708 20466
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7392 19378 7420 19790
rect 7484 19446 7512 20431
rect 7656 20402 7708 20408
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7668 19378 7696 20402
rect 7760 19922 7788 21354
rect 7944 21078 7972 23462
rect 8024 21684 8076 21690
rect 8024 21626 8076 21632
rect 8036 21350 8064 21626
rect 8024 21344 8076 21350
rect 8024 21286 8076 21292
rect 8036 21078 8064 21286
rect 7932 21072 7984 21078
rect 7932 21014 7984 21020
rect 8024 21072 8076 21078
rect 8024 21014 8076 21020
rect 8036 20058 8064 21014
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7392 18970 7420 19314
rect 7760 19174 7788 19858
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7288 18828 7340 18834
rect 7288 18770 7340 18776
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 7300 18290 7328 18770
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7484 18222 7512 18566
rect 7576 18426 7604 18838
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 7286 17912 7342 17921
rect 6920 17876 6972 17882
rect 7286 17847 7342 17856
rect 6920 17818 6972 17824
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6656 17338 6684 17614
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6276 17128 6328 17134
rect 6276 17070 6328 17076
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 6012 15366 6040 15982
rect 6288 15570 6316 17070
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6276 15564 6328 15570
rect 6196 15524 6276 15552
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6012 14958 6040 15302
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 6000 14952 6052 14958
rect 6052 14912 6132 14940
rect 6000 14894 6052 14900
rect 5552 14482 5580 14894
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 5080 13942 5132 13948
rect 5446 13968 5502 13977
rect 4356 13786 4476 13814
rect 4724 13786 4844 13814
rect 4908 13786 5028 13814
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4172 11694 4200 12378
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4264 10810 4292 12582
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 3700 10532 3752 10538
rect 3620 10492 3700 10520
rect 3700 10474 3752 10480
rect 3804 10526 4016 10554
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3712 9178 3740 9454
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3700 9172 3752 9178
rect 3700 9114 3752 9120
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 1766 54 2084 82
rect 3054 128 3110 480
rect 3804 134 3832 10526
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 3988 9518 4016 9930
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 4080 9178 4108 10066
rect 4160 9988 4212 9994
rect 4160 9930 4212 9936
rect 4172 9217 4200 9930
rect 4158 9208 4214 9217
rect 4068 9172 4120 9178
rect 4158 9143 4214 9152
rect 4068 9114 4120 9120
rect 4172 9083 4200 9143
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 7002 4016 8230
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 4356 2650 4384 13786
rect 4724 13326 4752 13786
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4436 12844 4488 12850
rect 4436 12786 4488 12792
rect 4448 10452 4476 12786
rect 4540 12782 4568 13194
rect 4908 12782 4936 13786
rect 5092 13462 5120 13942
rect 5446 13903 5502 13912
rect 5552 13870 5580 14418
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6012 14006 6040 14418
rect 6104 14278 6132 14912
rect 6196 14618 6224 15524
rect 6276 15506 6328 15512
rect 6276 15428 6328 15434
rect 6276 15370 6328 15376
rect 6288 14822 6316 15370
rect 6276 14816 6328 14822
rect 6276 14758 6328 14764
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6288 14414 6316 14758
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 5540 13864 5592 13870
rect 6104 13814 6132 14214
rect 6288 14074 6316 14350
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 6288 13870 6316 14010
rect 5540 13806 5592 13812
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 5092 13190 5120 13398
rect 5552 13394 5580 13806
rect 6012 13786 6132 13814
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4804 12300 4856 12306
rect 4856 12260 4936 12288
rect 4804 12242 4856 12248
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4632 11286 4660 12106
rect 4724 11694 4752 12106
rect 4908 11898 4936 12260
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4908 11694 4936 11834
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4908 11354 4936 11630
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 4712 11144 4764 11150
rect 4710 11112 4712 11121
rect 4764 11112 4766 11121
rect 4710 11047 4766 11056
rect 4724 10742 4752 11047
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4620 10464 4672 10470
rect 4448 10424 4620 10452
rect 4448 10266 4476 10424
rect 4620 10406 4672 10412
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 5000 10198 5028 12582
rect 6012 12442 6040 13786
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 13258 6224 13670
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6184 13252 6236 13258
rect 6184 13194 6236 13200
rect 6196 12646 6224 13194
rect 6380 12986 6408 13330
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6472 12918 6500 13330
rect 6460 12912 6512 12918
rect 6460 12854 6512 12860
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 5092 11558 5120 12242
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5460 11694 5488 12174
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11694 6040 12038
rect 6196 11898 6224 12582
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 5092 10130 5120 11494
rect 5184 11354 5212 11494
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5184 11218 5212 11290
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5368 10538 5396 10950
rect 5460 10810 5488 11290
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5276 10198 5304 10474
rect 5368 10266 5396 10474
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9518 5028 9998
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4540 9042 4568 9318
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4540 8294 4568 8978
rect 5000 8294 5028 9454
rect 5092 9382 5120 10066
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5276 9518 5304 9930
rect 5552 9926 5580 11630
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6104 11150 6132 11562
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6012 10606 6040 10950
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6104 10266 6132 11086
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5080 9376 5132 9382
rect 5080 9318 5132 9324
rect 5276 8838 5304 9454
rect 5552 9450 5580 9862
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5552 9110 5580 9386
rect 6012 9110 6040 9454
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4540 7954 4568 8230
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4540 7206 4568 7890
rect 5000 7886 5028 8230
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5000 7206 5028 7822
rect 5092 7342 5120 8774
rect 5552 8498 5580 9046
rect 6012 8838 6040 9046
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6012 8498 6040 8774
rect 6104 8634 6132 8978
rect 6196 8906 6224 9318
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6196 8498 6224 8842
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4540 1329 4568 7142
rect 5000 6798 5028 7142
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 5092 6662 5120 7278
rect 5368 6866 5396 8434
rect 6196 8090 6224 8434
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5460 7546 5488 7890
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5448 7268 5500 7274
rect 5552 7256 5580 7754
rect 6472 7750 6500 12038
rect 6564 10577 6592 16186
rect 6644 15496 6696 15502
rect 6748 15484 6776 17478
rect 6932 17338 6960 17818
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6696 15456 6776 15484
rect 6644 15438 6696 15444
rect 6656 14278 6684 15438
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6656 11286 6684 14214
rect 6840 13802 6868 14418
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 6932 13682 6960 17070
rect 7300 16153 7328 17847
rect 7392 17338 7420 18090
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7392 16658 7420 17274
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7392 16182 7420 16594
rect 7484 16590 7512 18158
rect 7760 18086 7788 19110
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7760 17882 7788 18022
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7760 16998 7788 17818
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7944 17134 7972 17478
rect 7932 17128 7984 17134
rect 8116 17128 8168 17134
rect 7932 17070 7984 17076
rect 8036 17088 8116 17116
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7380 16176 7432 16182
rect 7286 16144 7342 16153
rect 7380 16118 7432 16124
rect 7286 16079 7342 16088
rect 7300 16046 7328 16079
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7760 15978 7788 16458
rect 7944 16046 7972 17070
rect 8036 16794 8064 17088
rect 8116 17070 8168 17076
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8036 16454 8064 16730
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7012 14816 7064 14822
rect 7576 14804 7604 15846
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7668 14958 7696 15506
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7576 14776 7696 14804
rect 7012 14758 7064 14764
rect 6840 13654 6960 13682
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6550 10568 6606 10577
rect 6550 10503 6606 10512
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9654 6776 9862
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6656 8430 6684 9114
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6656 7954 6684 8366
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6748 7342 6776 9386
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 5724 7268 5776 7274
rect 5552 7228 5724 7256
rect 5448 7210 5500 7216
rect 5724 7210 5776 7216
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 5460 6934 5488 7210
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5736 6866 5764 7210
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 4185 5120 6598
rect 5368 6390 5396 6802
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5552 6118 5580 6734
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6458 6040 7210
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5078 4176 5134 4185
rect 5078 4111 5134 4120
rect 5552 2689 5580 6054
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5538 2680 5594 2689
rect 5644 2650 5672 2858
rect 5538 2615 5594 2624
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4526 1320 4582 1329
rect 4526 1255 4582 1264
rect 3054 76 3056 128
rect 3108 76 3110 128
rect 570 0 626 54
rect 1766 0 1822 54
rect 3054 0 3110 76
rect 3792 128 3844 134
rect 3792 70 3844 76
rect 4342 82 4398 480
rect 4632 82 4660 2450
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 4342 54 4660 82
rect 5630 82 5686 480
rect 6012 82 6040 2246
rect 5630 54 6040 82
rect 6840 82 6868 13654
rect 7024 13394 7052 14758
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13870 7512 14214
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7576 13530 7604 13874
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 11150 6960 12582
rect 7012 11280 7064 11286
rect 7012 11222 7064 11228
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6932 10810 6960 11086
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7024 10674 7052 11222
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 7546 7052 10406
rect 7116 10266 7144 10542
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7116 9178 7144 10066
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7208 5302 7236 12718
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7392 11762 7420 12310
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7392 11558 7420 11698
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7484 10169 7512 13262
rect 7668 12306 7696 14776
rect 7760 13530 7788 15914
rect 7944 15638 7972 15982
rect 8036 15910 8064 16390
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 7932 15632 7984 15638
rect 7984 15580 8064 15586
rect 7932 15574 8064 15580
rect 7944 15558 8064 15574
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7944 14958 7972 15438
rect 7932 14952 7984 14958
rect 7852 14912 7932 14940
rect 7852 13870 7880 14912
rect 7932 14894 7984 14900
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7944 13734 7972 14350
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12714 7788 13126
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7668 11830 7696 12242
rect 7656 11824 7708 11830
rect 7562 11792 7618 11801
rect 7656 11766 7708 11772
rect 7562 11727 7618 11736
rect 7576 11286 7604 11727
rect 7668 11354 7696 11766
rect 7760 11626 7788 12650
rect 7852 11830 7880 13670
rect 7944 13394 7972 13670
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7944 12646 7972 13330
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7944 11898 7972 12582
rect 8036 12238 8064 15558
rect 8220 13814 8248 19382
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8312 14278 8340 14894
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8312 13870 8340 14214
rect 8128 13786 8248 13814
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7760 11286 7788 11562
rect 7564 11280 7616 11286
rect 7564 11222 7616 11228
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7576 10742 7604 11222
rect 8128 11218 8156 13786
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8220 12102 8248 12718
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11694 8248 12038
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8220 10810 8248 11630
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 7564 10736 7616 10742
rect 7564 10678 7616 10684
rect 7656 10736 7708 10742
rect 7656 10678 7708 10684
rect 7470 10160 7526 10169
rect 7470 10095 7526 10104
rect 7668 9926 7696 10678
rect 8312 10198 8340 13466
rect 8404 10198 8432 24006
rect 8496 23186 8524 27492
rect 8944 24268 8996 24274
rect 8944 24210 8996 24216
rect 8956 23866 8984 24210
rect 8944 23860 8996 23866
rect 8944 23802 8996 23808
rect 9048 23798 9076 27526
rect 9402 27520 9458 27526
rect 10152 27526 10470 27554
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9232 24410 9260 24550
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9036 23792 9088 23798
rect 9036 23734 9088 23740
rect 9324 23474 9352 24550
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9402 23760 9458 23769
rect 9402 23695 9458 23704
rect 9416 23662 9444 23695
rect 9692 23662 9720 24346
rect 10152 23866 10180 27526
rect 10414 27520 10470 27526
rect 11072 27526 11482 27554
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10784 25152 10836 25158
rect 10784 25094 10836 25100
rect 10796 24954 10824 25094
rect 11072 24954 11100 27526
rect 11426 27520 11482 27526
rect 12438 27520 12494 28000
rect 13450 27532 13506 28000
rect 13450 27520 13452 27532
rect 11428 25356 11480 25362
rect 11428 25298 11480 25304
rect 11336 25288 11388 25294
rect 11336 25230 11388 25236
rect 10784 24948 10836 24954
rect 10784 24890 10836 24896
rect 11060 24948 11112 24954
rect 11060 24890 11112 24896
rect 10796 24750 10824 24890
rect 10784 24744 10836 24750
rect 10784 24686 10836 24692
rect 11244 24676 11296 24682
rect 11244 24618 11296 24624
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 10336 23866 10364 24210
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10888 23730 10916 24142
rect 10876 23724 10928 23730
rect 10876 23666 10928 23672
rect 9404 23656 9456 23662
rect 9404 23598 9456 23604
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 9232 23446 9352 23474
rect 8484 23180 8536 23186
rect 8484 23122 8536 23128
rect 8496 22778 8524 23122
rect 8484 22772 8536 22778
rect 8484 22714 8536 22720
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8680 21962 8708 22510
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 8668 21956 8720 21962
rect 8668 21898 8720 21904
rect 8956 21554 8984 21966
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8484 21412 8536 21418
rect 8484 21354 8536 21360
rect 8496 20262 8524 21354
rect 8864 21146 8892 21490
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8680 18970 8708 19314
rect 8772 19242 8800 19654
rect 8864 19378 8892 20334
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8760 19236 8812 19242
rect 8760 19178 8812 19184
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 9232 18358 9260 23446
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 11256 23322 11284 24618
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 11348 23254 11376 25230
rect 11440 24750 11468 25298
rect 11704 24880 11756 24886
rect 11704 24822 11756 24828
rect 11428 24744 11480 24750
rect 11428 24686 11480 24692
rect 11428 23520 11480 23526
rect 11428 23462 11480 23468
rect 11440 23254 11468 23462
rect 11336 23248 11388 23254
rect 11336 23190 11388 23196
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 9772 23180 9824 23186
rect 9772 23122 9824 23128
rect 9956 23180 10008 23186
rect 9956 23122 10008 23128
rect 9784 22710 9812 23122
rect 9772 22704 9824 22710
rect 9772 22646 9824 22652
rect 9404 22500 9456 22506
rect 9404 22442 9456 22448
rect 9416 20466 9444 22442
rect 9968 22438 9996 23122
rect 10324 22976 10376 22982
rect 10324 22918 10376 22924
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10336 22642 10364 22918
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 10796 22506 10824 22918
rect 11348 22778 11376 23190
rect 11440 22778 11468 23190
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11152 22704 11204 22710
rect 11152 22646 11204 22652
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 10968 22500 11020 22506
rect 10968 22442 11020 22448
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 9784 21690 9812 22102
rect 9772 21684 9824 21690
rect 9772 21626 9824 21632
rect 9680 21616 9732 21622
rect 9680 21558 9732 21564
rect 9692 21010 9720 21558
rect 9968 21554 9996 22374
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9692 20602 9720 20946
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9404 20460 9456 20466
rect 9404 20402 9456 20408
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9692 19990 9720 20198
rect 9680 19984 9732 19990
rect 9680 19926 9732 19932
rect 9404 19916 9456 19922
rect 9404 19858 9456 19864
rect 9416 19174 9444 19858
rect 9968 19718 9996 21490
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 10060 20806 10088 21422
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9968 19242 9996 19654
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9324 17814 9352 18226
rect 9312 17808 9364 17814
rect 9312 17750 9364 17756
rect 9036 17536 9088 17542
rect 9036 17478 9088 17484
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8588 15706 8616 16594
rect 8956 16046 8984 17070
rect 9048 16726 9076 17478
rect 9416 17202 9444 19110
rect 9600 18698 9628 19178
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9600 18290 9628 18634
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9232 16794 9260 17070
rect 9508 16794 9536 17682
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9036 16720 9088 16726
rect 9036 16662 9088 16668
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9508 16114 9536 16526
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8956 15434 8984 15982
rect 8944 15428 8996 15434
rect 8944 15370 8996 15376
rect 9140 15366 9168 15982
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9140 14958 9168 15302
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 8772 14414 8800 14894
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8772 14074 8800 14350
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8956 13870 8984 13942
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9586 7880 9862
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7288 9376 7340 9382
rect 7760 9353 7788 9386
rect 7288 9318 7340 9324
rect 7746 9344 7802 9353
rect 7300 8498 7328 9318
rect 7746 9279 7802 9288
rect 8128 9178 8156 10066
rect 8220 9722 8248 10066
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8220 9217 8248 9658
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8206 9208 8262 9217
rect 8116 9172 8168 9178
rect 8206 9143 8262 9152
rect 8116 9114 8168 9120
rect 8220 9110 8248 9143
rect 7932 9104 7984 9110
rect 7932 9046 7984 9052
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7760 6866 7788 8570
rect 7944 8090 7972 9046
rect 8312 9042 8340 9590
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8312 8634 8340 8978
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7760 6322 7788 6802
rect 7944 6798 7972 8026
rect 8128 8022 8156 8366
rect 8220 8022 8248 8502
rect 8404 8498 8432 9386
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8404 8362 8432 8434
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 6934 8156 7822
rect 8220 7546 8248 7958
rect 8404 7546 8432 8298
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7944 6458 7972 6734
rect 8404 6458 8432 7482
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7760 6225 7788 6258
rect 7746 6216 7802 6225
rect 7746 6151 7802 6160
rect 7944 5642 7972 6394
rect 8404 6186 8432 6394
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8496 5778 8524 13262
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8588 12442 8616 12582
rect 8956 12442 8984 13806
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9048 12782 9076 13262
rect 9140 13190 9168 14894
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9218 13832 9274 13841
rect 9218 13767 9274 13776
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 8588 12306 8616 12378
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8588 10810 8616 11154
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8588 8498 8616 8910
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8588 8090 8616 8434
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8680 6322 8708 12106
rect 9048 11762 9076 12718
rect 9140 12714 9168 13126
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9232 11218 9260 13767
rect 9324 13462 9352 14214
rect 9416 13938 9444 14962
rect 9600 14482 9628 18226
rect 9968 16522 9996 19178
rect 10060 19174 10088 20742
rect 10152 20330 10180 21286
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10704 21146 10732 21966
rect 10796 21690 10824 22442
rect 10980 22166 11008 22442
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10140 20324 10192 20330
rect 10140 20266 10192 20272
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10704 20058 10732 20402
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 11072 19514 11100 19926
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 11164 19446 11192 22646
rect 11440 22234 11468 22714
rect 11428 22228 11480 22234
rect 11428 22170 11480 22176
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11348 20330 11376 21082
rect 11440 20602 11468 22170
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 11428 20596 11480 20602
rect 11428 20538 11480 20544
rect 11336 20324 11388 20330
rect 11336 20266 11388 20272
rect 11532 19854 11560 22102
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 11624 21622 11652 22034
rect 11612 21616 11664 21622
rect 11612 21558 11664 21564
rect 11624 21350 11652 21558
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11624 20874 11652 21286
rect 11612 20868 11664 20874
rect 11612 20810 11664 20816
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11348 19514 11376 19790
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 11152 19440 11204 19446
rect 11152 19382 11204 19388
rect 11060 19304 11112 19310
rect 11164 19281 11192 19382
rect 11060 19246 11112 19252
rect 11150 19272 11206 19281
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 10152 18086 10180 18838
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10152 17882 10180 18022
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10152 17338 10180 17682
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10704 17202 10732 17478
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10152 16998 10180 17070
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10152 16794 10180 16934
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 10152 16182 10180 16730
rect 10140 16176 10192 16182
rect 10060 16136 10140 16164
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 9876 15638 9904 15982
rect 9864 15632 9916 15638
rect 9864 15574 9916 15580
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 14618 9720 15506
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9784 14822 9812 15370
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9680 14612 9732 14618
rect 9732 14572 9812 14600
rect 9680 14554 9732 14560
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9692 13530 9720 14010
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9784 12594 9812 14572
rect 9876 13326 9904 15574
rect 10060 15162 10088 16136
rect 10140 16118 10192 16124
rect 11072 16114 11100 19246
rect 11150 19207 11206 19216
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10152 14006 10180 15846
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10796 15570 10824 15982
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10796 15366 10824 15506
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14414 10732 14826
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10520 13870 10548 14214
rect 10704 14074 10732 14350
rect 10796 14278 10824 15302
rect 11072 15026 11100 15302
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10888 14550 10916 14758
rect 10876 14544 10928 14550
rect 10876 14486 10928 14492
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10888 14006 10916 14486
rect 10876 14000 10928 14006
rect 10796 13960 10876 13988
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 10336 12986 10364 13330
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10796 12918 10824 13960
rect 10876 13942 10928 13948
rect 11164 13841 11192 19207
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11256 16250 11284 18566
rect 11428 18216 11480 18222
rect 11428 18158 11480 18164
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11348 16794 11376 17614
rect 11440 17270 11468 18158
rect 11520 18148 11572 18154
rect 11520 18090 11572 18096
rect 11532 17814 11560 18090
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11532 17338 11560 17750
rect 11612 17604 11664 17610
rect 11612 17546 11664 17552
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11624 16590 11652 17546
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11624 15706 11652 16526
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11150 13832 11206 13841
rect 10968 13796 11020 13802
rect 11150 13767 11206 13776
rect 10968 13738 11020 13744
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10796 12646 10824 12854
rect 10888 12850 10916 13126
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10980 12753 11008 13738
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11624 12850 11652 13398
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 10966 12744 11022 12753
rect 10966 12679 11022 12688
rect 10784 12640 10836 12646
rect 9784 12566 9904 12594
rect 10784 12582 10836 12588
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9416 11694 9444 12378
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 8956 9722 8984 10950
rect 9034 10704 9090 10713
rect 9034 10639 9090 10648
rect 9048 10538 9076 10639
rect 9140 10606 9168 10950
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 9048 10266 9076 10474
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 9140 9654 9168 10542
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9692 10266 9720 10474
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9692 9586 9720 10202
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8772 7410 8800 7822
rect 8864 7546 8892 9318
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9692 8430 9720 8978
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 9784 7342 9812 12378
rect 9876 12306 9904 12566
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 9876 12170 9904 12242
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9876 11898 9904 12106
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 10060 11354 10088 12242
rect 10520 12170 10548 12242
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10428 11762 10456 12038
rect 10796 11898 10824 12582
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10796 11558 10824 11834
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10980 11354 11008 12242
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 11348 11286 11376 11494
rect 11440 11354 11468 12174
rect 11532 11558 11560 12310
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 9968 10470 9996 11154
rect 10428 10606 10456 11154
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 10060 9110 10088 9386
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 10060 8022 10088 9046
rect 10152 9042 10180 9998
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10704 8974 10732 11086
rect 11348 10810 11376 11222
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11348 10606 11376 10746
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 11348 10266 11376 10542
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 10980 9382 11008 10134
rect 11150 10024 11206 10033
rect 11150 9959 11206 9968
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10980 8838 11008 9318
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10612 8362 10640 8774
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10048 8016 10100 8022
rect 9968 7976 10048 8004
rect 9968 7478 9996 7976
rect 10048 7958 10100 7964
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8680 5914 8708 6258
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 8496 5370 8524 5714
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8496 4826 8524 5034
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8680 4690 8708 5238
rect 8772 5098 8800 6190
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8680 4282 8708 4626
rect 8772 4622 8800 5034
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 9140 4282 9168 5034
rect 9324 4758 9352 7142
rect 9784 7002 9812 7278
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9876 6730 9904 7210
rect 10060 6934 10088 7822
rect 10152 7002 10180 8298
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10336 7274 10364 7482
rect 10888 7410 10916 8434
rect 10980 8362 11008 8774
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10324 7268 10376 7274
rect 10324 7210 10376 7216
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 10888 6798 10916 7346
rect 10980 6934 11008 7686
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10520 6186 10548 6258
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9508 5370 9536 5646
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 10060 5234 10088 5850
rect 10888 5846 10916 6258
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10980 5914 11008 6054
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9312 4752 9364 4758
rect 9312 4694 9364 4700
rect 9404 4548 9456 4554
rect 9404 4490 9456 4496
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 8680 3369 8708 4218
rect 9416 4078 9444 4490
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8666 3360 8722 3369
rect 8666 3295 8722 3304
rect 8772 3194 8800 3878
rect 9416 3738 9444 4014
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9692 3670 9720 4966
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9784 4146 9812 4694
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9968 4486 9996 4558
rect 10152 4554 10180 5170
rect 10704 5030 10732 5782
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 11072 4758 11100 4966
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 9968 4282 9996 4422
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9784 3602 9812 4082
rect 10152 3942 10180 4218
rect 10888 4146 10916 4422
rect 11072 4282 11100 4694
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11164 4154 11192 9959
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11256 8090 11284 8978
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11348 6458 11376 6870
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11440 4154 11468 11018
rect 11532 10674 11560 11494
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11532 8498 11560 9046
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11716 6882 11744 24822
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 12072 24608 12124 24614
rect 12072 24550 12124 24556
rect 11980 23860 12032 23866
rect 11980 23802 12032 23808
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11808 20942 11836 23054
rect 11992 22574 12020 23802
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 11900 21010 11928 22170
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11900 20602 11928 20946
rect 11888 20596 11940 20602
rect 11992 20584 12020 22510
rect 12084 22098 12112 24550
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 12176 21146 12204 23462
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 12268 21962 12296 22034
rect 12256 21956 12308 21962
rect 12256 21898 12308 21904
rect 12268 21554 12296 21898
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 11992 20556 12112 20584
rect 11888 20538 11940 20544
rect 11796 18896 11848 18902
rect 11796 18838 11848 18844
rect 11808 18086 11836 18838
rect 11888 18352 11940 18358
rect 11888 18294 11940 18300
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11808 16726 11836 18022
rect 11900 17678 11928 18294
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11796 16720 11848 16726
rect 11796 16662 11848 16668
rect 11808 16250 11836 16662
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11808 14618 11836 15438
rect 11992 15162 12020 15574
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11808 14385 11836 14418
rect 11794 14376 11850 14385
rect 11794 14311 11850 14320
rect 12084 13814 12112 20556
rect 12176 19990 12204 21082
rect 12164 19984 12216 19990
rect 12164 19926 12216 19932
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 12268 17066 12296 18022
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12360 15502 12388 24686
rect 12452 24410 12480 27520
rect 13504 27520 13506 27532
rect 14462 27520 14518 28000
rect 14740 27532 14792 27538
rect 13452 27474 13504 27480
rect 13464 27443 13492 27474
rect 13544 25356 13596 25362
rect 13544 25298 13596 25304
rect 12992 25220 13044 25226
rect 12992 25162 13044 25168
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12636 24342 12664 25094
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12624 24336 12676 24342
rect 12624 24278 12676 24284
rect 12532 24132 12584 24138
rect 12532 24074 12584 24080
rect 12544 23730 12572 24074
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12532 23588 12584 23594
rect 12636 23576 12664 24278
rect 12584 23548 12664 23576
rect 12532 23530 12584 23536
rect 12622 23488 12678 23497
rect 12622 23423 12678 23432
rect 12636 22778 12664 23423
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12728 19922 12756 24550
rect 12808 24336 12860 24342
rect 12808 24278 12860 24284
rect 12820 22982 12848 24278
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 12912 23798 12940 24142
rect 12900 23792 12952 23798
rect 12900 23734 12952 23740
rect 12900 23248 12952 23254
rect 12900 23190 12952 23196
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12912 22234 12940 23190
rect 12900 22228 12952 22234
rect 12900 22170 12952 22176
rect 12900 21004 12952 21010
rect 12900 20946 12952 20952
rect 12912 20466 12940 20946
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12728 18970 12756 19858
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12820 18970 12848 19110
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12820 18290 12848 18702
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12544 17202 12572 17546
rect 12636 17542 12664 18226
rect 12820 17814 12848 18226
rect 12808 17808 12860 17814
rect 12808 17750 12860 17756
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12820 17338 12848 17750
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12544 16561 12572 16934
rect 12636 16726 12664 17002
rect 12820 16794 12848 17138
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12624 16720 12676 16726
rect 12624 16662 12676 16668
rect 12530 16552 12586 16561
rect 12530 16487 12586 16496
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12452 15638 12480 15914
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12348 15496 12400 15502
rect 12544 15484 12572 16487
rect 12900 15904 12952 15910
rect 12900 15846 12952 15852
rect 12348 15438 12400 15444
rect 12452 15456 12572 15484
rect 12624 15496 12676 15502
rect 12360 15094 12388 15438
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12268 14074 12296 14486
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 11992 13786 12112 13814
rect 12164 13796 12216 13802
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11808 12918 11836 13194
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11808 11150 11836 12854
rect 11900 12442 11928 13262
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11992 12322 12020 13786
rect 12164 13738 12216 13744
rect 12176 13530 12204 13738
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 11900 12294 12020 12322
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 10266 11836 11086
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11900 10033 11928 12294
rect 12084 12238 12112 12378
rect 12268 12238 12296 12582
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12268 11762 12296 12174
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12360 11354 12388 11766
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12452 11268 12480 15456
rect 12624 15438 12676 15444
rect 12636 14550 12664 15438
rect 12912 15366 12940 15846
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12912 14890 12940 15302
rect 12900 14884 12952 14890
rect 12900 14826 12952 14832
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12544 13802 12572 14214
rect 12636 13802 12664 14282
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12636 13530 12664 13738
rect 13004 13530 13032 25162
rect 13556 24818 13584 25298
rect 14476 24886 14504 27520
rect 14740 27474 14792 27480
rect 15292 27532 15344 27538
rect 15382 27520 15438 28000
rect 16394 27520 16450 28000
rect 17406 27520 17462 28000
rect 18418 27554 18474 28000
rect 17880 27526 18474 27554
rect 15292 27474 15344 27480
rect 14556 25356 14608 25362
rect 14556 25298 14608 25304
rect 14568 24954 14596 25298
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 14096 24880 14148 24886
rect 14096 24822 14148 24828
rect 14464 24880 14516 24886
rect 14464 24822 14516 24828
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13096 18902 13124 24754
rect 13556 24721 13584 24754
rect 13542 24712 13598 24721
rect 13542 24647 13598 24656
rect 14108 24274 14136 24822
rect 14280 24608 14332 24614
rect 14280 24550 14332 24556
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14004 23792 14056 23798
rect 14108 23780 14136 24210
rect 14056 23752 14136 23780
rect 14004 23734 14056 23740
rect 14292 23730 14320 24550
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 14372 23724 14424 23730
rect 14372 23666 14424 23672
rect 14556 23724 14608 23730
rect 14556 23666 14608 23672
rect 13176 23588 13228 23594
rect 13176 23530 13228 23536
rect 14188 23588 14240 23594
rect 14188 23530 14240 23536
rect 13188 23118 13216 23530
rect 14200 23474 14228 23530
rect 14108 23446 14228 23474
rect 14108 23322 14136 23446
rect 14384 23322 14412 23666
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 13268 23248 13320 23254
rect 13268 23190 13320 23196
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13188 22166 13216 23054
rect 13280 22982 13308 23190
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13280 22778 13308 22918
rect 13268 22772 13320 22778
rect 13268 22714 13320 22720
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 13728 22500 13780 22506
rect 13728 22442 13780 22448
rect 13740 22234 13768 22442
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 13176 22160 13228 22166
rect 13176 22102 13228 22108
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 13188 21690 13216 22102
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13280 21554 13308 22034
rect 13648 21690 13676 22102
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13360 21412 13412 21418
rect 13360 21354 13412 21360
rect 13176 21072 13228 21078
rect 13176 21014 13228 21020
rect 13188 20330 13216 21014
rect 13176 20324 13228 20330
rect 13176 20266 13228 20272
rect 13188 19990 13216 20266
rect 13372 20058 13400 21354
rect 13648 20602 13676 21626
rect 13740 21146 13768 22170
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13176 19984 13228 19990
rect 13176 19926 13228 19932
rect 13912 19984 13964 19990
rect 13912 19926 13964 19932
rect 13924 19378 13952 19926
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 13832 18834 13860 19178
rect 13924 18970 13952 19314
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13082 18184 13138 18193
rect 13082 18119 13138 18128
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12544 12714 12572 13126
rect 13004 12986 13032 13466
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12544 11665 12572 12650
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12530 11656 12586 11665
rect 12530 11591 12586 11600
rect 12452 11240 12572 11268
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11886 10024 11942 10033
rect 11886 9959 11942 9968
rect 11992 9178 12020 10406
rect 12348 10192 12400 10198
rect 12348 10134 12400 10140
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12084 9722 12112 9998
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12360 9518 12388 10134
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12360 9178 12388 9454
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 12268 8022 12296 8298
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11900 7546 11928 7822
rect 12268 7546 12296 7958
rect 12452 7546 12480 9318
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 11716 6854 11836 6882
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11716 6458 11744 6734
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11532 4690 11560 6122
rect 11808 5778 11836 6854
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11532 4282 11560 4626
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 10692 4140 10744 4146
rect 10876 4140 10928 4146
rect 10744 4100 10824 4128
rect 10692 4082 10744 4088
rect 10796 3942 10824 4100
rect 10876 4082 10928 4088
rect 11072 4126 11192 4154
rect 11348 4126 11468 4154
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10796 3738 10824 3878
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9784 3194 9812 3538
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 8772 2990 8800 3130
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 6918 82 6974 480
rect 6840 54 6974 82
rect 4342 0 4398 54
rect 5630 0 5686 54
rect 6918 0 6974 54
rect 8114 96 8170 480
rect 9324 82 9352 2790
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10980 2650 11008 2790
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 9402 82 9458 480
rect 9324 54 9458 82
rect 8114 0 8170 40
rect 9402 0 9458 54
rect 10690 82 10746 480
rect 10796 82 10824 2246
rect 11072 134 11100 4126
rect 11348 3194 11376 4126
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11348 2990 11376 3130
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 10690 54 10824 82
rect 11060 128 11112 134
rect 11060 70 11112 76
rect 11978 128 12034 480
rect 12544 134 12572 11240
rect 12636 11150 12664 12106
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10674 12756 10950
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12728 10062 12756 10610
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12636 9178 12664 9386
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12728 8566 12756 9998
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12728 7750 12756 8298
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12728 7546 12756 7686
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12728 5370 12756 5714
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12820 4154 12848 10406
rect 12912 7274 12940 12922
rect 13096 9674 13124 18119
rect 13556 17814 13584 18294
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 13544 17808 13596 17814
rect 13544 17750 13596 17756
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13280 15026 13308 15302
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13280 14550 13308 14962
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 13280 13938 13308 14486
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13372 13814 13400 17478
rect 13464 17270 13492 17750
rect 13452 17264 13504 17270
rect 13452 17206 13504 17212
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13464 16250 13492 16594
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13556 14822 13584 15506
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13372 13786 13492 13814
rect 13556 13802 13584 14758
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13372 12442 13400 13262
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13372 11762 13400 12378
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13096 9646 13216 9674
rect 13188 7478 13216 9646
rect 13280 9586 13308 10542
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 13280 6934 13308 9522
rect 13372 9450 13400 9862
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 8362 13400 9386
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13372 8022 13400 8298
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13096 6254 13124 6598
rect 13176 6452 13228 6458
rect 13280 6440 13308 6870
rect 13228 6412 13308 6440
rect 13176 6394 13228 6400
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13096 5914 13124 6190
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 12636 4126 12848 4154
rect 12636 2922 12664 4126
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 13464 2650 13492 13786
rect 13544 13796 13596 13802
rect 13544 13738 13596 13744
rect 13544 13456 13596 13462
rect 13596 13416 13676 13444
rect 13544 13398 13596 13404
rect 13648 12850 13676 13416
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13648 12646 13676 12786
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 12306 13676 12582
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13648 11898 13676 12242
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13740 11121 13768 18294
rect 13832 18222 13860 18770
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13832 17814 13860 18158
rect 13912 17876 13964 17882
rect 14016 17864 14044 22374
rect 14108 22166 14136 22646
rect 14384 22642 14412 23258
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14096 22160 14148 22166
rect 14096 22102 14148 22108
rect 14108 21554 14136 22102
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14292 21350 14320 21558
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14108 20602 14136 20878
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 14108 19281 14136 19450
rect 14200 19310 14228 19994
rect 14188 19304 14240 19310
rect 14094 19272 14150 19281
rect 14188 19246 14240 19252
rect 14094 19207 14150 19216
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 14108 18086 14136 18770
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 13964 17836 14044 17864
rect 13912 17818 13964 17824
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 13924 13814 13952 17818
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 14016 14006 14044 14418
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 13832 13786 13952 13814
rect 13832 13705 13860 13786
rect 13818 13696 13874 13705
rect 13818 13631 13874 13640
rect 13726 11112 13782 11121
rect 13726 11047 13782 11056
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13740 9722 13768 10066
rect 13728 9716 13780 9722
rect 13556 9664 13728 9674
rect 13556 9658 13780 9664
rect 13556 9646 13768 9658
rect 13556 8634 13584 9646
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13648 8090 13676 8910
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13832 8022 13860 13631
rect 14108 13394 14136 18022
rect 14292 14822 14320 21286
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14292 13512 14320 14758
rect 14384 13938 14412 19110
rect 14464 18692 14516 18698
rect 14464 18634 14516 18640
rect 14476 18358 14504 18634
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14568 18204 14596 23666
rect 14648 19236 14700 19242
rect 14648 19178 14700 19184
rect 14660 18970 14688 19178
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14660 18290 14688 18906
rect 14752 18426 14780 27474
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15304 24954 15332 27474
rect 15396 25362 15424 27520
rect 15384 25356 15436 25362
rect 15384 25298 15436 25304
rect 15292 24948 15344 24954
rect 15292 24890 15344 24896
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 16408 23866 16436 27520
rect 17420 23866 17448 27520
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 17408 23860 17460 23866
rect 17408 23802 17460 23808
rect 17880 23769 17908 27526
rect 18418 27520 18474 27526
rect 19430 27520 19486 28000
rect 20442 27520 20498 28000
rect 21454 27520 21510 28000
rect 22374 27520 22430 28000
rect 23386 27520 23442 28000
rect 24398 27554 24454 28000
rect 24228 27526 24454 27554
rect 17866 23760 17922 23769
rect 17866 23695 17922 23704
rect 18604 23724 18656 23730
rect 17316 23656 17368 23662
rect 17316 23598 17368 23604
rect 16120 23180 16172 23186
rect 16120 23122 16172 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 16132 22778 16160 23122
rect 16120 22772 16172 22778
rect 16120 22714 16172 22720
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 14924 22432 14976 22438
rect 14924 22374 14976 22380
rect 15384 22432 15436 22438
rect 15384 22374 15436 22380
rect 14936 22030 14964 22374
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 14936 21146 14964 21422
rect 14924 21140 14976 21146
rect 14844 21100 14924 21128
rect 14844 20058 14872 21100
rect 14924 21082 14976 21088
rect 15396 21010 15424 22374
rect 15488 21690 15516 22510
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15660 21956 15712 21962
rect 15660 21898 15712 21904
rect 15476 21684 15528 21690
rect 15476 21626 15528 21632
rect 15568 21412 15620 21418
rect 15568 21354 15620 21360
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15106 20496 15162 20505
rect 15580 20466 15608 21354
rect 15672 21146 15700 21898
rect 15856 21418 15884 22034
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 15844 21412 15896 21418
rect 15844 21354 15896 21360
rect 16040 21146 16068 21966
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16500 21486 16528 21830
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 15660 21140 15712 21146
rect 15660 21082 15712 21088
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 15106 20431 15162 20440
rect 15568 20460 15620 20466
rect 15120 20398 15148 20431
rect 15568 20402 15620 20408
rect 15108 20392 15160 20398
rect 15108 20334 15160 20340
rect 16408 20330 16436 21082
rect 15384 20324 15436 20330
rect 15384 20266 15436 20272
rect 16396 20324 16448 20330
rect 16396 20266 16448 20272
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15396 19378 15424 20266
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14476 18176 14596 18204
rect 14476 16153 14504 18176
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14568 17134 14596 17750
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14462 16144 14518 16153
rect 14462 16079 14518 16088
rect 14568 16046 14596 16934
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14384 13530 14412 13874
rect 14200 13484 14320 13512
rect 14372 13524 14424 13530
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14108 12918 14136 13330
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13924 10266 13952 11494
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14016 10470 14044 11154
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14016 10130 14044 10406
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13924 9110 13952 9658
rect 14016 9110 14044 10066
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 13924 8634 13952 9046
rect 14108 8906 14136 12854
rect 14200 11286 14228 13484
rect 14372 13466 14424 13472
rect 14278 13424 14334 13433
rect 14278 13359 14334 13368
rect 14292 12986 14320 13359
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14188 11280 14240 11286
rect 14384 11234 14412 13466
rect 14188 11222 14240 11228
rect 14200 10742 14228 11222
rect 14292 11206 14412 11234
rect 14188 10736 14240 10742
rect 14188 10678 14240 10684
rect 14292 10198 14320 11206
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14384 10810 14412 11086
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14568 10713 14596 15982
rect 14752 14482 14780 18362
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 15212 17678 15240 18090
rect 15396 18086 15424 18294
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15396 16980 15424 18022
rect 15488 17882 15516 20198
rect 16408 20058 16436 20266
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16500 19922 16528 21286
rect 16960 20058 16988 21286
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 15568 19304 15620 19310
rect 15568 19246 15620 19252
rect 15580 18902 15608 19246
rect 16132 18970 16160 19858
rect 16304 19236 16356 19242
rect 16304 19178 16356 19184
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16224 18222 16252 18702
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15672 17338 15700 18022
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 16224 17202 16252 18158
rect 16316 17814 16344 19178
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16592 18970 16620 19110
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 17132 18148 17184 18154
rect 17132 18090 17184 18096
rect 16304 17808 16356 17814
rect 16304 17750 16356 17756
rect 16316 17338 16344 17750
rect 17144 17542 17172 18090
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15476 16992 15528 16998
rect 15396 16952 15476 16980
rect 15476 16934 15528 16940
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15304 16561 15332 16594
rect 15290 16552 15346 16561
rect 15290 16487 15346 16496
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14844 16046 14872 16390
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16250 15332 16487
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14844 14958 14872 15982
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 15028 15706 15056 15914
rect 15488 15910 15516 16934
rect 16040 16454 16068 17070
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 16776 16794 16804 17002
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 16028 16448 16080 16454
rect 16028 16390 16080 16396
rect 15856 16046 15884 16390
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14844 14618 14872 14894
rect 15488 14822 15516 15846
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14844 14074 14872 14554
rect 15488 14550 15516 14758
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14844 13870 14872 14010
rect 15304 13938 15332 14350
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14646 13424 14702 13433
rect 14646 13359 14702 13368
rect 14660 12889 14688 13359
rect 14646 12880 14702 12889
rect 14646 12815 14702 12824
rect 14844 11762 14872 13670
rect 15304 13530 15332 13874
rect 15488 13734 15516 14486
rect 15856 13734 15884 15982
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15844 13728 15896 13734
rect 15948 13705 15976 13806
rect 15844 13670 15896 13676
rect 15934 13696 15990 13705
rect 15934 13631 15990 13640
rect 15948 13530 15976 13631
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 16040 13462 16068 16390
rect 16960 16250 16988 16662
rect 17052 16250 17080 16934
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 16224 15706 16252 15914
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16500 14618 16528 14894
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16396 13864 16448 13870
rect 17144 13814 17172 17478
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17236 14550 17264 16458
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 16396 13806 16448 13812
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 16408 13394 16436 13806
rect 17052 13786 17172 13814
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15948 12986 15976 13330
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 16500 12850 16528 13194
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 15660 12708 15712 12714
rect 15660 12650 15712 12656
rect 15028 12442 15056 12650
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15396 11898 15424 12378
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15672 11762 15700 12650
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14554 10704 14610 10713
rect 14844 10674 14872 10950
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15672 10674 15700 11698
rect 15948 11694 15976 12310
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15948 11286 15976 11630
rect 16224 11558 16252 12582
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15948 10810 15976 11222
rect 16224 11014 16252 11494
rect 16592 11354 16620 12106
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16856 11620 16908 11626
rect 16856 11562 16908 11568
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16868 11014 16896 11562
rect 16960 11286 16988 12038
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 14554 10639 14610 10648
rect 14832 10668 14884 10674
rect 14280 10192 14332 10198
rect 14280 10134 14332 10140
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14200 9178 14228 9386
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14568 9042 14596 10639
rect 14832 10610 14884 10616
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15948 10266 15976 10746
rect 16224 10538 16252 10950
rect 16762 10568 16818 10577
rect 16212 10532 16264 10538
rect 16762 10503 16818 10512
rect 16212 10474 16264 10480
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 14096 8900 14148 8906
rect 14096 8842 14148 8848
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8634 15332 8978
rect 15396 8838 15424 9998
rect 15948 9722 15976 10202
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15948 9178 15976 9454
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15752 8900 15804 8906
rect 15752 8842 15804 8848
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14200 7562 14228 7890
rect 14292 7750 14320 8298
rect 15396 8090 15424 8774
rect 15764 8430 15792 8842
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15948 8294 15976 9114
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16316 8430 16344 8978
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 16316 8090 16344 8366
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15844 7948 15896 7954
rect 15844 7890 15896 7896
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14200 7534 14320 7562
rect 14292 7410 14320 7534
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14292 7313 14320 7346
rect 14278 7304 14334 7313
rect 14278 7239 14334 7248
rect 14660 7002 14688 7686
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15672 7206 15700 7890
rect 15856 7546 15884 7890
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13832 6458 13860 6802
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 13818 3360 13874 3369
rect 13818 3295 13874 3304
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13832 2514 13860 3295
rect 13176 2508 13228 2514
rect 13176 2450 13228 2456
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 13188 2417 13216 2450
rect 13174 2408 13230 2417
rect 13174 2343 13230 2352
rect 13188 2310 13216 2343
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 11978 76 11980 128
rect 12032 76 12034 128
rect 10690 0 10746 54
rect 11978 0 12034 76
rect 12532 128 12584 134
rect 12532 70 12584 76
rect 13266 128 13322 480
rect 13266 76 13268 128
rect 13320 76 13322 128
rect 13266 0 13322 76
rect 14554 82 14610 480
rect 14660 82 14688 6326
rect 15672 6225 15700 7142
rect 15658 6216 15714 6225
rect 15658 6151 15714 6160
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15764 2514 15792 7278
rect 16776 4154 16804 10503
rect 16868 10266 16896 10950
rect 16960 10810 16988 11222
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 9110 16896 9318
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 16868 8634 16896 9046
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 17052 8566 17080 13786
rect 17236 13530 17264 14486
rect 17328 13814 17356 23598
rect 17408 22160 17460 22166
rect 17408 22102 17460 22108
rect 17420 21350 17448 22102
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17592 21412 17644 21418
rect 17592 21354 17644 21360
rect 17408 21344 17460 21350
rect 17408 21286 17460 21292
rect 17604 19514 17632 21354
rect 17696 21078 17724 21966
rect 17776 21344 17828 21350
rect 17776 21286 17828 21292
rect 17788 21146 17816 21286
rect 17776 21140 17828 21146
rect 17776 21082 17828 21088
rect 17684 21072 17736 21078
rect 17684 21014 17736 21020
rect 17696 20466 17724 21014
rect 17880 20534 17908 23695
rect 18604 23666 18656 23672
rect 18512 23656 18564 23662
rect 18512 23598 18564 23604
rect 18328 22092 18380 22098
rect 18328 22034 18380 22040
rect 18340 21418 18368 22034
rect 18144 21412 18196 21418
rect 18144 21354 18196 21360
rect 18328 21412 18380 21418
rect 18328 21354 18380 21360
rect 18156 20942 18184 21354
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 17868 20528 17920 20534
rect 17868 20470 17920 20476
rect 17684 20460 17736 20466
rect 17684 20402 17736 20408
rect 18156 20330 18184 20742
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 18328 20324 18380 20330
rect 18328 20266 18380 20272
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17512 16658 17540 17818
rect 17604 17746 17632 19450
rect 17788 18884 17816 20198
rect 18156 20058 18184 20266
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18340 19990 18368 20266
rect 18328 19984 18380 19990
rect 18248 19944 18328 19972
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17880 19514 17908 19790
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 18248 18970 18276 19944
rect 18328 19926 18380 19932
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 18340 18970 18368 19178
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18328 18964 18380 18970
rect 18328 18906 18380 18912
rect 17868 18896 17920 18902
rect 17788 18856 17868 18884
rect 17868 18838 17920 18844
rect 17880 18426 17908 18838
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 18064 17882 18092 18702
rect 18248 18154 18276 18906
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18432 18290 18460 18702
rect 18524 18698 18552 23598
rect 18616 23322 18644 23666
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 19444 22778 19472 27520
rect 20166 26480 20222 26489
rect 20166 26415 20222 26424
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19984 23588 20036 23594
rect 19984 23530 20036 23536
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19156 22432 19208 22438
rect 19156 22374 19208 22380
rect 19168 22234 19196 22374
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19156 22228 19208 22234
rect 19156 22170 19208 22176
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19536 21146 19564 21286
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19524 21140 19576 21146
rect 19524 21082 19576 21088
rect 18972 21072 19024 21078
rect 18972 21014 19024 21020
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18892 19990 18920 20402
rect 18984 20262 19012 21014
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 19260 19990 19288 20878
rect 19536 20466 19564 21082
rect 19524 20460 19576 20466
rect 19524 20402 19576 20408
rect 19522 20360 19578 20369
rect 19340 20324 19392 20330
rect 19522 20295 19578 20304
rect 19340 20266 19392 20272
rect 18880 19984 18932 19990
rect 18880 19926 18932 19932
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 18788 19372 18840 19378
rect 18892 19360 18920 19926
rect 19352 19514 19380 20266
rect 19536 20262 19564 20295
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 19514 19472 19654
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 18840 19332 18920 19360
rect 18788 19314 18840 19320
rect 19338 19272 19394 19281
rect 19338 19207 19394 19216
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 19260 18358 19288 18770
rect 19352 18698 19380 19207
rect 19444 18766 19472 19450
rect 19720 19310 19748 19858
rect 19708 19304 19760 19310
rect 19706 19272 19708 19281
rect 19760 19272 19762 19281
rect 19706 19207 19762 19216
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19248 18352 19300 18358
rect 19248 18294 19300 18300
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18236 18148 18288 18154
rect 18236 18090 18288 18096
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 18432 17814 18460 18226
rect 18420 17808 18472 17814
rect 18420 17750 18472 17756
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 17604 16998 17632 17682
rect 17592 16992 17644 16998
rect 17592 16934 17644 16940
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17512 16182 17540 16594
rect 17500 16176 17552 16182
rect 17500 16118 17552 16124
rect 17408 15632 17460 15638
rect 17408 15574 17460 15580
rect 17420 15366 17448 15574
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17420 15162 17448 15302
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17420 14278 17448 14486
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17420 14074 17448 14214
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17328 13786 17448 13814
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17144 11150 17172 12718
rect 17328 12628 17356 13330
rect 17420 12918 17448 13786
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17408 12640 17460 12646
rect 17328 12600 17408 12628
rect 17408 12582 17460 12588
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17236 11762 17264 12038
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17420 11626 17448 12582
rect 17512 12442 17540 12582
rect 17604 12442 17632 16934
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17316 11620 17368 11626
rect 17316 11562 17368 11568
rect 17408 11620 17460 11626
rect 17408 11562 17460 11568
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17144 10266 17172 11086
rect 17328 11082 17356 11562
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17696 10418 17724 16934
rect 17788 16454 17816 17682
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18616 17066 18644 17478
rect 18984 17202 19012 17478
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18604 17060 18656 17066
rect 18604 17002 18656 17008
rect 18616 16794 18644 17002
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18892 16726 18920 17070
rect 18696 16720 18748 16726
rect 18696 16662 18748 16668
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 17788 15094 17816 16390
rect 18064 16114 18092 16390
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17776 15088 17828 15094
rect 17776 15030 17828 15036
rect 17788 13870 17816 15030
rect 17880 14550 17908 15302
rect 17972 15162 18000 15438
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18156 15026 18184 15302
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 18156 14618 18184 14826
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 17868 14544 17920 14550
rect 17868 14486 17920 14492
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 18064 13530 18092 14486
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18156 13802 18184 14350
rect 18248 14346 18276 16050
rect 18340 15978 18368 16186
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 18432 15434 18460 16526
rect 18708 16250 18736 16662
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18892 16114 18920 16662
rect 18984 16114 19012 17138
rect 19168 16998 19196 17682
rect 19156 16992 19208 16998
rect 19156 16934 19208 16940
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18972 16108 19024 16114
rect 18972 16050 19024 16056
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18892 15638 18920 15846
rect 18880 15632 18932 15638
rect 18880 15574 18932 15580
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 18432 15026 18460 15370
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18236 14340 18288 14346
rect 18236 14282 18288 14288
rect 18248 13938 18276 14282
rect 18340 14074 18368 14826
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18234 13832 18290 13841
rect 18144 13796 18196 13802
rect 18340 13802 18368 14010
rect 18432 13841 18460 14554
rect 18892 14550 18920 15574
rect 19260 14550 19288 18294
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 19248 14544 19300 14550
rect 19248 14486 19300 14492
rect 18892 14074 18920 14486
rect 19248 14340 19300 14346
rect 19248 14282 19300 14288
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18418 13832 18474 13841
rect 18234 13767 18290 13776
rect 18328 13796 18380 13802
rect 18144 13738 18196 13744
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 18248 13462 18276 13767
rect 18418 13767 18474 13776
rect 18328 13738 18380 13744
rect 19260 13462 19288 14282
rect 19352 13814 19380 18090
rect 19536 18086 19564 19110
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19536 17882 19564 18022
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19996 17338 20024 23530
rect 20180 21690 20208 26415
rect 20456 23866 20484 27520
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 21468 23633 21496 27520
rect 22388 23798 22416 27520
rect 23400 24410 23428 27520
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 24228 23866 24256 27526
rect 24398 27520 24454 27526
rect 25410 27520 25466 28000
rect 26422 27532 26478 28000
rect 26422 27520 26424 27532
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24674 24712 24730 24721
rect 24674 24647 24730 24656
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24216 23860 24268 23866
rect 24216 23802 24268 23808
rect 22376 23792 22428 23798
rect 22376 23734 22428 23740
rect 21454 23624 21510 23633
rect 21454 23559 21510 23568
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24122 22400 24178 22409
rect 24122 22335 24178 22344
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 20180 21486 20208 21626
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 20076 21412 20128 21418
rect 20076 21354 20128 21360
rect 20088 19378 20116 21354
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20548 20942 20576 21286
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20352 20868 20404 20874
rect 20352 20810 20404 20816
rect 20364 20330 20392 20810
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20352 20324 20404 20330
rect 20352 20266 20404 20272
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20076 19236 20128 19242
rect 20076 19178 20128 19184
rect 20088 18970 20116 19178
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 20364 18290 20392 20266
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19522 17232 19578 17241
rect 19522 17167 19578 17176
rect 19536 16794 19564 17167
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19536 15960 19564 16730
rect 20718 16144 20774 16153
rect 19984 16108 20036 16114
rect 20718 16079 20774 16088
rect 19984 16050 20036 16056
rect 19616 15972 19668 15978
rect 19536 15932 19616 15960
rect 19616 15914 19668 15920
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19444 14822 19472 15506
rect 19996 15026 20024 16050
rect 20076 15972 20128 15978
rect 20076 15914 20128 15920
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19812 14890 19840 14962
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19800 14884 19852 14890
rect 19800 14826 19852 14832
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19536 14278 19564 14826
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 20088 14618 20116 15914
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19812 14074 19840 14214
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19352 13786 19564 13814
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19444 13530 19472 13670
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18156 12850 18184 13126
rect 18524 12986 18552 13398
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19444 12986 19472 13262
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 17960 12776 18012 12782
rect 17774 12744 17830 12753
rect 17960 12718 18012 12724
rect 17774 12679 17830 12688
rect 17788 12374 17816 12679
rect 17972 12646 18000 12718
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17788 11286 17816 12310
rect 17880 11558 17908 12310
rect 18248 11626 18276 12650
rect 18512 12164 18564 12170
rect 18512 12106 18564 12112
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 18248 11354 18276 11562
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17604 10390 17724 10418
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17236 8974 17264 9522
rect 17328 8974 17356 9998
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 17236 8090 17264 8910
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17604 7313 17632 10390
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17696 9518 17724 10202
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17880 9110 17908 10950
rect 18432 10674 18460 12038
rect 18524 11626 18552 12106
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18800 11898 18828 12038
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18892 11665 18920 12038
rect 18984 11830 19012 12786
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 18972 11688 19024 11694
rect 18878 11656 18934 11665
rect 18512 11620 18564 11626
rect 18972 11630 19024 11636
rect 18878 11591 18934 11600
rect 18512 11562 18564 11568
rect 18420 10668 18472 10674
rect 18420 10610 18472 10616
rect 18236 10532 18288 10538
rect 18288 10492 18368 10520
rect 18236 10474 18288 10480
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17972 10266 18000 10406
rect 18340 10266 18368 10492
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18340 9722 18368 10202
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18340 9450 18368 9658
rect 18524 9586 18552 11562
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18708 10810 18736 11086
rect 18696 10804 18748 10810
rect 18696 10746 18748 10752
rect 18708 10198 18736 10746
rect 18984 10577 19012 11630
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 19076 10742 19104 11222
rect 19168 11014 19196 12786
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19260 11762 19288 12242
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19444 11354 19472 12242
rect 19432 11348 19484 11354
rect 19352 11308 19432 11336
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 18970 10568 19026 10577
rect 18970 10503 19026 10512
rect 19076 10266 19104 10678
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 18696 10192 18748 10198
rect 18696 10134 18748 10140
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19260 9722 19288 9998
rect 19248 9716 19300 9722
rect 19248 9658 19300 9664
rect 19260 9625 19288 9658
rect 19246 9616 19302 9625
rect 18512 9580 18564 9586
rect 19246 9551 19302 9560
rect 18512 9522 18564 9528
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18248 9178 18276 9386
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 17866 8528 17922 8537
rect 17866 8463 17922 8472
rect 17880 8430 17908 8463
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17590 7304 17646 7313
rect 17590 7239 17646 7248
rect 17880 6866 17908 8366
rect 18800 8294 18828 8978
rect 19352 8498 19380 11308
rect 19432 11290 19484 11296
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 19444 10169 19472 10542
rect 19430 10160 19486 10169
rect 19430 10095 19486 10104
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 18788 8288 18840 8294
rect 18788 8230 18840 8236
rect 18800 7449 18828 8230
rect 18786 7440 18842 7449
rect 18786 7375 18842 7384
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 16776 4126 16896 4154
rect 16868 2514 16896 4126
rect 19536 2650 19564 13786
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19800 11280 19852 11286
rect 19800 11222 19852 11228
rect 19812 10810 19840 11222
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4154 20024 14486
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20074 13968 20130 13977
rect 20074 13903 20130 13912
rect 20088 13870 20116 13903
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 20088 12753 20116 13670
rect 20180 13190 20208 14214
rect 20272 13433 20300 14758
rect 20732 13814 20760 16079
rect 20824 14482 20852 20470
rect 21364 16448 21416 16454
rect 21364 16390 21416 16396
rect 21376 16114 21404 16390
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20824 14006 20852 14418
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20732 13786 20852 13814
rect 20258 13424 20314 13433
rect 20824 13394 20852 13786
rect 20258 13359 20314 13368
rect 20812 13388 20864 13394
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20074 12744 20130 12753
rect 20074 12679 20130 12688
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 20180 9625 20208 12582
rect 20272 11218 20300 13359
rect 20812 13330 20864 13336
rect 20824 12986 20852 13330
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 21192 12889 21220 14894
rect 24136 13814 24164 22335
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 17128 24268 17134
rect 24216 17070 24268 17076
rect 24228 14385 24256 17070
rect 24688 16658 24716 24647
rect 25424 21690 25452 27520
rect 26476 27520 26478 27532
rect 27434 27520 27490 28000
rect 26424 27474 26476 27480
rect 26436 27443 26464 27474
rect 27342 24848 27398 24857
rect 27448 24834 27476 27520
rect 27398 24806 27476 24834
rect 27342 24783 27398 24792
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25134 20632 25190 20641
rect 25134 20567 25190 20576
rect 25148 20534 25176 20567
rect 25136 20528 25188 20534
rect 25136 20470 25188 20476
rect 27620 17264 27672 17270
rect 27620 17206 27672 17212
rect 27632 16969 27660 17206
rect 27618 16960 27674 16969
rect 27618 16895 27674 16904
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16250 24716 16594
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24766 14648 24822 14657
rect 24766 14583 24822 14592
rect 24214 14376 24270 14385
rect 24780 14346 24808 14583
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24214 14311 24270 14320
rect 24768 14340 24820 14346
rect 24768 14282 24820 14288
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 25056 14074 25084 14418
rect 25044 14068 25096 14074
rect 25044 14010 25096 14016
rect 24136 13786 24256 13814
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23860 13297 23888 13330
rect 23846 13288 23902 13297
rect 23846 13223 23902 13232
rect 23860 12986 23888 13223
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 21178 12880 21234 12889
rect 21178 12815 21234 12824
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 21468 11558 21496 12242
rect 23860 11898 23888 12242
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23860 11801 23888 11834
rect 23846 11792 23902 11801
rect 23846 11727 23902 11736
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 21376 10810 21404 11154
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21468 10033 21496 11494
rect 24044 11218 24072 13126
rect 24124 12096 24176 12102
rect 24124 12038 24176 12044
rect 24136 11694 24164 12038
rect 24124 11688 24176 11694
rect 24124 11630 24176 11636
rect 24032 11212 24084 11218
rect 24032 11154 24084 11160
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 21454 10024 21510 10033
rect 21454 9959 21510 9968
rect 20166 9616 20222 9625
rect 20166 9551 20222 9560
rect 19996 4126 20116 4154
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 20088 2514 20116 4126
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 15752 2508 15804 2514
rect 15752 2450 15804 2456
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 20626 2408 20682 2417
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14554 54 14688 82
rect 15488 82 15516 2314
rect 15750 82 15806 480
rect 15488 54 15806 82
rect 16776 82 16804 2314
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 17038 82 17094 480
rect 16776 54 17094 82
rect 18064 82 18092 2246
rect 18326 82 18382 480
rect 18708 105 18736 2246
rect 18064 54 18382 82
rect 14554 0 14610 54
rect 15750 0 15806 54
rect 17038 0 17094 54
rect 18326 0 18382 54
rect 18694 96 18750 105
rect 19444 82 19472 2382
rect 20626 2343 20682 2352
rect 19614 82 19670 480
rect 19444 54 19670 82
rect 20640 82 20668 2343
rect 20902 82 20958 480
rect 20640 54 20958 82
rect 21744 82 21772 3878
rect 22098 82 22154 480
rect 22204 134 22232 10950
rect 24228 2514 24256 13786
rect 26240 13796 26292 13802
rect 26240 13738 26292 13744
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24766 12472 24822 12481
rect 24766 12407 24822 12416
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24780 11898 24808 12407
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 25504 11620 25556 11626
rect 25504 11562 25556 11568
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24780 11257 24808 11290
rect 24766 11248 24822 11257
rect 24676 11212 24728 11218
rect 24766 11183 24822 11192
rect 24676 11154 24728 11160
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24688 10810 24716 11154
rect 24676 10804 24728 10810
rect 24676 10746 24728 10752
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 25516 7041 25544 11562
rect 25502 7032 25558 7041
rect 25502 6967 25558 6976
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 26056 2440 26108 2446
rect 26056 2382 26108 2388
rect 24860 2372 24912 2378
rect 24860 2314 24912 2320
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 21744 54 22154 82
rect 22192 128 22244 134
rect 22192 70 22244 76
rect 23386 128 23442 480
rect 23386 76 23388 128
rect 23440 76 23442 128
rect 18694 31 18750 40
rect 19614 0 19670 54
rect 20902 0 20958 54
rect 22098 0 22154 54
rect 23386 0 23442 76
rect 24674 82 24730 480
rect 24872 82 24900 2314
rect 24674 54 24900 82
rect 25962 82 26018 480
rect 26068 82 26096 2382
rect 26252 134 26280 13738
rect 27710 7440 27766 7449
rect 27710 7375 27766 7384
rect 27618 7304 27674 7313
rect 27618 7239 27674 7248
rect 27632 5001 27660 7239
rect 27618 4992 27674 5001
rect 27618 4927 27674 4936
rect 27724 1057 27752 7375
rect 27710 1048 27766 1057
rect 27710 983 27766 992
rect 25962 54 26096 82
rect 26240 128 26292 134
rect 26240 70 26292 76
rect 27250 128 27306 480
rect 27250 76 27252 128
rect 27304 76 27306 128
rect 24674 0 24730 54
rect 25962 0 26018 54
rect 27250 0 27306 76
<< via2 >>
rect 18 24248 74 24304
rect 18 19760 74 19816
rect 1122 26696 1178 26752
rect 1214 25200 1270 25256
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 1582 22208 1638 22264
rect 1582 17176 1638 17232
rect 1582 16632 1638 16688
rect 1306 15952 1362 16008
rect 1214 13640 1270 13696
rect 2226 13912 2282 13968
rect 2410 13912 2466 13968
rect 2134 12960 2190 13016
rect 110 6568 166 6624
rect 2778 20712 2834 20768
rect 3054 18128 3110 18184
rect 2686 10104 2742 10160
rect 2042 9288 2098 9344
rect 1858 7520 1914 7576
rect 1306 5616 1362 5672
rect 4802 20304 4858 20360
rect 3606 13504 3662 13560
rect 3882 13232 3938 13288
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 7470 20440 7526 20496
rect 7286 17856 7342 17912
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 4158 9152 4214 9208
rect 5446 13912 5502 13968
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 4710 11092 4712 11112
rect 4712 11092 4764 11112
rect 4764 11092 4766 11112
rect 4710 11056 4766 11092
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 7286 16088 7342 16144
rect 6550 10512 6606 10568
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5078 4120 5134 4176
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5538 2624 5594 2680
rect 4526 1264 4582 1320
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7562 11736 7618 11792
rect 7470 10104 7526 10160
rect 9402 23704 9458 23760
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 7746 9288 7802 9344
rect 8206 9152 8262 9208
rect 7746 6160 7802 6216
rect 9218 13776 9274 13832
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 11150 19216 11206 19272
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 11150 13776 11206 13832
rect 10966 12688 11022 12744
rect 9034 10648 9090 10704
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 11150 9968 11206 10024
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 8666 3304 8722 3360
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 11794 14320 11850 14376
rect 12622 23432 12678 23488
rect 12530 16496 12586 16552
rect 13542 24656 13598 24712
rect 13082 18128 13138 18184
rect 12530 11600 12586 11656
rect 11886 9968 11942 10024
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 8114 40 8170 96
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 14094 19216 14150 19272
rect 13818 13640 13874 13696
rect 13726 11056 13782 11112
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 17866 23704 17922 23760
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15106 20440 15162 20496
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14462 16088 14518 16144
rect 14278 13368 14334 13424
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15290 16496 15346 16552
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14646 13368 14702 13424
rect 14646 12824 14702 12880
rect 15934 13640 15990 13696
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14554 10648 14610 10704
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 16762 10512 16818 10568
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14278 7248 14334 7304
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 13818 3304 13874 3360
rect 13174 2352 13230 2408
rect 15658 6160 15714 6216
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 20166 26424 20222 26480
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19522 20304 19578 20360
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19338 19216 19394 19272
rect 19706 19252 19708 19272
rect 19708 19252 19760 19272
rect 19760 19252 19762 19272
rect 19706 19216 19762 19252
rect 18234 13776 18290 13832
rect 18418 13776 18474 13832
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24674 24656 24730 24712
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 21454 23568 21510 23624
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24122 22344 24178 22400
rect 19522 17176 19578 17232
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20718 16088 20774 16144
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 17774 12688 17830 12744
rect 18878 11600 18934 11656
rect 18970 10512 19026 10568
rect 19246 9560 19302 9616
rect 17866 8472 17922 8528
rect 17590 7248 17646 7304
rect 19430 10104 19486 10160
rect 18786 7384 18842 7440
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 20074 13912 20130 13968
rect 20258 13368 20314 13424
rect 20074 12688 20130 12744
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 27342 24792 27398 24848
rect 25134 20576 25190 20632
rect 27618 16904 27674 16960
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24766 14592 24822 14648
rect 24214 14320 24270 14376
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 23846 13232 23902 13288
rect 21178 12824 21234 12880
rect 23846 11736 23902 11792
rect 21454 9968 21510 10024
rect 20166 9560 20222 9616
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 18694 40 18750 96
rect 20626 2352 20682 2408
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24766 12416 24822 12472
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24766 11192 24822 11248
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 25502 6976 25558 7032
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 27710 7384 27766 7440
rect 27618 7248 27674 7304
rect 27618 4936 27674 4992
rect 27710 992 27766 1048
<< metal3 >>
rect 0 27208 480 27328
rect 62 26754 122 27208
rect 27520 26936 28000 27056
rect 1117 26754 1183 26757
rect 62 26752 1183 26754
rect 62 26696 1122 26752
rect 1178 26696 1183 26752
rect 62 26694 1183 26696
rect 1117 26691 1183 26694
rect 20161 26482 20227 26485
rect 27662 26482 27722 26936
rect 20161 26480 27722 26482
rect 20161 26424 20166 26480
rect 20222 26424 27722 26480
rect 20161 26422 27722 26424
rect 20161 26419 20227 26422
rect 0 25712 480 25832
rect 62 25258 122 25712
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 1209 25258 1275 25261
rect 62 25256 1275 25258
rect 62 25200 1214 25256
rect 1270 25200 1275 25256
rect 62 25198 1275 25200
rect 1209 25195 1275 25198
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 27520 24896 28000 25016
rect 27337 24850 27403 24853
rect 19290 24848 27403 24850
rect 19290 24792 27342 24848
rect 27398 24792 27403 24848
rect 19290 24790 27403 24792
rect 13537 24714 13603 24717
rect 19290 24714 19350 24790
rect 27337 24787 27403 24790
rect 13537 24712 19350 24714
rect 13537 24656 13542 24712
rect 13598 24656 19350 24712
rect 13537 24654 19350 24656
rect 24669 24714 24735 24717
rect 27662 24714 27722 24896
rect 24669 24712 27722 24714
rect 24669 24656 24674 24712
rect 24730 24656 27722 24712
rect 24669 24654 27722 24656
rect 13537 24651 13603 24654
rect 24669 24651 24735 24654
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24304 480 24336
rect 0 24248 18 24304
rect 74 24248 480 24304
rect 0 24216 480 24248
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 9397 23762 9463 23765
rect 17861 23762 17927 23765
rect 9397 23760 17927 23762
rect 9397 23704 9402 23760
rect 9458 23704 17866 23760
rect 17922 23704 17927 23760
rect 9397 23702 17927 23704
rect 9397 23699 9463 23702
rect 17861 23699 17927 23702
rect 21449 23626 21515 23629
rect 13770 23624 21515 23626
rect 13770 23568 21454 23624
rect 21510 23568 21515 23624
rect 13770 23566 21515 23568
rect 12617 23490 12683 23493
rect 13770 23490 13830 23566
rect 21449 23563 21515 23566
rect 12617 23488 13830 23490
rect 12617 23432 12622 23488
rect 12678 23432 13830 23488
rect 12617 23430 13830 23432
rect 12617 23427 12683 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 5610 22880 5930 22881
rect 0 22720 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 27520 22856 28000 22976
rect 24277 22815 24597 22816
rect 62 22266 122 22720
rect 24117 22402 24183 22405
rect 27662 22402 27722 22856
rect 24117 22400 27722 22402
rect 24117 22344 24122 22400
rect 24178 22344 27722 22400
rect 24117 22342 27722 22344
rect 24117 22339 24183 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 1577 22266 1643 22269
rect 62 22264 1643 22266
rect 62 22208 1582 22264
rect 1638 22208 1643 22264
rect 62 22206 1643 22208
rect 1577 22203 1643 22206
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21224 480 21344
rect 10277 21248 10597 21249
rect 62 20770 122 21224
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 27520 20952 28000 21072
rect 2773 20770 2839 20773
rect 62 20768 2839 20770
rect 62 20712 2778 20768
rect 2834 20712 2839 20768
rect 62 20710 2839 20712
rect 2773 20707 2839 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 25129 20634 25195 20637
rect 27662 20634 27722 20952
rect 25129 20632 27722 20634
rect 25129 20576 25134 20632
rect 25190 20576 27722 20632
rect 25129 20574 27722 20576
rect 25129 20571 25195 20574
rect 7465 20498 7531 20501
rect 15101 20498 15167 20501
rect 7465 20496 15167 20498
rect 7465 20440 7470 20496
rect 7526 20440 15106 20496
rect 15162 20440 15167 20496
rect 7465 20438 15167 20440
rect 7465 20435 7531 20438
rect 15101 20435 15167 20438
rect 4797 20362 4863 20365
rect 19517 20362 19583 20365
rect 4797 20360 19583 20362
rect 4797 20304 4802 20360
rect 4858 20304 19522 20360
rect 19578 20304 19583 20360
rect 4797 20302 19583 20304
rect 4797 20299 4863 20302
rect 19517 20299 19583 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 19816 480 19848
rect 0 19760 18 19816
rect 74 19760 480 19816
rect 0 19728 480 19760
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 11145 19274 11211 19277
rect 14089 19274 14155 19277
rect 11145 19272 14155 19274
rect 11145 19216 11150 19272
rect 11206 19216 14094 19272
rect 14150 19216 14155 19272
rect 11145 19214 14155 19216
rect 11145 19211 11211 19214
rect 14089 19211 14155 19214
rect 19333 19274 19399 19277
rect 19701 19274 19767 19277
rect 19333 19272 19767 19274
rect 19333 19216 19338 19272
rect 19394 19216 19706 19272
rect 19762 19216 19767 19272
rect 19333 19214 19767 19216
rect 19333 19211 19399 19214
rect 19701 19211 19767 19214
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 27520 18912 28000 19032
rect 5610 18528 5930 18529
rect 0 18368 480 18488
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 62 17914 122 18368
rect 3049 18186 3115 18189
rect 13077 18186 13143 18189
rect 27662 18186 27722 18912
rect 3049 18184 27722 18186
rect 3049 18128 3054 18184
rect 3110 18128 13082 18184
rect 13138 18128 27722 18184
rect 3049 18126 27722 18128
rect 3049 18123 3115 18126
rect 13077 18123 13143 18126
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 7281 17914 7347 17917
rect 62 17912 7347 17914
rect 62 17856 7286 17912
rect 7342 17856 7347 17912
rect 62 17854 7347 17856
rect 7281 17851 7347 17854
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 1577 17234 1643 17237
rect 19517 17234 19583 17237
rect 1577 17232 19583 17234
rect 1577 17176 1582 17232
rect 1638 17176 19522 17232
rect 19578 17176 19583 17232
rect 1577 17174 19583 17176
rect 1577 17171 1643 17174
rect 19517 17171 19583 17174
rect 0 16964 480 16992
rect 0 16900 60 16964
rect 124 16900 480 16964
rect 0 16872 480 16900
rect 27520 16960 28000 16992
rect 27520 16904 27618 16960
rect 27674 16904 28000 16960
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 27520 16872 28000 16904
rect 19610 16831 19930 16832
rect 54 16628 60 16692
rect 124 16690 130 16692
rect 1577 16690 1643 16693
rect 124 16688 1643 16690
rect 124 16632 1582 16688
rect 1638 16632 1643 16688
rect 124 16630 1643 16632
rect 124 16628 130 16630
rect 1577 16627 1643 16630
rect 12525 16554 12591 16557
rect 15285 16554 15351 16557
rect 12525 16552 15351 16554
rect 12525 16496 12530 16552
rect 12586 16496 15290 16552
rect 15346 16496 15351 16552
rect 12525 16494 15351 16496
rect 12525 16491 12591 16494
rect 15285 16491 15351 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 7281 16146 7347 16149
rect 14457 16146 14523 16149
rect 20713 16146 20779 16149
rect 7281 16144 20779 16146
rect 7281 16088 7286 16144
rect 7342 16088 14462 16144
rect 14518 16088 20718 16144
rect 20774 16088 20779 16144
rect 7281 16086 20779 16088
rect 7281 16083 7347 16086
rect 14457 16083 14523 16086
rect 20713 16083 20779 16086
rect 1301 16010 1367 16013
rect 62 16008 1367 16010
rect 62 15952 1306 16008
rect 1362 15952 1367 16008
rect 62 15950 1367 15952
rect 62 15496 122 15950
rect 1301 15947 1367 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 0 15376 480 15496
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 27520 14968 28000 15088
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 24761 14650 24827 14653
rect 27662 14650 27722 14968
rect 24761 14648 27722 14650
rect 24761 14592 24766 14648
rect 24822 14592 27722 14648
rect 24761 14590 27722 14592
rect 24761 14587 24827 14590
rect 11789 14378 11855 14381
rect 24209 14378 24275 14381
rect 11789 14376 24275 14378
rect 11789 14320 11794 14376
rect 11850 14320 24214 14376
rect 24270 14320 24275 14376
rect 11789 14318 24275 14320
rect 11789 14315 11855 14318
rect 24209 14315 24275 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13880 480 14000
rect 2221 13970 2287 13973
rect 2405 13970 2471 13973
rect 2221 13968 2471 13970
rect 2221 13912 2226 13968
rect 2282 13912 2410 13968
rect 2466 13912 2471 13968
rect 2221 13910 2471 13912
rect 2221 13907 2287 13910
rect 2405 13907 2471 13910
rect 5441 13970 5507 13973
rect 20069 13970 20135 13973
rect 5441 13968 20135 13970
rect 5441 13912 5446 13968
rect 5502 13912 20074 13968
rect 20130 13912 20135 13968
rect 5441 13910 20135 13912
rect 5441 13907 5507 13910
rect 20069 13907 20135 13910
rect 62 13698 122 13880
rect 9213 13834 9279 13837
rect 11145 13834 11211 13837
rect 9213 13832 11211 13834
rect 9213 13776 9218 13832
rect 9274 13776 11150 13832
rect 11206 13776 11211 13832
rect 9213 13774 11211 13776
rect 9213 13771 9279 13774
rect 11145 13771 11211 13774
rect 18229 13834 18295 13837
rect 18413 13834 18479 13837
rect 18229 13832 18479 13834
rect 18229 13776 18234 13832
rect 18290 13776 18418 13832
rect 18474 13776 18479 13832
rect 18229 13774 18479 13776
rect 18229 13771 18295 13774
rect 18413 13771 18479 13774
rect 1209 13698 1275 13701
rect 62 13696 1275 13698
rect 62 13640 1214 13696
rect 1270 13640 1275 13696
rect 62 13638 1275 13640
rect 1209 13635 1275 13638
rect 13813 13698 13879 13701
rect 15929 13698 15995 13701
rect 13813 13696 15995 13698
rect 13813 13640 13818 13696
rect 13874 13640 15934 13696
rect 15990 13640 15995 13696
rect 13813 13638 15995 13640
rect 13813 13635 13879 13638
rect 15929 13635 15995 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3601 13562 3667 13565
rect 3601 13560 4170 13562
rect 3601 13504 3606 13560
rect 3662 13504 4170 13560
rect 3601 13502 4170 13504
rect 3601 13499 3667 13502
rect 4110 13426 4170 13502
rect 14273 13426 14339 13429
rect 4110 13424 14339 13426
rect 4110 13368 14278 13424
rect 14334 13368 14339 13424
rect 4110 13366 14339 13368
rect 14273 13363 14339 13366
rect 14641 13426 14707 13429
rect 20253 13426 20319 13429
rect 14641 13424 20319 13426
rect 14641 13368 14646 13424
rect 14702 13368 20258 13424
rect 20314 13368 20319 13424
rect 14641 13366 20319 13368
rect 14641 13363 14707 13366
rect 20253 13363 20319 13366
rect 3877 13290 3943 13293
rect 23841 13290 23907 13293
rect 3877 13288 23907 13290
rect 3877 13232 3882 13288
rect 3938 13232 23846 13288
rect 23902 13232 23907 13288
rect 3877 13230 23907 13232
rect 3877 13227 3943 13230
rect 23841 13227 23907 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 2129 13018 2195 13021
rect 62 13016 4170 13018
rect 62 12960 2134 13016
rect 2190 12960 4170 13016
rect 62 12958 4170 12960
rect 62 12504 122 12958
rect 2129 12955 2195 12958
rect 4110 12882 4170 12958
rect 27520 12928 28000 13048
rect 14641 12882 14707 12885
rect 21173 12882 21239 12885
rect 4110 12880 14707 12882
rect 4110 12824 14646 12880
rect 14702 12824 14707 12880
rect 4110 12822 14707 12824
rect 14641 12819 14707 12822
rect 14782 12880 21239 12882
rect 14782 12824 21178 12880
rect 21234 12824 21239 12880
rect 14782 12822 21239 12824
rect 10961 12746 11027 12749
rect 14782 12746 14842 12822
rect 21173 12819 21239 12822
rect 10961 12744 14842 12746
rect 10961 12688 10966 12744
rect 11022 12688 14842 12744
rect 10961 12686 14842 12688
rect 17769 12746 17835 12749
rect 20069 12746 20135 12749
rect 17769 12744 20135 12746
rect 17769 12688 17774 12744
rect 17830 12688 20074 12744
rect 20130 12688 20135 12744
rect 17769 12686 20135 12688
rect 10961 12683 11027 12686
rect 17769 12683 17835 12686
rect 20069 12683 20135 12686
rect 10277 12544 10597 12545
rect 0 12384 480 12504
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 24761 12474 24827 12477
rect 27662 12474 27722 12928
rect 24761 12472 27722 12474
rect 24761 12416 24766 12472
rect 24822 12416 27722 12472
rect 24761 12414 27722 12416
rect 24761 12411 24827 12414
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 7557 11794 7623 11797
rect 23841 11794 23907 11797
rect 7557 11792 23907 11794
rect 7557 11736 7562 11792
rect 7618 11736 23846 11792
rect 23902 11736 23907 11792
rect 7557 11734 23907 11736
rect 7557 11731 7623 11734
rect 23841 11731 23907 11734
rect 12525 11658 12591 11661
rect 18873 11658 18939 11661
rect 12525 11656 18939 11658
rect 12525 11600 12530 11656
rect 12586 11600 18878 11656
rect 18934 11600 18939 11656
rect 12525 11598 18939 11600
rect 12525 11595 12591 11598
rect 18873 11595 18939 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 54 11188 60 11252
rect 124 11250 130 11252
rect 24761 11250 24827 11253
rect 27654 11250 27660 11252
rect 124 11190 4768 11250
rect 124 11188 130 11190
rect 4708 11117 4768 11190
rect 24761 11248 27660 11250
rect 24761 11192 24766 11248
rect 24822 11192 27660 11248
rect 24761 11190 27660 11192
rect 24761 11187 24827 11190
rect 27654 11188 27660 11190
rect 27724 11188 27730 11252
rect 4705 11114 4771 11117
rect 13721 11114 13787 11117
rect 4705 11112 13787 11114
rect 4705 11056 4710 11112
rect 4766 11056 13726 11112
rect 13782 11056 13787 11112
rect 4705 11054 13787 11056
rect 4705 11051 4771 11054
rect 13721 11051 13787 11054
rect 0 10980 480 11008
rect 0 10916 60 10980
rect 124 10916 480 10980
rect 0 10888 480 10916
rect 27520 10980 28000 11008
rect 27520 10916 27660 10980
rect 27724 10916 28000 10980
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 27520 10888 28000 10916
rect 24277 10847 24597 10848
rect 9029 10706 9095 10709
rect 14549 10706 14615 10709
rect 9029 10704 14615 10706
rect 9029 10648 9034 10704
rect 9090 10648 14554 10704
rect 14610 10648 14615 10704
rect 9029 10646 14615 10648
rect 9029 10643 9095 10646
rect 14549 10643 14615 10646
rect 6545 10570 6611 10573
rect 16757 10570 16823 10573
rect 18965 10570 19031 10573
rect 6545 10568 19031 10570
rect 6545 10512 6550 10568
rect 6606 10512 16762 10568
rect 16818 10512 18970 10568
rect 19026 10512 19031 10568
rect 6545 10510 19031 10512
rect 6545 10507 6611 10510
rect 16757 10507 16823 10510
rect 18965 10507 19031 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 2681 10162 2747 10165
rect 62 10160 2747 10162
rect 62 10104 2686 10160
rect 2742 10104 2747 10160
rect 62 10102 2747 10104
rect 62 9648 122 10102
rect 2681 10099 2747 10102
rect 7465 10162 7531 10165
rect 19425 10162 19491 10165
rect 7465 10160 19491 10162
rect 7465 10104 7470 10160
rect 7526 10104 19430 10160
rect 19486 10104 19491 10160
rect 7465 10102 19491 10104
rect 7465 10099 7531 10102
rect 19425 10099 19491 10102
rect 11145 10026 11211 10029
rect 11881 10026 11947 10029
rect 21449 10026 21515 10029
rect 11145 10024 21515 10026
rect 11145 9968 11150 10024
rect 11206 9968 11886 10024
rect 11942 9968 21454 10024
rect 21510 9968 21515 10024
rect 11145 9966 21515 9968
rect 11145 9963 11211 9966
rect 11881 9963 11947 9966
rect 21449 9963 21515 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 0 9528 480 9648
rect 19241 9618 19307 9621
rect 20161 9618 20227 9621
rect 27654 9618 27660 9620
rect 19241 9616 27660 9618
rect 19241 9560 19246 9616
rect 19302 9560 20166 9616
rect 20222 9560 27660 9616
rect 19241 9558 27660 9560
rect 19241 9555 19307 9558
rect 20161 9555 20227 9558
rect 27654 9556 27660 9558
rect 27724 9556 27730 9620
rect 2037 9346 2103 9349
rect 7741 9346 7807 9349
rect 2037 9344 7807 9346
rect 2037 9288 2042 9344
rect 2098 9288 7746 9344
rect 7802 9288 7807 9344
rect 2037 9286 7807 9288
rect 2037 9283 2103 9286
rect 7741 9283 7807 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 4153 9210 4219 9213
rect 8201 9210 8267 9213
rect 4153 9208 8267 9210
rect 4153 9152 4158 9208
rect 4214 9152 8206 9208
rect 8262 9152 8267 9208
rect 4153 9150 8267 9152
rect 4153 9147 4219 9150
rect 8201 9147 8267 9150
rect 27520 8848 28000 8968
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 17861 8530 17927 8533
rect 27662 8530 27722 8848
rect 17861 8528 27722 8530
rect 17861 8472 17866 8528
rect 17922 8472 27722 8528
rect 17861 8470 27722 8472
rect 17861 8467 17927 8470
rect 10277 8192 10597 8193
rect 0 8032 480 8152
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 62 7578 122 8032
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 1853 7578 1919 7581
rect 62 7576 1919 7578
rect 62 7520 1858 7576
rect 1914 7520 1919 7576
rect 62 7518 1919 7520
rect 1853 7515 1919 7518
rect 18781 7442 18847 7445
rect 27705 7442 27771 7445
rect 18781 7440 27771 7442
rect 18781 7384 18786 7440
rect 18842 7384 27710 7440
rect 27766 7384 27771 7440
rect 18781 7382 27771 7384
rect 18781 7379 18847 7382
rect 27705 7379 27771 7382
rect 14273 7306 14339 7309
rect 17585 7306 17651 7309
rect 27613 7306 27679 7309
rect 14273 7304 27679 7306
rect 14273 7248 14278 7304
rect 14334 7248 17590 7304
rect 17646 7248 27618 7304
rect 27674 7248 27679 7304
rect 14273 7246 27679 7248
rect 14273 7243 14339 7246
rect 17585 7243 17651 7246
rect 27613 7243 27679 7246
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 25497 7034 25563 7037
rect 27520 7034 28000 7064
rect 25497 7032 28000 7034
rect 25497 6976 25502 7032
rect 25558 6976 28000 7032
rect 25497 6974 28000 6976
rect 25497 6971 25563 6974
rect 27520 6944 28000 6974
rect 0 6624 480 6656
rect 0 6568 110 6624
rect 166 6568 480 6624
rect 0 6536 480 6568
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 7741 6218 7807 6221
rect 15653 6218 15719 6221
rect 7741 6216 15719 6218
rect 7741 6160 7746 6216
rect 7802 6160 15658 6216
rect 15714 6160 15719 6216
rect 7741 6158 15719 6160
rect 7741 6155 7807 6158
rect 15653 6155 15719 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 1301 5674 1367 5677
rect 62 5672 1367 5674
rect 62 5616 1306 5672
rect 1362 5616 1367 5672
rect 62 5614 1367 5616
rect 62 5160 122 5614
rect 1301 5611 1367 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 0 5040 480 5160
rect 27520 4992 28000 5024
rect 27520 4936 27618 4992
rect 27674 4936 28000 4992
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 27520 4904 28000 4936
rect 19610 4863 19930 4864
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 5073 4178 5139 4181
rect 62 4176 5139 4178
rect 62 4120 5078 4176
rect 5134 4120 5139 4176
rect 62 4118 5139 4120
rect 62 3664 122 4118
rect 5073 4115 5139 4118
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 0 3544 480 3664
rect 8661 3362 8727 3365
rect 13813 3362 13879 3365
rect 8661 3360 13879 3362
rect 8661 3304 8666 3360
rect 8722 3304 13818 3360
rect 13874 3304 13879 3360
rect 8661 3302 13879 3304
rect 8661 3299 8727 3302
rect 13813 3299 13879 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 27520 2956 28000 2984
rect 27520 2892 27660 2956
rect 27724 2892 28000 2956
rect 27520 2864 28000 2892
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 5533 2682 5599 2685
rect 62 2680 5599 2682
rect 62 2624 5538 2680
rect 5594 2624 5599 2680
rect 62 2622 5599 2624
rect 62 2168 122 2622
rect 5533 2619 5599 2622
rect 13169 2410 13235 2413
rect 20621 2410 20687 2413
rect 13169 2408 20687 2410
rect 13169 2352 13174 2408
rect 13230 2352 20626 2408
rect 20682 2352 20687 2408
rect 13169 2350 20687 2352
rect 13169 2347 13235 2350
rect 20621 2347 20687 2350
rect 5610 2208 5930 2209
rect 0 2048 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 4521 1322 4587 1325
rect 62 1320 4587 1322
rect 62 1264 4526 1320
rect 4582 1264 4587 1320
rect 62 1262 4587 1264
rect 62 808 122 1262
rect 4521 1259 4587 1262
rect 27520 1048 28000 1080
rect 27520 992 27710 1048
rect 27766 992 28000 1048
rect 27520 960 28000 992
rect 0 688 480 808
rect 8109 98 8175 101
rect 18689 98 18755 101
rect 8109 96 18755 98
rect 8109 40 8114 96
rect 8170 40 18694 96
rect 18750 40 18755 96
rect 8109 38 18755 40
rect 8109 35 8175 38
rect 18689 35 18755 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 60 16900 124 16964
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 60 16628 124 16692
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 60 11188 124 11252
rect 27660 11188 27724 11252
rect 60 10916 124 10980
rect 27660 10916 27724 10980
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 27660 9556 27724 9620
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 27660 2892 27724 2956
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 59 16964 125 16965
rect 59 16900 60 16964
rect 124 16900 125 16964
rect 59 16899 125 16900
rect 62 16693 122 16899
rect 59 16692 125 16693
rect 59 16628 60 16692
rect 124 16628 125 16692
rect 59 16627 125 16628
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 59 11252 125 11253
rect 59 11188 60 11252
rect 124 11188 125 11252
rect 59 11187 125 11188
rect 62 10981 122 11187
rect 59 10980 125 10981
rect 59 10916 60 10980
rect 124 10916 125 10980
rect 59 10915 125 10916
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 27659 11252 27725 11253
rect 27659 11188 27660 11252
rect 27724 11188 27725 11252
rect 27659 11187 27725 11188
rect 27662 10981 27722 11187
rect 27659 10980 27725 10981
rect 27659 10916 27660 10980
rect 27724 10916 27725 10980
rect 27659 10915 27725 10916
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 27659 9620 27725 9621
rect 27659 9556 27660 9620
rect 27724 9556 27725 9620
rect 27659 9555 27725 9556
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 27662 2957 27722 9555
rect 27659 2956 27725 2957
rect 27659 2892 27660 2956
rect 27724 2892 27725 2956
rect 27659 2891 27725 2892
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_38 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_42
timestamp 1586364061
transform 1 0 4968 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_49
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_53 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5980 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_1_51
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_61 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_59
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _205_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_87 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 774 592
use scs8hd_decap_4  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 406 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_104
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_92
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_95
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_108
timestamp 1586364061
transform 1 0 11040 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 774 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _214_
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_128
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_132
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_142
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _212_
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__214__A
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_154
timestamp 1586364061
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _211_
timestamp 1586364061
transform 1 0 16836 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__212__A
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__211__A
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_163
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_167
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_175
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_179
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_185
timestamp 1586364061
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_195
timestamp 1586364061
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_204
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_239
timestamp 1586364061
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_234
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _221_
timestamp 1586364061
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_243
timestamp 1586364061
transform 1 0 23460 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__221__A
timestamp 1586364061
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_275
timestamp 1586364061
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_8  _177_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_91
timestamp 1586364061
transform 1 0 9476 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_118
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_130
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_150
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_3_83
timestamp 1586364061
transform 1 0 8740 0 1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_92
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_96
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_204
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_210
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_214
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_226
timestamp 1586364061
transform 1 0 21896 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_238
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_76
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_8  _178_
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_12  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_133
timestamp 1586364061
transform 1 0 13340 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_251
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_263
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  FILLER_5_70
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_109
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_128
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_140
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_152
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_164
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_5_176
timestamp 1586364061
transform 1 0 17296 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_182
timestamp 1586364061
transform 1 0 17848 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_19
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__077__C
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_70
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 130 592
use scs8hd_buf_1  _128_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_73
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_77
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_96
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_107
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_113
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_109
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _195_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_121
timestamp 1586364061
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_117
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_6_118
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_128
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__217__A
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _217_
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13708 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_139
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_133
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_163
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_18
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use scs8hd_or3_4  _077_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_40
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_8_70
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 314 592
use scs8hd_nor2_4  _129_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 10120 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_97
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_101
timestamp 1586364061
transform 1 0 10396 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11132 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_118
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 314 592
use scs8hd_inv_8  _075_
timestamp 1586364061
transform 1 0 5060 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_52
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_56
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_60
timestamp 1586364061
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_65
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_69
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_111
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_115
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_126
timestamp 1586364061
transform 1 0 12696 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_130
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_137
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_141
timestamp 1586364061
transform 1 0 14076 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_144
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_152
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_160
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_172
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 866 592
use scs8hd_buf_1  _158_
timestamp 1586364061
transform 1 0 4508 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_40
timestamp 1586364061
transform 1 0 4784 0 -1 8160
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__C
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_61
timestamp 1586364061
transform 1 0 6716 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_72
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_88
timestamp 1586364061
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_108
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_112
timestamp 1586364061
transform 1 0 11408 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_120
timestamp 1586364061
transform 1 0 12144 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_134
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_138
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_163
timestamp 1586364061
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_173
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_176
timestamp 1586364061
transform 1 0 17296 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_188
timestamp 1586364061
transform 1 0 18400 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_200
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_10_212
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _078_
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_22
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_26
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_35
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 5060 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_52
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use scs8hd_or3_4  _096_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__093__C
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_56
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_91
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_99
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_111
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_115
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_119
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_134
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_172
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_176
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_187
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_205
timestamp 1586364061
transform 1 0 19964 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_229
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_11_241
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__081__C
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_12
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_16
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _156_
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_29
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_8  _076_
timestamp 1586364061
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 5520 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_46
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_50
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use scs8hd_or3_4  _093_
timestamp 1586364061
transform 1 0 6072 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_63
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 590 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_2  FILLER_12_104
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_138
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_142
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_146
timestamp 1586364061
transform 1 0 14536 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_150
timestamp 1586364061
transform 1 0 14904 0 -1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_167
timestamp 1586364061
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_171
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_183
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_187
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_16
timestamp 1586364061
transform 1 0 2576 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_12
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_inv_8  _114_
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 866 592
use scs8hd_or3_4  _081_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_24
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_20
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _136_
timestamp 1586364061
transform 1 0 2944 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_35
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_39
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_40
timestamp 1586364061
transform 1 0 4784 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_36
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_52
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_or3_4  _099_
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 866 592
use scs8hd_or3_4  _090_
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 6624 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_67
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_63
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_65
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_buf_1  _097_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_69
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_89
timestamp 1586364061
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_85
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1050 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_104
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_114
timestamp 1586364061
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_110
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_112
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_108
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_120
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_116
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_127
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_135
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_149
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_155
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_172
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_172
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_175
timestamp 1586364061
transform 1 0 17204 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_194
timestamp 1586364061
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_187
timestamp 1586364061
transform 1 0 18308 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_198
timestamp 1586364061
transform 1 0 19320 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_210
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_198
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_210
timestamp 1586364061
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_13_222
timestamp 1586364061
transform 1 0 21528 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_234
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_242
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_or3_4  _104_
timestamp 1586364061
transform 1 0 1472 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_13
timestamp 1586364061
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_17
timestamp 1586364061
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_21
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_25
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _185_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_78
timestamp 1586364061
transform 1 0 8280 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _181_
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_94
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_102
timestamp 1586364061
transform 1 0 10488 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14904 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_146
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_163
timestamp 1586364061
transform 1 0 16100 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_169
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_204
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_222
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_234
timestamp 1586364061
transform 1 0 22632 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_242
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 24564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_253
timestamp 1586364061
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_inv_8  _103_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_12
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_16
timestamp 1586364061
transform 1 0 2576 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 2944 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_35
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__172__C
timestamp 1586364061
transform 1 0 4508 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_39
timestamp 1586364061
transform 1 0 4692 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__C
timestamp 1586364061
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_54
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_58
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_75
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_78
timestamp 1586364061
transform 1 0 8280 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_109
timestamp 1586364061
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_122
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_126
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_130
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_149
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_165
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_169
timestamp 1586364061
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_182
timestamp 1586364061
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_203
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  FILLER_16_211
timestamp 1586364061
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_2  _223_
timestamp 1586364061
transform 1 0 21344 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_219
timestamp 1586364061
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_236
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_16_248
timestamp 1586364061
transform 1 0 23920 0 -1 11424
box -38 -48 590 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_254
timestamp 1586364061
transform 1 0 24472 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_259
timestamp 1586364061
transform 1 0 24932 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_271
timestamp 1586364061
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_14.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2668 0 1 11424
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_6
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_10
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_14
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__172__D
timestamp 1586364061
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_28
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_34
timestamp 1586364061
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _171_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4416 0 1 11424
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _116_
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__164__C
timestamp 1586364061
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__B
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_65
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_69
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _167_
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 1602 592
use scs8hd_decap_3  FILLER_17_73
timestamp 1586364061
transform 1 0 7820 0 1 11424
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_97
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_137
timestamp 1586364061
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_141
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_160
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_163
timestamp 1586364061
transform 1 0 16100 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_199
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_204
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_215
timestamp 1586364061
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_219
timestamp 1586364061
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_223
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_235
timestamp 1586364061
transform 1 0 22724 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_243
timestamp 1586364061
transform 1 0 23460 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_249
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 590 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_259
timestamp 1586364061
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_263
timestamp 1586364061
transform 1 0 25300 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_275
timestamp 1586364061
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _082_
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_8  _186_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _172_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_49
timestamp 1586364061
transform 1 0 5612 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_53
timestamp 1586364061
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _164_
timestamp 1586364061
transform 1 0 7268 0 -1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__164__D
timestamp 1586364061
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__D
timestamp 1586364061
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_57
timestamp 1586364061
transform 1 0 6348 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_63
timestamp 1586364061
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _163_
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__167__D
timestamp 1586364061
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_114
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_8  _182_
timestamp 1586364061
transform 1 0 13524 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_127
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_131
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_144
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_148
timestamp 1586364061
transform 1 0 14720 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_151
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_160
timestamp 1586364061
transform 1 0 15824 0 -1 12512
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15916 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_172
timestamp 1586364061
transform 1 0 16928 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_176
timestamp 1586364061
transform 1 0 17296 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17664 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_189
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_193
timestamp 1586364061
transform 1 0 18860 0 -1 12512
box -38 -48 406 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_218
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_230
timestamp 1586364061
transform 1 0 22264 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_242
timestamp 1586364061
transform 1 0 23368 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_247
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_259
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_271
timestamp 1586364061
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_17
timestamp 1586364061
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_13
timestamp 1586364061
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_12
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 -1 13600
box -38 -48 866 592
use scs8hd_or3_4  _115_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_20_25
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_21
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_33
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_29
timestamp 1586364061
transform 1 0 3772 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _179_
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__D
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_49
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_45
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_50
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_46
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__C
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 222 592
use scs8hd_or3_4  _135_
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_conb_1  _192_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_64
timestamp 1586364061
transform 1 0 6992 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_69
timestamp 1586364061
transform 1 0 7452 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_65
timestamp 1586364061
transform 1 0 7084 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 7544 0 1 12512
box -38 -48 222 592
use scs8hd_or3_4  _137_
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 866 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use scs8hd_nor4_4  _168_
timestamp 1586364061
transform 1 0 8096 0 1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__D
timestamp 1586364061
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_72
timestamp 1586364061
transform 1 0 7728 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_88
timestamp 1586364061
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_97
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_93
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_104
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__C
timestamp 1586364061
transform 1 0 10212 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10396 0 -1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_12.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_20_108
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_116
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_140
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_138
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_1  FILLER_20_150
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_146
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_145
timestamp 1586364061
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_158
timestamp 1586364061
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_167
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_162
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_171
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_183
timestamp 1586364061
transform 1 0 17940 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_179
timestamp 1586364061
transform 1 0 17572 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_196
timestamp 1586364061
transform 1 0 19136 0 -1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_204
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_208
timestamp 1586364061
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_215
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_219
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_223
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_235
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_19_243
timestamp 1586364061
transform 1 0 23460 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_249
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_247
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_261
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_273
timestamp 1586364061
transform 1 0 26220 0 1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_14
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3128 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_18
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 130 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 314 592
use scs8hd_buf_1  _126_
timestamp 1586364061
transform 1 0 5704 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__C
timestamp 1586364061
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_38
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_42
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_46
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 6900 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 7360 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__D
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_70
timestamp 1586364061
transform 1 0 7544 0 1 13600
box -38 -48 222 592
use scs8hd_nor4_4  _169_
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use scs8hd_or3_4  _117_
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_91
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_108
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_116
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_138
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_142
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_153
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_157
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_170
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_21_176
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_180
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20608 0 1 13600
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_204
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_215
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_219
timestamp 1586364061
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_223
timestamp 1586364061
transform 1 0 21620 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_235
timestamp 1586364061
transform 1 0 22724 0 1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_21_243
timestamp 1586364061
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__210__A
timestamp 1586364061
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_253
timestamp 1586364061
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_258
timestamp 1586364061
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_262
timestamp 1586364061
transform 1 0 25208 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_266
timestamp 1586364061
transform 1 0 25576 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_274
timestamp 1586364061
transform 1 0 26312 0 1 13600
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1472 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_22_24
timestamp 1586364061
transform 1 0 3312 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_28
timestamp 1586364061
transform 1 0 3680 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use scs8hd_nor4_4  _165_
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_22_53
timestamp 1586364061
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_8  _125_
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__C
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_57
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 406 592
use scs8hd_conb_1  _196_
timestamp 1586364061
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_76
timestamp 1586364061
transform 1 0 8096 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 10120 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_96
timestamp 1586364061
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_100
timestamp 1586364061
transform 1 0 10304 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_115
timestamp 1586364061
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_119
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_132
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_136
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_143
timestamp 1586364061
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_147
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_165
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_169
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_173
timestamp 1586364061
transform 1 0 17020 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_200
timestamp 1586364061
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_204
timestamp 1586364061
transform 1 0 19872 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_22_212
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_218
timestamp 1586364061
transform 1 0 21160 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_230
timestamp 1586364061
transform 1 0 22264 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_242
timestamp 1586364061
transform 1 0 23368 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_2  _210_
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_254
timestamp 1586364061
transform 1 0 24472 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_259
timestamp 1586364061
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_271
timestamp 1586364061
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_conb_1  _190_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_10.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 1050 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_6
timestamp 1586364061
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_10
timestamp 1586364061
transform 1 0 2024 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_14
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_28
timestamp 1586364061
transform 1 0 3680 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_34
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use scs8hd_nor4_4  _166_
timestamp 1586364061
transform 1 0 4416 0 1 14688
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _079_
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__B
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_65
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_69
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 130 592
use scs8hd_nor4_4  _170_
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_23_72
timestamp 1586364061
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_23_119
timestamp 1586364061
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_142
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 14444 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_158
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_173
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_210
timestamp 1586364061
transform 1 0 20424 0 1 14688
box -38 -48 774 592
use scs8hd_buf_1  _118_
timestamp 1586364061
transform 1 0 21160 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_221
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_225
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_23_237
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_23_243
timestamp 1586364061
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_19
timestamp 1586364061
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use scs8hd_or3_4  _146_
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_45
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_49
timestamp 1586364061
transform 1 0 5612 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__D
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__C
timestamp 1586364061
transform 1 0 9292 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_79
timestamp 1586364061
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_87
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use scs8hd_or3_4  _106_
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_110
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_115
timestamp 1586364061
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _184_
timestamp 1586364061
transform 1 0 13432 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_130
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 15824 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_143
timestamp 1586364061
transform 1 0 14260 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_171
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_179
timestamp 1586364061
transform 1 0 17572 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_191
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_195
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _198_
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_218
timestamp 1586364061
transform 1 0 21160 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_230
timestamp 1586364061
transform 1 0 22264 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_242
timestamp 1586364061
transform 1 0 23368 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_254
timestamp 1586364061
transform 1 0 24472 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_24_266
timestamp 1586364061
transform 1 0 25576 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_274
timestamp 1586364061
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__159__D
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_14
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_nor4_4  _159_
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__C
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_18
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_52
timestamp 1586364061
transform 1 0 5888 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_67
timestamp 1586364061
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_nor4_4  _162_
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_96
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _183_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_117
timestamp 1586364061
transform 1 0 11868 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_140
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 130 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_152
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_156
timestamp 1586364061
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_194
timestamp 1586364061
transform 1 0 18952 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19688 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_198
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_211
timestamp 1586364061
transform 1 0 20516 0 1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_228
timestamp 1586364061
transform 1 0 22080 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_253
timestamp 1586364061
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_7
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_2  _216_
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_16
timestamp 1586364061
transform 1 0 2576 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_12
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__216__A
timestamp 1586364061
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use scs8hd_inv_8  _180_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_26
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_22
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__D
timestamp 1586364061
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_1  _160_
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 1050 592
use scs8hd_nor4_4  _157_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1602 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5520 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_49
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_41
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_45
timestamp 1586364061
transform 1 0 5244 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_61
timestamp 1586364061
transform 1 0 6716 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_69
timestamp 1586364061
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_65
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 6900 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_77
timestamp 1586364061
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__D
timestamp 1586364061
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_buf_1  _107_
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 314 592
use scs8hd_nor4_4  _161_
timestamp 1586364061
transform 1 0 8004 0 1 16864
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_27_96
timestamp 1586364061
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_92
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10304 0 1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9752 0 -1 16864
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_27_115
timestamp 1586364061
transform 1 0 11684 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_111
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_109
timestamp 1586364061
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_119
timestamp 1586364061
transform 1 0 12052 0 1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_122
timestamp 1586364061
transform 1 0 12328 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_8  _176_
timestamp 1586364061
transform 1 0 13064 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_139
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_140
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_155
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_157
timestamp 1586364061
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_161
timestamp 1586364061
transform 1 0 15916 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_165
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_177
timestamp 1586364061
transform 1 0 17388 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_27_178
timestamp 1586364061
transform 1 0 17480 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_181
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_181
timestamp 1586364061
transform 1 0 17756 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17940 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_194
timestamp 1586364061
transform 1 0 18952 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_194
timestamp 1586364061
transform 1 0 18952 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 16864
box -38 -48 866 592
use scs8hd_fill_1  FILLER_27_202
timestamp 1586364061
transform 1 0 19688 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_198
timestamp 1586364061
transform 1 0 19320 0 1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_26_204
timestamp 1586364061
transform 1 0 19872 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_206
timestamp 1586364061
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_212
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_210
timestamp 1586364061
transform 1 0 20424 0 1 16864
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_221
timestamp 1586364061
transform 1 0 21436 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_222
timestamp 1586364061
transform 1 0 21528 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_233
timestamp 1586364061
transform 1 0 22540 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_26_245
timestamp 1586364061
transform 1 0 23644 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_27_234
timestamp 1586364061
transform 1 0 22632 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_242
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_253
timestamp 1586364061
transform 1 0 24380 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_258
timestamp 1586364061
transform 1 0 24840 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_253
timestamp 1586364061
transform 1 0 24380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_259
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_263
timestamp 1586364061
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_270
timestamp 1586364061
transform 1 0 25944 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_275
timestamp 1586364061
transform 1 0 26404 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _154_
timestamp 1586364061
transform 1 0 1932 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_12
timestamp 1586364061
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_16
timestamp 1586364061
transform 1 0 2576 0 -1 17952
box -38 -48 406 592
use scs8hd_buf_1  _155_
timestamp 1586364061
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 17952
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_track_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_36
timestamp 1586364061
transform 1 0 4416 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_40
timestamp 1586364061
transform 1 0 4784 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_46
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__161__C
timestamp 1586364061
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_59
timestamp 1586364061
transform 1 0 6532 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_79
timestamp 1586364061
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_83
timestamp 1586364061
transform 1 0 8740 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_87
timestamp 1586364061
transform 1 0 9108 0 -1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_90
timestamp 1586364061
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_102
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_106
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_121
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_138
timestamp 1586364061
transform 1 0 13800 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_148
timestamp 1586364061
transform 1 0 14720 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_171
timestamp 1586364061
transform 1 0 16836 0 -1 17952
box -38 -48 590 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19136 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_188
timestamp 1586364061
transform 1 0 18400 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_192
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_199
timestamp 1586364061
transform 1 0 19412 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_203
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_211
timestamp 1586364061
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_1  _147_
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_6
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_10
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_17
timestamp 1586364061
transform 1 0 2668 0 1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3404 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_22
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_36
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_40
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_84
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use scs8hd_inv_8  _175_
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_132
timestamp 1586364061
transform 1 0 13248 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_138
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_142
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 406 592
use scs8hd_conb_1  _194_
timestamp 1586364061
transform 1 0 16468 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_163
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_29_166
timestamp 1586364061
transform 1 0 16376 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_210
timestamp 1586364061
transform 1 0 20424 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_222
timestamp 1586364061
transform 1 0 21528 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_29_234
timestamp 1586364061
transform 1 0 22632 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_242
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_10.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_8  _173_
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_18
timestamp 1586364061
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_41
timestamp 1586364061
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_46
timestamp 1586364061
transform 1 0 5336 0 -1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_60
timestamp 1586364061
transform 1 0 6624 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_64
timestamp 1586364061
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_77
timestamp 1586364061
transform 1 0 8188 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_81
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_85
timestamp 1586364061
transform 1 0 8924 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_89
timestamp 1586364061
transform 1 0 9292 0 -1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11500 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_110
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_122
timestamp 1586364061
transform 1 0 12328 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_128
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_150
timestamp 1586364061
transform 1 0 14904 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_159
timestamp 1586364061
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16192 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16008 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_175
timestamp 1586364061
transform 1 0 17204 0 -1 19040
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17940 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18952 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_192
timestamp 1586364061
transform 1 0 18768 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_196
timestamp 1586364061
transform 1 0 19136 0 -1 19040
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19504 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_203
timestamp 1586364061
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_30_207
timestamp 1586364061
transform 1 0 20148 0 -1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_30_213
timestamp 1586364061
transform 1 0 20700 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_11
timestamp 1586364061
transform 1 0 2116 0 1 19040
box -38 -48 314 592
use scs8hd_decap_4  FILLER_31_16
timestamp 1586364061
transform 1 0 2576 0 1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3496 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3312 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_22
timestamp 1586364061
transform 1 0 3128 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_35
timestamp 1586364061
transform 1 0 4324 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_53
timestamp 1586364061
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_71
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8372 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_75
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_88
timestamp 1586364061
transform 1 0 9200 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_92
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_105
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_109
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_113
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 314 592
use scs8hd_nor2_4  _098_
timestamp 1586364061
transform 1 0 13892 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 13708 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 13340 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_131
timestamp 1586364061
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15548 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_148
timestamp 1586364061
transform 1 0 14720 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_154
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_168
timestamp 1586364061
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_172
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_176
timestamp 1586364061
transform 1 0 17296 0 1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_195
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_199
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_212
timestamp 1586364061
transform 1 0 20608 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_224
timestamp 1586364061
transform 1 0 21712 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_31_236
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_inv_8  _174_
timestamp 1586364061
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  FILLER_32_11
timestamp 1586364061
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_23
timestamp 1586364061
transform 1 0 3220 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 130 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 5796 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_42
timestamp 1586364061
transform 1 0 4968 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_50
timestamp 1586364061
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_60
timestamp 1586364061
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 -1 20128
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10948 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_97
timestamp 1586364061
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_101
timestamp 1586364061
transform 1 0 10396 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_116
timestamp 1586364061
transform 1 0 11776 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_124
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_137
timestamp 1586364061
transform 1 0 13708 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16008 0 -1 20128
box -38 -48 1050 592
use scs8hd_decap_12  FILLER_32_173
timestamp 1586364061
transform 1 0 17020 0 -1 20128
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_194
timestamp 1586364061
transform 1 0 18952 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_198
timestamp 1586364061
transform 1 0 19320 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_32_205
timestamp 1586364061
transform 1 0 19964 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_209
timestamp 1586364061
transform 1 0 20332 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_conb_1  _197_
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_218
timestamp 1586364061
transform 1 0 21160 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_230
timestamp 1586364061
transform 1 0 22264 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_242
timestamp 1586364061
transform 1 0 23368 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_254
timestamp 1586364061
transform 1 0 24472 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_266
timestamp 1586364061
transform 1 0 25576 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_274
timestamp 1586364061
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_buf_2  _219_
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__219__A
timestamp 1586364061
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2576 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_7
timestamp 1586364061
transform 1 0 1748 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_23
timestamp 1586364061
transform 1 0 3220 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_19
timestamp 1586364061
transform 1 0 2852 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_18
timestamp 1586364061
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use scs8hd_conb_1  _193_
timestamp 1586364061
transform 1 0 2944 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_35
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_31
timestamp 1586364061
transform 1 0 3956 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3128 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 5980 0 -1 21216
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_48
timestamp 1586364061
transform 1 0 5520 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_52
timestamp 1586364061
transform 1 0 5888 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_41
timestamp 1586364061
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_45
timestamp 1586364061
transform 1 0 5244 0 -1 21216
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_55
timestamp 1586364061
transform 1 0 6164 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_64
timestamp 1586364061
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_76
timestamp 1586364061
transform 1 0 8096 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_72
timestamp 1586364061
transform 1 0 7728 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_86
timestamp 1586364061
transform 1 0 9016 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_34_82
timestamp 1586364061
transform 1 0 8648 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_89
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7820 0 -1 21216
box -38 -48 866 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 8464 0 1 20128
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_96
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_95
timestamp 1586364061
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_101
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10212 0 -1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10212 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10948 0 -1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_114
timestamp 1586364061
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_118
timestamp 1586364061
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_118
timestamp 1586364061
transform 1 0 11960 0 -1 21216
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 21216
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12880 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14076 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_139
timestamp 1586364061
transform 1 0 13892 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_126
timestamp 1586364061
transform 1 0 12696 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_33_143
timestamp 1586364061
transform 1 0 14260 0 1 20128
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_34_151
timestamp 1586364061
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_150
timestamp 1586364061
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15088 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 15456 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_34_158
timestamp 1586364061
transform 1 0 15640 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16100 0 1 20128
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15916 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_174
timestamp 1586364061
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_178
timestamp 1586364061
transform 1 0 17480 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_174
timestamp 1586364061
transform 1 0 17112 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_186
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_34_181
timestamp 1586364061
transform 1 0 17756 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17572 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_193
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_197
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_210
timestamp 1586364061
transform 1 0 20424 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_34_200
timestamp 1586364061
transform 1 0 19504 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_204
timestamp 1586364061
transform 1 0 19872 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_34_212
timestamp 1586364061
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_222
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_234
timestamp 1586364061
transform 1 0 22632 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_242
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_258
timestamp 1586364061
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_262
timestamp 1586364061
transform 1 0 25208 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_274
timestamp 1586364061
transform 1 0 26312 0 1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2024 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_9
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_12
timestamp 1586364061
transform 1 0 2208 0 1 21216
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_35_24
timestamp 1586364061
transform 1 0 3312 0 1 21216
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5704 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_43
timestamp 1586364061
transform 1 0 5060 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_47
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_52
timestamp 1586364061
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_73
timestamp 1586364061
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_77
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10212 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_90
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_95
timestamp 1586364061
transform 1 0 9844 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12972 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_127
timestamp 1586364061
transform 1 0 12788 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_140
timestamp 1586364061
transform 1 0 13984 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_144
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_158
timestamp 1586364061
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_162
timestamp 1586364061
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_193
timestamp 1586364061
transform 1 0 18860 0 1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_198
timestamp 1586364061
transform 1 0 19320 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_204
timestamp 1586364061
transform 1 0 19872 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_35_248
timestamp 1586364061
transform 1 0 23920 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_252
timestamp 1586364061
transform 1 0 24288 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_264
timestamp 1586364061
transform 1 0 25392 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_fill_1  FILLER_35_276
timestamp 1586364061
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2024 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_9
timestamp 1586364061
transform 1 0 1932 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_13
timestamp 1586364061
transform 1 0 2300 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_25
timestamp 1586364061
transform 1 0 3404 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_6  FILLER_36_36
timestamp 1586364061
transform 1 0 4416 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_42
timestamp 1586364061
transform 1 0 4968 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_46
timestamp 1586364061
transform 1 0 5336 0 -1 22304
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6072 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_57
timestamp 1586364061
transform 1 0 6348 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_61
timestamp 1586364061
transform 1 0 6716 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_64
timestamp 1586364061
transform 1 0 6992 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 8648 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_74
timestamp 1586364061
transform 1 0 7912 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_8  FILLER_36_84
timestamp 1586364061
transform 1 0 8832 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 590 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 11776 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_36_108
timestamp 1586364061
transform 1 0 11040 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13340 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13156 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_125
timestamp 1586364061
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_142
timestamp 1586364061
transform 1 0 14168 0 -1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_146
timestamp 1586364061
transform 1 0 14536 0 -1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_36_152
timestamp 1586364061
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_163
timestamp 1586364061
transform 1 0 16100 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_168
timestamp 1586364061
transform 1 0 16560 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_36_176
timestamp 1586364061
transform 1 0 17296 0 -1 22304
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17572 0 -1 22304
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19136 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_188
timestamp 1586364061
transform 1 0 18400 0 -1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_199
timestamp 1586364061
transform 1 0 19412 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_36_211
timestamp 1586364061
transform 1 0 20516 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_43
timestamp 1586364061
transform 1 0 5060 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_46
timestamp 1586364061
transform 1 0 5336 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_53
timestamp 1586364061
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_57
timestamp 1586364061
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_71
timestamp 1586364061
transform 1 0 7636 0 1 22304
box -38 -48 406 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 8648 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 8096 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_75
timestamp 1586364061
transform 1 0 8004 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_78
timestamp 1586364061
transform 1 0 8280 0 1 22304
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_91
timestamp 1586364061
transform 1 0 9476 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _224_
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_108
timestamp 1586364061
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_112
timestamp 1586364061
transform 1 0 11408 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_116
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 12972 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_127
timestamp 1586364061
transform 1 0 12788 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_131
timestamp 1586364061
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use scs8hd_nor2_4  _108_
timestamp 1586364061
transform 1 0 15088 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 14904 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_144
timestamp 1586364061
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_148
timestamp 1586364061
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16100 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_161
timestamp 1586364061
transform 1 0 15916 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_165
timestamp 1586364061
transform 1 0 16284 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_37_177
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 590 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 18492 0 1 22304
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_193
timestamp 1586364061
transform 1 0 18860 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_197
timestamp 1586364061
transform 1 0 19228 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_209
timestamp 1586364061
transform 1 0 20332 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_221
timestamp 1586364061
transform 1 0 21436 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_37_233
timestamp 1586364061
transform 1 0 22540 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_37_241
timestamp 1586364061
transform 1 0 23276 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_38_47
timestamp 1586364061
transform 1 0 5428 0 -1 23392
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_64
timestamp 1586364061
transform 1 0 6992 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_84
timestamp 1586364061
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_106
timestamp 1586364061
transform 1 0 10856 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_119
timestamp 1586364061
transform 1 0 12052 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_123
timestamp 1586364061
transform 1 0 12420 0 -1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_126
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_136
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_142
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14352 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_38_146
timestamp 1586364061
transform 1 0 14536 0 -1 23392
box -38 -48 590 592
use scs8hd_fill_1  FILLER_38_152
timestamp 1586364061
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_157
timestamp 1586364061
transform 1 0 15548 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_169
timestamp 1586364061
transform 1 0 16652 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_181
timestamp 1586364061
transform 1 0 17756 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_193
timestamp 1586364061
transform 1 0 18860 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_205
timestamp 1586364061
transform 1 0 19964 0 -1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_38_213
timestamp 1586364061
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_17
timestamp 1586364061
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_6
timestamp 1586364061
transform 1 0 1656 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_21
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_40_30
timestamp 1586364061
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_6  FILLER_39_32
timestamp 1586364061
transform 1 0 4048 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_28
timestamp 1586364061
transform 1 0 3680 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_18
timestamp 1586364061
transform 1 0 2760 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4600 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5060 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_41
timestamp 1586364061
transform 1 0 4876 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_45
timestamp 1586364061
transform 1 0 5244 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 6992 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 7544 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_57
timestamp 1586364061
transform 1 0 6348 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_68
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 24480
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_72
timestamp 1586364061
transform 1 0 7728 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_83
timestamp 1586364061
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_87
timestamp 1586364061
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_40_84
timestamp 1586364061
transform 1 0 8832 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_97
timestamp 1586364061
transform 1 0 10028 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_97
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_91
timestamp 1586364061
transform 1 0 9476 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 9844 0 -1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 9660 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_40_107
timestamp 1586364061
transform 1 0 10948 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  FILLER_40_102
timestamp 1586364061
transform 1 0 10488 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_101
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 -1 24480
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_114
timestamp 1586364061
transform 1 0 11592 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _200_
timestamp 1586364061
transform 1 0 11224 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 -1 24480
box -38 -48 866 592
use scs8hd_buf_2  _220_
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__220__A
timestamp 1586364061
transform 1 0 13800 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_136
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_133
timestamp 1586364061
transform 1 0 13340 0 -1 24480
box -38 -48 774 592
use scs8hd_buf_2  _215_
timestamp 1586364061
transform 1 0 15548 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_149
timestamp 1586364061
transform 1 0 14812 0 1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_145
timestamp 1586364061
transform 1 0 14444 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _213_
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__215__A
timestamp 1586364061
transform 1 0 16100 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__213__A
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_161
timestamp 1586364061
transform 1 0 15916 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_165
timestamp 1586364061
transform 1 0 16284 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_173
timestamp 1586364061
transform 1 0 17020 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_177
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _225_
timestamp 1586364061
transform 1 0 18492 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 19044 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_193
timestamp 1586364061
transform 1 0 18860 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _222_
timestamp 1586364061
transform 1 0 20056 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_197
timestamp 1586364061
transform 1 0 19228 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_39_205
timestamp 1586364061
transform 1 0 19964 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_210
timestamp 1586364061
transform 1 0 20424 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_214
timestamp 1586364061
transform 1 0 20792 0 1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _218_
timestamp 1586364061
transform 1 0 21160 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__218__A
timestamp 1586364061
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_222
timestamp 1586364061
transform 1 0 21528 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_226
timestamp 1586364061
transform 1 0 21896 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_39_238
timestamp 1586364061
transform 1 0 23000 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8832 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use scs8hd_decap_8  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_82
timestamp 1586364061
transform 1 0 8648 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_87
timestamp 1586364061
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 10856 0 1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 10672 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_91
timestamp 1586364061
transform 1 0 9476 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_102
timestamp 1586364061
transform 1 0 10488 0 1 24480
box -38 -48 222 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11408 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_114
timestamp 1586364061
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_118
timestamp 1586364061
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_132
timestamp 1586364061
transform 1 0 13248 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_136
timestamp 1586364061
transform 1 0 13616 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_151
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_163
timestamp 1586364061
transform 1 0 16100 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_175
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_conb_1  _199_
timestamp 1586364061
transform 1 0 10396 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 590 592
use scs8hd_fill_1  FILLER_42_100
timestamp 1586364061
transform 1 0 10304 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_104
timestamp 1586364061
transform 1 0 10672 0 -1 25568
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 25568
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_115
timestamp 1586364061
transform 1 0 11684 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_1  FILLER_42_123
timestamp 1586364061
transform 1 0 12420 0 -1 25568
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_12.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 25568
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13156 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_6  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_8  FILLER_42_134
timestamp 1586364061
transform 1 0 13432 0 -1 25568
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_145
timestamp 1586364061
transform 1 0 14444 0 -1 25568
box -38 -48 774 592
use scs8hd_fill_2  FILLER_42_153
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 688 480 808 6 address[0]
port 0 nsew default input
rlabel metal3 s 0 2048 480 2168 6 address[1]
port 1 nsew default input
rlabel metal3 s 0 3544 480 3664 6 address[2]
port 2 nsew default input
rlabel metal2 s 478 27520 534 28000 6 address[3]
port 3 nsew default input
rlabel metal3 s 0 5040 480 5160 6 address[4]
port 4 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 address[5]
port 5 nsew default input
rlabel metal2 s 3054 0 3110 480 6 address[6]
port 6 nsew default input
rlabel metal3 s 0 8032 480 8152 6 bottom_left_grid_pin_11_
port 7 nsew default input
rlabel metal2 s 3422 27520 3478 28000 6 bottom_left_grid_pin_13_
port 8 nsew default input
rlabel metal2 s 4434 27520 4490 28000 6 bottom_left_grid_pin_15_
port 9 nsew default input
rlabel metal3 s 27520 960 28000 1080 6 bottom_left_grid_pin_1_
port 10 nsew default input
rlabel metal2 s 4342 0 4398 480 6 bottom_left_grid_pin_3_
port 11 nsew default input
rlabel metal3 s 0 6536 480 6656 6 bottom_left_grid_pin_5_
port 12 nsew default input
rlabel metal2 s 5630 0 5686 480 6 bottom_left_grid_pin_7_
port 13 nsew default input
rlabel metal2 s 2410 27520 2466 28000 6 bottom_left_grid_pin_9_
port 14 nsew default input
rlabel metal2 s 5446 27520 5502 28000 6 bottom_right_grid_pin_11_
port 15 nsew default input
rlabel metal3 s 27520 2864 28000 2984 6 chanx_right_in[0]
port 16 nsew default input
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_in[1]
port 17 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chanx_right_in[2]
port 18 nsew default input
rlabel metal2 s 6458 27520 6514 28000 6 chanx_right_in[3]
port 19 nsew default input
rlabel metal2 s 7470 27520 7526 28000 6 chanx_right_in[4]
port 20 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chanx_right_in[5]
port 21 nsew default input
rlabel metal3 s 27520 6944 28000 7064 6 chanx_right_in[6]
port 22 nsew default input
rlabel metal3 s 27520 8848 28000 8968 6 chanx_right_in[7]
port 23 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_right_in[8]
port 24 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chanx_right_out[0]
port 25 nsew default tristate
rlabel metal2 s 9402 27520 9458 28000 6 chanx_right_out[1]
port 26 nsew default tristate
rlabel metal2 s 10414 27520 10470 28000 6 chanx_right_out[2]
port 27 nsew default tristate
rlabel metal2 s 9402 0 9458 480 6 chanx_right_out[3]
port 28 nsew default tristate
rlabel metal2 s 11426 27520 11482 28000 6 chanx_right_out[4]
port 29 nsew default tristate
rlabel metal3 s 27520 10888 28000 11008 6 chanx_right_out[5]
port 30 nsew default tristate
rlabel metal2 s 10690 0 10746 480 6 chanx_right_out[6]
port 31 nsew default tristate
rlabel metal3 s 27520 12928 28000 13048 6 chanx_right_out[7]
port 32 nsew default tristate
rlabel metal2 s 12438 27520 12494 28000 6 chanx_right_out[8]
port 33 nsew default tristate
rlabel metal3 s 0 10888 480 11008 6 chany_bottom_in[0]
port 34 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[1]
port 35 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chany_bottom_in[2]
port 36 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chany_bottom_in[3]
port 37 nsew default input
rlabel metal2 s 13450 27520 13506 28000 6 chany_bottom_in[4]
port 38 nsew default input
rlabel metal2 s 14462 27520 14518 28000 6 chany_bottom_in[5]
port 39 nsew default input
rlabel metal2 s 13266 0 13322 480 6 chany_bottom_in[6]
port 40 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 chany_bottom_in[7]
port 41 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chany_bottom_in[8]
port 42 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_out[0]
port 43 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chany_bottom_out[1]
port 44 nsew default tristate
rlabel metal2 s 16394 27520 16450 28000 6 chany_bottom_out[2]
port 45 nsew default tristate
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_out[3]
port 46 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_bottom_out[4]
port 47 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[5]
port 48 nsew default tristate
rlabel metal2 s 18326 0 18382 480 6 chany_bottom_out[6]
port 49 nsew default tristate
rlabel metal3 s 27520 14968 28000 15088 6 chany_bottom_out[7]
port 50 nsew default tristate
rlabel metal3 s 27520 16872 28000 16992 6 chany_bottom_out[8]
port 51 nsew default tristate
rlabel metal3 s 27520 18912 28000 19032 6 chany_top_in[0]
port 52 nsew default input
rlabel metal3 s 0 18368 480 18488 6 chany_top_in[1]
port 53 nsew default input
rlabel metal3 s 0 19728 480 19848 6 chany_top_in[2]
port 54 nsew default input
rlabel metal3 s 27520 20952 28000 21072 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 19614 0 19670 480 6 chany_top_in[4]
port 56 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 18418 27520 18474 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 20902 0 20958 480 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 22098 0 22154 480 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 19430 27520 19486 28000 6 chany_top_out[0]
port 61 nsew default tristate
rlabel metal2 s 20442 27520 20498 28000 6 chany_top_out[1]
port 62 nsew default tristate
rlabel metal2 s 21454 27520 21510 28000 6 chany_top_out[2]
port 63 nsew default tristate
rlabel metal2 s 23386 0 23442 480 6 chany_top_out[3]
port 64 nsew default tristate
rlabel metal2 s 22374 27520 22430 28000 6 chany_top_out[4]
port 65 nsew default tristate
rlabel metal2 s 24674 0 24730 480 6 chany_top_out[5]
port 66 nsew default tristate
rlabel metal2 s 23386 27520 23442 28000 6 chany_top_out[6]
port 67 nsew default tristate
rlabel metal3 s 0 22720 480 22840 6 chany_top_out[7]
port 68 nsew default tristate
rlabel metal2 s 24398 27520 24454 28000 6 chany_top_out[8]
port 69 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 data_in
port 70 nsew default input
rlabel metal2 s 570 0 626 480 6 enable
port 71 nsew default input
rlabel metal3 s 0 24216 480 24336 6 right_bottom_grid_pin_12_
port 72 nsew default input
rlabel metal3 s 27520 22856 28000 22976 6 right_top_grid_pin_10_
port 73 nsew default input
rlabel metal2 s 27250 0 27306 480 6 top_left_grid_pin_11_
port 74 nsew default input
rlabel metal3 s 27520 26936 28000 27056 6 top_left_grid_pin_13_
port 75 nsew default input
rlabel metal3 s 0 25712 480 25832 6 top_left_grid_pin_15_
port 76 nsew default input
rlabel metal2 s 25410 27520 25466 28000 6 top_left_grid_pin_1_
port 77 nsew default input
rlabel metal2 s 26422 27520 26478 28000 6 top_left_grid_pin_3_
port 78 nsew default input
rlabel metal3 s 27520 24896 28000 25016 6 top_left_grid_pin_5_
port 79 nsew default input
rlabel metal2 s 25962 0 26018 480 6 top_left_grid_pin_7_
port 80 nsew default input
rlabel metal2 s 27434 27520 27490 28000 6 top_left_grid_pin_9_
port 81 nsew default input
rlabel metal3 s 0 27208 480 27328 6 top_right_grid_pin_11_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
