VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 123.000 BY 123.000 ;
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 119.000 85.470 123.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 119.000 88.690 123.000 ;
    END
  END SC_OUT_TOP
  PIN Test_en_E_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 34.040 123.000 34.640 ;
    END
  END Test_en_E_in
  PIN Test_en_E_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 31.320 123.000 31.920 ;
    END
  END Test_en_E_out
  PIN Test_en_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END Test_en_W_in
  PIN Test_en_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END Test_en_W_out
  PIN bottom_width_0_height_0__pin_50_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END bottom_width_0_height_0__pin_50_
  PIN bottom_width_0_height_0__pin_51_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END bottom_width_0_height_0__pin_51_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 27.920 123.000 28.520 ;
    END
  END ccff_tail
  PIN clk_0_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 119.000 91.910 123.000 ;
    END
  END clk_0_N_in
  PIN clk_0_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END clk_0_S_in
  PIN prog_clk_0_E_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 40.840 123.000 41.440 ;
    END
  END prog_clk_0_E_out
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 37.440 123.000 38.040 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_0_N_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 119.000 95.130 123.000 ;
    END
  END prog_clk_0_N_out
  PIN prog_clk_0_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END prog_clk_0_S_in
  PIN prog_clk_0_S_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END prog_clk_0_S_out
  PIN prog_clk_0_W_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END prog_clk_0_W_out
  PIN right_width_0_height_0__pin_16_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 44.240 123.000 44.840 ;
    END
  END right_width_0_height_0__pin_16_
  PIN right_width_0_height_0__pin_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 47.640 123.000 48.240 ;
    END
  END right_width_0_height_0__pin_17_
  PIN right_width_0_height_0__pin_18_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 51.040 123.000 51.640 ;
    END
  END right_width_0_height_0__pin_18_
  PIN right_width_0_height_0__pin_19_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 54.440 123.000 55.040 ;
    END
  END right_width_0_height_0__pin_19_
  PIN right_width_0_height_0__pin_20_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 57.840 123.000 58.440 ;
    END
  END right_width_0_height_0__pin_20_
  PIN right_width_0_height_0__pin_21_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 61.240 123.000 61.840 ;
    END
  END right_width_0_height_0__pin_21_
  PIN right_width_0_height_0__pin_22_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 63.960 123.000 64.560 ;
    END
  END right_width_0_height_0__pin_22_
  PIN right_width_0_height_0__pin_23_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 67.360 123.000 67.960 ;
    END
  END right_width_0_height_0__pin_23_
  PIN right_width_0_height_0__pin_24_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 70.760 123.000 71.360 ;
    END
  END right_width_0_height_0__pin_24_
  PIN right_width_0_height_0__pin_25_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 74.160 123.000 74.760 ;
    END
  END right_width_0_height_0__pin_25_
  PIN right_width_0_height_0__pin_26_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 77.560 123.000 78.160 ;
    END
  END right_width_0_height_0__pin_26_
  PIN right_width_0_height_0__pin_27_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 80.960 123.000 81.560 ;
    END
  END right_width_0_height_0__pin_27_
  PIN right_width_0_height_0__pin_28_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 84.360 123.000 84.960 ;
    END
  END right_width_0_height_0__pin_28_
  PIN right_width_0_height_0__pin_29_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 87.760 123.000 88.360 ;
    END
  END right_width_0_height_0__pin_29_
  PIN right_width_0_height_0__pin_30_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 91.160 123.000 91.760 ;
    END
  END right_width_0_height_0__pin_30_
  PIN right_width_0_height_0__pin_31_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 93.880 123.000 94.480 ;
    END
  END right_width_0_height_0__pin_31_
  PIN right_width_0_height_0__pin_42_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 1.400 123.000 2.000 ;
    END
  END right_width_0_height_0__pin_42_lower
  PIN right_width_0_height_0__pin_42_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 97.280 123.000 97.880 ;
    END
  END right_width_0_height_0__pin_42_upper
  PIN right_width_0_height_0__pin_43_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 4.120 123.000 4.720 ;
    END
  END right_width_0_height_0__pin_43_lower
  PIN right_width_0_height_0__pin_43_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 100.680 123.000 101.280 ;
    END
  END right_width_0_height_0__pin_43_upper
  PIN right_width_0_height_0__pin_44_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 7.520 123.000 8.120 ;
    END
  END right_width_0_height_0__pin_44_lower
  PIN right_width_0_height_0__pin_44_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 104.080 123.000 104.680 ;
    END
  END right_width_0_height_0__pin_44_upper
  PIN right_width_0_height_0__pin_45_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 10.920 123.000 11.520 ;
    END
  END right_width_0_height_0__pin_45_lower
  PIN right_width_0_height_0__pin_45_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 107.480 123.000 108.080 ;
    END
  END right_width_0_height_0__pin_45_upper
  PIN right_width_0_height_0__pin_46_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 14.320 123.000 14.920 ;
    END
  END right_width_0_height_0__pin_46_lower
  PIN right_width_0_height_0__pin_46_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 110.880 123.000 111.480 ;
    END
  END right_width_0_height_0__pin_46_upper
  PIN right_width_0_height_0__pin_47_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 17.720 123.000 18.320 ;
    END
  END right_width_0_height_0__pin_47_lower
  PIN right_width_0_height_0__pin_47_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 114.280 123.000 114.880 ;
    END
  END right_width_0_height_0__pin_47_upper
  PIN right_width_0_height_0__pin_48_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 21.120 123.000 21.720 ;
    END
  END right_width_0_height_0__pin_48_lower
  PIN right_width_0_height_0__pin_48_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 117.680 123.000 118.280 ;
    END
  END right_width_0_height_0__pin_48_upper
  PIN right_width_0_height_0__pin_49_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 24.520 123.000 25.120 ;
    END
  END right_width_0_height_0__pin_49_lower
  PIN right_width_0_height_0__pin_49_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.000 121.080 123.000 121.680 ;
    END
  END right_width_0_height_0__pin_49_upper
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 119.000 27.510 123.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 119.000 59.710 123.000 ;
    END
  END top_width_0_height_0__pin_10_
  PIN top_width_0_height_0__pin_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 119.000 62.930 123.000 ;
    END
  END top_width_0_height_0__pin_11_
  PIN top_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 119.000 66.150 123.000 ;
    END
  END top_width_0_height_0__pin_12_
  PIN top_width_0_height_0__pin_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 119.000 69.370 123.000 ;
    END
  END top_width_0_height_0__pin_13_
  PIN top_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 119.000 72.590 123.000 ;
    END
  END top_width_0_height_0__pin_14_
  PIN top_width_0_height_0__pin_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 119.000 75.810 123.000 ;
    END
  END top_width_0_height_0__pin_15_
  PIN top_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 119.000 30.730 123.000 ;
    END
  END top_width_0_height_0__pin_1_
  PIN top_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 119.000 33.950 123.000 ;
    END
  END top_width_0_height_0__pin_2_
  PIN top_width_0_height_0__pin_32_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 119.000 79.030 123.000 ;
    END
  END top_width_0_height_0__pin_32_
  PIN top_width_0_height_0__pin_33_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 119.000 82.250 123.000 ;
    END
  END top_width_0_height_0__pin_33_
  PIN top_width_0_height_0__pin_34_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 119.000 98.350 123.000 ;
    END
  END top_width_0_height_0__pin_34_lower
  PIN top_width_0_height_0__pin_34_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 119.000 1.750 123.000 ;
    END
  END top_width_0_height_0__pin_34_upper
  PIN top_width_0_height_0__pin_35_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 119.000 101.570 123.000 ;
    END
  END top_width_0_height_0__pin_35_lower
  PIN top_width_0_height_0__pin_35_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 119.000 4.970 123.000 ;
    END
  END top_width_0_height_0__pin_35_upper
  PIN top_width_0_height_0__pin_36_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 119.000 104.790 123.000 ;
    END
  END top_width_0_height_0__pin_36_lower
  PIN top_width_0_height_0__pin_36_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 119.000 8.190 123.000 ;
    END
  END top_width_0_height_0__pin_36_upper
  PIN top_width_0_height_0__pin_37_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 119.000 108.010 123.000 ;
    END
  END top_width_0_height_0__pin_37_lower
  PIN top_width_0_height_0__pin_37_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 119.000 11.410 123.000 ;
    END
  END top_width_0_height_0__pin_37_upper
  PIN top_width_0_height_0__pin_38_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 119.000 111.230 123.000 ;
    END
  END top_width_0_height_0__pin_38_lower
  PIN top_width_0_height_0__pin_38_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 119.000 14.630 123.000 ;
    END
  END top_width_0_height_0__pin_38_upper
  PIN top_width_0_height_0__pin_39_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 119.000 114.450 123.000 ;
    END
  END top_width_0_height_0__pin_39_lower
  PIN top_width_0_height_0__pin_39_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 119.000 17.850 123.000 ;
    END
  END top_width_0_height_0__pin_39_upper
  PIN top_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 119.000 37.170 123.000 ;
    END
  END top_width_0_height_0__pin_3_
  PIN top_width_0_height_0__pin_40_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 119.000 117.670 123.000 ;
    END
  END top_width_0_height_0__pin_40_lower
  PIN top_width_0_height_0__pin_40_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 119.000 21.070 123.000 ;
    END
  END top_width_0_height_0__pin_40_upper
  PIN top_width_0_height_0__pin_41_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 119.000 120.890 123.000 ;
    END
  END top_width_0_height_0__pin_41_lower
  PIN top_width_0_height_0__pin_41_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 119.000 24.290 123.000 ;
    END
  END top_width_0_height_0__pin_41_upper
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 119.000 40.390 123.000 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 119.000 43.610 123.000 ;
    END
  END top_width_0_height_0__pin_5_
  PIN top_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 119.000 46.830 123.000 ;
    END
  END top_width_0_height_0__pin_6_
  PIN top_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 119.000 50.050 123.000 ;
    END
  END top_width_0_height_0__pin_7_
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 119.000 53.270 123.000 ;
    END
  END top_width_0_height_0__pin_8_
  PIN top_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 119.000 56.490 123.000 ;
    END
  END top_width_0_height_0__pin_9_
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 98.020 10.640 99.620 111.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 60.700 10.640 62.300 111.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.380 10.640 24.980 111.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 79.360 10.640 80.960 111.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 42.040 10.640 43.640 111.760 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 118.075 111.605 ;
      LAYER met1 ;
        RECT 1.450 10.640 120.910 112.500 ;
      LAYER met2 ;
        RECT 2.030 118.720 4.410 121.565 ;
        RECT 5.250 118.720 7.630 121.565 ;
        RECT 8.470 118.720 10.850 121.565 ;
        RECT 11.690 118.720 14.070 121.565 ;
        RECT 14.910 118.720 17.290 121.565 ;
        RECT 18.130 118.720 20.510 121.565 ;
        RECT 21.350 118.720 23.730 121.565 ;
        RECT 24.570 118.720 26.950 121.565 ;
        RECT 27.790 118.720 30.170 121.565 ;
        RECT 31.010 118.720 33.390 121.565 ;
        RECT 34.230 118.720 36.610 121.565 ;
        RECT 37.450 118.720 39.830 121.565 ;
        RECT 40.670 118.720 43.050 121.565 ;
        RECT 43.890 118.720 46.270 121.565 ;
        RECT 47.110 118.720 49.490 121.565 ;
        RECT 50.330 118.720 52.710 121.565 ;
        RECT 53.550 118.720 55.930 121.565 ;
        RECT 56.770 118.720 59.150 121.565 ;
        RECT 59.990 118.720 62.370 121.565 ;
        RECT 63.210 118.720 65.590 121.565 ;
        RECT 66.430 118.720 68.810 121.565 ;
        RECT 69.650 118.720 72.030 121.565 ;
        RECT 72.870 118.720 75.250 121.565 ;
        RECT 76.090 118.720 78.470 121.565 ;
        RECT 79.310 118.720 81.690 121.565 ;
        RECT 82.530 118.720 84.910 121.565 ;
        RECT 85.750 118.720 88.130 121.565 ;
        RECT 88.970 118.720 91.350 121.565 ;
        RECT 92.190 118.720 94.570 121.565 ;
        RECT 95.410 118.720 97.790 121.565 ;
        RECT 98.630 118.720 101.010 121.565 ;
        RECT 101.850 118.720 104.230 121.565 ;
        RECT 105.070 118.720 107.450 121.565 ;
        RECT 108.290 118.720 110.670 121.565 ;
        RECT 111.510 118.720 113.890 121.565 ;
        RECT 114.730 118.720 117.110 121.565 ;
        RECT 117.950 118.720 120.330 121.565 ;
        RECT 1.480 4.280 120.880 118.720 ;
        RECT 1.480 1.515 9.930 4.280 ;
        RECT 10.770 1.515 30.170 4.280 ;
        RECT 31.010 1.515 50.870 4.280 ;
        RECT 51.710 1.515 71.110 4.280 ;
        RECT 71.950 1.515 91.810 4.280 ;
        RECT 92.650 1.515 112.050 4.280 ;
        RECT 112.890 1.515 120.880 4.280 ;
      LAYER met3 ;
        RECT 4.000 120.680 118.600 121.545 ;
        RECT 4.000 118.680 119.000 120.680 ;
        RECT 4.000 117.280 118.600 118.680 ;
        RECT 4.000 115.280 119.000 117.280 ;
        RECT 4.000 113.880 118.600 115.280 ;
        RECT 4.000 111.880 119.000 113.880 ;
        RECT 4.000 110.480 118.600 111.880 ;
        RECT 4.000 108.480 119.000 110.480 ;
        RECT 4.000 107.800 118.600 108.480 ;
        RECT 4.400 107.080 118.600 107.800 ;
        RECT 4.400 106.400 119.000 107.080 ;
        RECT 4.000 105.080 119.000 106.400 ;
        RECT 4.000 103.680 118.600 105.080 ;
        RECT 4.000 101.680 119.000 103.680 ;
        RECT 4.000 100.280 118.600 101.680 ;
        RECT 4.000 98.280 119.000 100.280 ;
        RECT 4.000 96.880 118.600 98.280 ;
        RECT 4.000 94.880 119.000 96.880 ;
        RECT 4.000 93.480 118.600 94.880 ;
        RECT 4.000 92.160 119.000 93.480 ;
        RECT 4.000 90.760 118.600 92.160 ;
        RECT 4.000 88.760 119.000 90.760 ;
        RECT 4.000 87.360 118.600 88.760 ;
        RECT 4.000 85.360 119.000 87.360 ;
        RECT 4.000 83.960 118.600 85.360 ;
        RECT 4.000 81.960 119.000 83.960 ;
        RECT 4.000 80.560 118.600 81.960 ;
        RECT 4.000 78.560 119.000 80.560 ;
        RECT 4.000 77.200 118.600 78.560 ;
        RECT 4.400 77.160 118.600 77.200 ;
        RECT 4.400 75.800 119.000 77.160 ;
        RECT 4.000 75.160 119.000 75.800 ;
        RECT 4.000 73.760 118.600 75.160 ;
        RECT 4.000 71.760 119.000 73.760 ;
        RECT 4.000 70.360 118.600 71.760 ;
        RECT 4.000 68.360 119.000 70.360 ;
        RECT 4.000 66.960 118.600 68.360 ;
        RECT 4.000 64.960 119.000 66.960 ;
        RECT 4.000 63.560 118.600 64.960 ;
        RECT 4.000 62.240 119.000 63.560 ;
        RECT 4.000 60.840 118.600 62.240 ;
        RECT 4.000 58.840 119.000 60.840 ;
        RECT 4.000 57.440 118.600 58.840 ;
        RECT 4.000 55.440 119.000 57.440 ;
        RECT 4.000 54.040 118.600 55.440 ;
        RECT 4.000 52.040 119.000 54.040 ;
        RECT 4.000 50.640 118.600 52.040 ;
        RECT 4.000 48.640 119.000 50.640 ;
        RECT 4.000 47.240 118.600 48.640 ;
        RECT 4.000 46.600 119.000 47.240 ;
        RECT 4.400 45.240 119.000 46.600 ;
        RECT 4.400 45.200 118.600 45.240 ;
        RECT 4.000 43.840 118.600 45.200 ;
        RECT 4.000 41.840 119.000 43.840 ;
        RECT 4.000 40.440 118.600 41.840 ;
        RECT 4.000 38.440 119.000 40.440 ;
        RECT 4.000 37.040 118.600 38.440 ;
        RECT 4.000 35.040 119.000 37.040 ;
        RECT 4.000 33.640 118.600 35.040 ;
        RECT 4.000 32.320 119.000 33.640 ;
        RECT 4.000 30.920 118.600 32.320 ;
        RECT 4.000 28.920 119.000 30.920 ;
        RECT 4.000 27.520 118.600 28.920 ;
        RECT 4.000 25.520 119.000 27.520 ;
        RECT 4.000 24.120 118.600 25.520 ;
        RECT 4.000 22.120 119.000 24.120 ;
        RECT 4.000 20.720 118.600 22.120 ;
        RECT 4.000 18.720 119.000 20.720 ;
        RECT 4.000 17.320 118.600 18.720 ;
        RECT 4.000 16.000 119.000 17.320 ;
        RECT 4.400 15.320 119.000 16.000 ;
        RECT 4.400 14.600 118.600 15.320 ;
        RECT 4.000 13.920 118.600 14.600 ;
        RECT 4.000 11.920 119.000 13.920 ;
        RECT 4.000 10.520 118.600 11.920 ;
        RECT 4.000 8.520 119.000 10.520 ;
        RECT 4.000 7.120 118.600 8.520 ;
        RECT 4.000 5.120 119.000 7.120 ;
        RECT 4.000 3.720 118.600 5.120 ;
        RECT 4.000 2.400 119.000 3.720 ;
        RECT 4.000 1.535 118.600 2.400 ;
      LAYER met4 ;
        RECT 96.895 41.655 97.225 46.065 ;
  END
END grid_clb
END LIBRARY

