VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__0_
  CLASS BLOCK ;
  FOREIGN cbx_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 80.000 ;
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 2.400 ;
    END
  END bottom_grid_pin_0_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 2.400 1.320 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 2.400 21.040 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 2.400 25.120 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 2.400 27.160 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.400 29.200 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 2.400 31.240 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 2.400 35.320 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.400 37.360 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 2.400 39.400 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 2.400 2.680 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 2.400 6.760 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 2.400 14.920 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 2.400 16.960 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.400 19.000 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.400 41.440 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 2.400 61.160 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 2.400 65.240 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 2.400 67.280 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 2.400 69.320 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 2.400 71.360 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 2.400 75.440 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 2.400 77.480 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 2.400 79.520 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 2.400 42.800 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 2.400 44.840 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 2.400 46.880 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 2.400 48.920 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 2.400 50.960 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 2.400 53.000 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 2.400 55.040 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.400 57.080 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 0.720 200.000 1.320 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 20.440 200.000 21.040 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 22.480 200.000 23.080 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 24.520 200.000 25.120 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 26.560 200.000 27.160 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 28.600 200.000 29.200 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 30.640 200.000 31.240 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 32.680 200.000 33.280 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 34.720 200.000 35.320 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 36.760 200.000 37.360 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 38.800 200.000 39.400 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 2.080 200.000 2.680 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 4.120 200.000 4.720 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 6.160 200.000 6.760 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 8.200 200.000 8.800 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 10.240 200.000 10.840 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 12.280 200.000 12.880 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 14.320 200.000 14.920 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 16.360 200.000 16.960 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 197.600 18.400 200.000 19.000 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 40.840 200.000 41.440 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 60.560 200.000 61.160 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 62.600 200.000 63.200 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 64.640 200.000 65.240 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 66.680 200.000 67.280 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 68.720 200.000 69.320 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 70.760 200.000 71.360 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 72.800 200.000 73.400 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 74.840 200.000 75.440 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 76.880 200.000 77.480 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 78.920 200.000 79.520 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 42.200 200.000 42.800 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 44.240 200.000 44.840 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 46.280 200.000 46.880 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 48.320 200.000 48.920 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 50.360 200.000 50.960 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 52.400 200.000 53.000 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 54.440 200.000 55.040 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 56.480 200.000 57.080 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 197.600 58.520 200.000 59.120 ;
    END
  END chanx_right_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 2.400 ;
    END
  END prog_clk
  PIN top_grid_pin_16_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.070 77.600 6.350 80.000 ;
    END
  END top_grid_pin_16_
  PIN top_grid_pin_17_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 77.600 18.770 80.000 ;
    END
  END top_grid_pin_17_
  PIN top_grid_pin_18_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 30.910 77.600 31.190 80.000 ;
    END
  END top_grid_pin_18_
  PIN top_grid_pin_19_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 43.330 77.600 43.610 80.000 ;
    END
  END top_grid_pin_19_
  PIN top_grid_pin_20_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.750 77.600 56.030 80.000 ;
    END
  END top_grid_pin_20_
  PIN top_grid_pin_21_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 77.600 68.450 80.000 ;
    END
  END top_grid_pin_21_
  PIN top_grid_pin_22_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 77.600 81.330 80.000 ;
    END
  END top_grid_pin_22_
  PIN top_grid_pin_23_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.470 77.600 93.750 80.000 ;
    END
  END top_grid_pin_23_
  PIN top_grid_pin_24_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 77.600 106.170 80.000 ;
    END
  END top_grid_pin_24_
  PIN top_grid_pin_25_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.310 77.600 118.590 80.000 ;
    END
  END top_grid_pin_25_
  PIN top_grid_pin_26_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 77.600 131.010 80.000 ;
    END
  END top_grid_pin_26_
  PIN top_grid_pin_27_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 143.610 77.600 143.890 80.000 ;
    END
  END top_grid_pin_27_
  PIN top_grid_pin_28_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 156.030 77.600 156.310 80.000 ;
    END
  END top_grid_pin_28_
  PIN top_grid_pin_29_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.450 77.600 168.730 80.000 ;
    END
  END top_grid_pin_29_
  PIN top_grid_pin_30_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.870 77.600 181.150 80.000 ;
    END
  END top_grid_pin_30_
  PIN top_grid_pin_31_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 193.290 77.600 193.570 80.000 ;
    END
  END top_grid_pin_31_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 38.055 10.640 39.655 68.240 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 71.385 10.640 72.985 68.240 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 68.085 ;
      LAYER met1 ;
        RECT 5.520 10.640 194.120 70.340 ;
      LAYER met2 ;
        RECT 6.630 77.320 18.210 79.405 ;
        RECT 19.050 77.320 30.630 79.405 ;
        RECT 31.470 77.320 43.050 79.405 ;
        RECT 43.890 77.320 55.470 79.405 ;
        RECT 56.310 77.320 67.890 79.405 ;
        RECT 68.730 77.320 80.770 79.405 ;
        RECT 81.610 77.320 93.190 79.405 ;
        RECT 94.030 77.320 105.610 79.405 ;
        RECT 106.450 77.320 118.030 79.405 ;
        RECT 118.870 77.320 130.450 79.405 ;
        RECT 131.290 77.320 143.330 79.405 ;
        RECT 144.170 77.320 155.750 79.405 ;
        RECT 156.590 77.320 168.170 79.405 ;
        RECT 169.010 77.320 180.590 79.405 ;
        RECT 181.430 77.320 193.010 79.405 ;
        RECT 6.080 2.680 193.570 77.320 ;
        RECT 6.080 0.835 24.650 2.680 ;
        RECT 25.490 0.835 74.330 2.680 ;
        RECT 75.170 0.835 124.470 2.680 ;
        RECT 125.310 0.835 174.610 2.680 ;
        RECT 175.450 0.835 193.570 2.680 ;
      LAYER met3 ;
        RECT 2.800 78.520 197.200 79.385 ;
        RECT 2.400 77.880 197.600 78.520 ;
        RECT 2.800 76.480 197.200 77.880 ;
        RECT 2.400 75.840 197.600 76.480 ;
        RECT 2.800 74.440 197.200 75.840 ;
        RECT 2.400 73.800 197.600 74.440 ;
        RECT 2.800 72.400 197.200 73.800 ;
        RECT 2.400 71.760 197.600 72.400 ;
        RECT 2.800 70.360 197.200 71.760 ;
        RECT 2.400 69.720 197.600 70.360 ;
        RECT 2.800 68.320 197.200 69.720 ;
        RECT 2.400 67.680 197.600 68.320 ;
        RECT 2.800 66.280 197.200 67.680 ;
        RECT 2.400 65.640 197.600 66.280 ;
        RECT 2.800 64.240 197.200 65.640 ;
        RECT 2.400 63.600 197.600 64.240 ;
        RECT 2.800 62.200 197.200 63.600 ;
        RECT 2.400 61.560 197.600 62.200 ;
        RECT 2.800 60.160 197.200 61.560 ;
        RECT 2.400 59.520 197.600 60.160 ;
        RECT 2.800 58.120 197.200 59.520 ;
        RECT 2.400 57.480 197.600 58.120 ;
        RECT 2.800 56.080 197.200 57.480 ;
        RECT 2.400 55.440 197.600 56.080 ;
        RECT 2.800 54.040 197.200 55.440 ;
        RECT 2.400 53.400 197.600 54.040 ;
        RECT 2.800 52.000 197.200 53.400 ;
        RECT 2.400 51.360 197.600 52.000 ;
        RECT 2.800 49.960 197.200 51.360 ;
        RECT 2.400 49.320 197.600 49.960 ;
        RECT 2.800 47.920 197.200 49.320 ;
        RECT 2.400 47.280 197.600 47.920 ;
        RECT 2.800 45.880 197.200 47.280 ;
        RECT 2.400 45.240 197.600 45.880 ;
        RECT 2.800 43.840 197.200 45.240 ;
        RECT 2.400 43.200 197.600 43.840 ;
        RECT 2.800 40.440 197.200 43.200 ;
        RECT 2.400 39.800 197.600 40.440 ;
        RECT 2.800 38.400 197.200 39.800 ;
        RECT 2.400 37.760 197.600 38.400 ;
        RECT 2.800 36.360 197.200 37.760 ;
        RECT 2.400 35.720 197.600 36.360 ;
        RECT 2.800 34.320 197.200 35.720 ;
        RECT 2.400 33.680 197.600 34.320 ;
        RECT 2.800 32.280 197.200 33.680 ;
        RECT 2.400 31.640 197.600 32.280 ;
        RECT 2.800 30.240 197.200 31.640 ;
        RECT 2.400 29.600 197.600 30.240 ;
        RECT 2.800 28.200 197.200 29.600 ;
        RECT 2.400 27.560 197.600 28.200 ;
        RECT 2.800 26.160 197.200 27.560 ;
        RECT 2.400 25.520 197.600 26.160 ;
        RECT 2.800 24.120 197.200 25.520 ;
        RECT 2.400 23.480 197.600 24.120 ;
        RECT 2.800 22.080 197.200 23.480 ;
        RECT 2.400 21.440 197.600 22.080 ;
        RECT 2.800 20.040 197.200 21.440 ;
        RECT 2.400 19.400 197.600 20.040 ;
        RECT 2.800 18.000 197.200 19.400 ;
        RECT 2.400 17.360 197.600 18.000 ;
        RECT 2.800 15.960 197.200 17.360 ;
        RECT 2.400 15.320 197.600 15.960 ;
        RECT 2.800 13.920 197.200 15.320 ;
        RECT 2.400 13.280 197.600 13.920 ;
        RECT 2.800 11.880 197.200 13.280 ;
        RECT 2.400 11.240 197.600 11.880 ;
        RECT 2.800 9.840 197.200 11.240 ;
        RECT 2.400 9.200 197.600 9.840 ;
        RECT 2.800 7.800 197.200 9.200 ;
        RECT 2.400 7.160 197.600 7.800 ;
        RECT 2.800 5.760 197.200 7.160 ;
        RECT 2.400 5.120 197.600 5.760 ;
        RECT 2.800 3.720 197.200 5.120 ;
        RECT 2.400 3.080 197.600 3.720 ;
        RECT 2.800 0.855 197.200 3.080 ;
      LAYER met4 ;
        RECT 22.870 10.640 37.655 68.240 ;
        RECT 40.055 10.640 70.985 68.240 ;
        RECT 73.385 10.640 180.450 68.240 ;
      LAYER met5 ;
        RECT 22.660 24.700 180.660 60.300 ;
  END
END cbx_1__0_
END LIBRARY

