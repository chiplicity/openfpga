magic
tech EFS8A
magscale 1 2
timestamp 1603810449
<< locali >>
rect 154825 389675 154859 389777
rect 145165 389539 145199 389641
rect 164393 389607 164427 389777
rect 167279 389573 167337 389607
rect 186507 389437 186565 389471
rect 135505 389335 135539 389437
rect 193465 388927 193499 389369
rect 249033 385595 249067 395149
rect 97325 350371 97359 351969
rect 186289 350983 186323 351833
rect 285005 350371 285039 351561
rect 75429 331603 75463 334765
rect 75429 330107 75463 331569
rect 75521 331671 75555 334697
rect 75981 334527 76015 344081
rect 75521 330175 75555 331637
rect 96865 329155 96899 329257
rect 87205 329019 87239 329121
rect 106433 329087 106467 329257
rect 186415 329053 186565 329087
rect 205735 329053 205977 329087
rect 109227 328985 109377 329019
rect 116185 328883 116219 328985
rect 119405 328883 119439 328985
rect 193465 328883 193499 328985
rect 203033 328883 203067 329053
rect 219685 329019 219719 329189
rect 266973 328951 267007 339321
rect 299725 331399 299759 331501
rect 309293 331399 309327 331569
rect 290065 329223 290099 329325
rect 283107 329189 283257 329223
rect 299633 329019 299667 329325
rect 319045 329087 319079 329189
rect 250447 327489 250631 327523
rect 250597 327251 250631 327489
rect 265317 327387 265351 328917
rect 256393 327251 256427 327353
rect 243789 327115 243823 327217
rect 152099 326401 152467 326435
rect 152433 326367 152467 326401
rect 157585 326367 157619 326673
rect 164485 326299 164519 326673
rect 256485 326367 256519 327217
rect 60249 319431 60283 320145
rect 64297 319635 64331 320417
rect 340389 320179 340423 320485
rect 341401 319975 341435 320281
rect 65033 319431 65067 319873
rect 352901 306987 352935 316541
rect 352993 279379 353027 290973
rect 342321 274687 342355 275061
rect 343333 274823 343367 275129
rect 156849 266119 156883 266629
rect 73957 262719 73991 263433
rect 74049 263399 74083 264385
rect 176445 246059 176479 246161
rect 77545 233003 77579 233105
rect 95393 233003 95427 233105
rect 96773 233003 96807 233173
rect 96865 233003 96899 233105
rect 101649 233003 101683 233105
rect 105145 232799 105179 233105
rect 250045 233105 250137 233139
rect 250045 233071 250079 233105
rect 222479 233037 222571 233071
rect 222537 233003 222571 233037
rect 114713 232799 114747 232901
rect 116185 232799 116219 232901
rect 120969 232799 121003 232969
rect 244525 232799 244559 232969
rect 358329 231031 358363 239293
rect 341953 224707 341987 225149
rect 345909 224775 345943 225421
rect 347933 223075 347967 225081
rect 348025 224775 348059 225081
rect 34857 213895 34891 220457
rect 369185 216479 369219 224129
rect 369921 221375 369955 229025
rect 34857 204715 34891 206857
rect 368725 192407 368759 195229
rect 348025 180847 348059 181697
rect 252253 172415 252287 172585
rect 252345 172279 252379 172585
rect 71657 168879 71691 169389
rect 271297 160651 271331 160753
rect 358605 156435 358639 163337
rect 76073 142087 76107 143957
rect 87113 143855 87147 143957
rect 302485 142087 302519 142189
rect 309385 142087 309419 142257
rect 318953 142155 318987 142257
rect 76073 140183 76107 142053
rect 157401 139571 157435 139673
rect 77545 139367 77579 139469
rect 87113 139299 87147 139469
rect 109285 139367 109319 139401
rect 109227 139333 109319 139367
rect 118485 139163 118519 139469
rect 124465 139163 124499 139333
rect 134125 139027 134159 139333
rect 143693 139027 143727 139129
rect 157585 138823 157619 139605
rect 158781 139571 158815 139877
rect 158045 139163 158079 139401
rect 162737 138823 162771 139673
rect 253357 139027 253391 139401
rect 253449 138959 253483 139333
rect 254093 139095 254127 139469
rect 254035 139061 254127 139095
rect 336801 130731 336835 131105
rect 345299 130833 345391 130867
rect 345357 130663 345391 130833
rect 51601 113731 51635 115125
rect 51693 107475 51727 108257
rect 51693 104075 51727 107441
rect 358329 95847 358363 105333
rect 26485 87007 26519 87449
rect 35961 87007 35995 87517
rect 36145 87143 36179 87449
rect 45713 87143 45747 87517
rect 45805 87143 45839 87381
rect 45897 87075 45931 87449
rect 51509 86123 51543 89013
rect 56109 87143 56143 87381
rect 65033 87075 65067 87449
rect 339929 86735 339963 86905
rect 64481 78983 64515 79153
rect 63929 78575 63963 78881
rect 67057 78507 67091 78745
rect 358421 76467 358455 86021
rect 88217 57155 88251 66709
rect 317573 57155 317607 66709
rect 193465 53211 193499 53313
rect 186749 53075 186783 53177
rect 203033 53143 203067 53313
rect 205793 53143 205827 53313
rect 174145 52871 174179 52973
rect 183713 52871 183747 53041
rect 96773 48519 96807 50933
rect 116185 47703 116219 47805
rect 109377 47635 109411 47669
rect 109227 47601 109411 47635
rect 95485 47431 95519 47533
rect 105053 47431 105087 47601
rect 125753 47567 125787 47805
rect 125845 47635 125879 47805
rect 135413 47703 135447 47805
rect 125879 47465 126029 47499
rect 317481 46139 317515 55013
rect 289973 45595 290007 46037
rect 298253 45595 298287 46037
rect 298345 45663 298379 45833
rect 283165 45527 283199 45561
rect 283107 45493 283199 45527
rect 278565 45323 278599 45493
rect 317113 37843 317147 44813
rect 358421 37843 358455 40597
rect 358237 18531 358271 28085
<< viali >>
rect 249033 395149 249067 395183
rect 154825 389777 154859 389811
rect 145165 389641 145199 389675
rect 154825 389641 154859 389675
rect 164393 389777 164427 389811
rect 164393 389573 164427 389607
rect 167245 389573 167279 389607
rect 167337 389573 167371 389607
rect 145165 389505 145199 389539
rect 135505 389437 135539 389471
rect 186473 389437 186507 389471
rect 186565 389437 186599 389471
rect 135505 389301 135539 389335
rect 193465 389369 193499 389403
rect 193465 388893 193499 388927
rect 249033 385561 249067 385595
rect 97325 351969 97359 352003
rect 186289 351833 186323 351867
rect 186289 350949 186323 350983
rect 285005 351561 285039 351595
rect 97325 350337 97359 350371
rect 285005 350337 285039 350371
rect 75981 344081 76015 344115
rect 75429 334765 75463 334799
rect 75429 331569 75463 331603
rect 75521 334697 75555 334731
rect 75981 334493 76015 334527
rect 266973 339321 267007 339355
rect 75521 331637 75555 331671
rect 75521 330141 75555 330175
rect 75429 330073 75463 330107
rect 96865 329257 96899 329291
rect 87205 329121 87239 329155
rect 96865 329121 96899 329155
rect 106433 329257 106467 329291
rect 219685 329189 219719 329223
rect 106433 329053 106467 329087
rect 186381 329053 186415 329087
rect 186565 329053 186599 329087
rect 203033 329053 203067 329087
rect 205701 329053 205735 329087
rect 205977 329053 206011 329087
rect 87205 328985 87239 329019
rect 109193 328985 109227 329019
rect 109377 328985 109411 329019
rect 116185 328985 116219 329019
rect 116185 328849 116219 328883
rect 119405 328985 119439 329019
rect 119405 328849 119439 328883
rect 193465 328985 193499 329019
rect 193465 328849 193499 328883
rect 219685 328985 219719 329019
rect 309293 331569 309327 331603
rect 299725 331501 299759 331535
rect 299725 331365 299759 331399
rect 309293 331365 309327 331399
rect 290065 329325 290099 329359
rect 283073 329189 283107 329223
rect 283257 329189 283291 329223
rect 290065 329189 290099 329223
rect 299633 329325 299667 329359
rect 319045 329189 319079 329223
rect 319045 329053 319079 329087
rect 299633 328985 299667 329019
rect 203033 328849 203067 328883
rect 265317 328917 265351 328951
rect 266973 328917 267007 328951
rect 250413 327489 250447 327523
rect 243789 327217 243823 327251
rect 250597 327217 250631 327251
rect 256393 327353 256427 327387
rect 265317 327353 265351 327387
rect 256393 327217 256427 327251
rect 256485 327217 256519 327251
rect 243789 327081 243823 327115
rect 157585 326673 157619 326707
rect 152065 326401 152099 326435
rect 152433 326333 152467 326367
rect 157585 326333 157619 326367
rect 164485 326673 164519 326707
rect 256485 326333 256519 326367
rect 164485 326265 164519 326299
rect 340389 320485 340423 320519
rect 64297 320417 64331 320451
rect 60249 320145 60283 320179
rect 340389 320145 340423 320179
rect 341401 320281 341435 320315
rect 341401 319941 341435 319975
rect 64297 319601 64331 319635
rect 65033 319873 65067 319907
rect 60249 319397 60283 319431
rect 65033 319397 65067 319431
rect 352901 316541 352935 316575
rect 352901 306953 352935 306987
rect 352993 290973 353027 291007
rect 352993 279345 353027 279379
rect 343333 275129 343367 275163
rect 342321 275061 342355 275095
rect 343333 274789 343367 274823
rect 342321 274653 342355 274687
rect 156849 266629 156883 266663
rect 156849 266085 156883 266119
rect 74049 264385 74083 264419
rect 73957 263433 73991 263467
rect 74049 263365 74083 263399
rect 73957 262685 73991 262719
rect 176445 246161 176479 246195
rect 176445 246025 176479 246059
rect 358329 239293 358363 239327
rect 96773 233173 96807 233207
rect 77545 233105 77579 233139
rect 77545 232969 77579 233003
rect 95393 233105 95427 233139
rect 95393 232969 95427 233003
rect 96773 232969 96807 233003
rect 96865 233105 96899 233139
rect 96865 232969 96899 233003
rect 101649 233105 101683 233139
rect 101649 232969 101683 233003
rect 105145 233105 105179 233139
rect 250137 233105 250171 233139
rect 222445 233037 222479 233071
rect 250045 233037 250079 233071
rect 120969 232969 121003 233003
rect 222537 232969 222571 233003
rect 244525 232969 244559 233003
rect 105145 232765 105179 232799
rect 114713 232901 114747 232935
rect 114713 232765 114747 232799
rect 116185 232901 116219 232935
rect 116185 232765 116219 232799
rect 120969 232765 121003 232799
rect 244525 232765 244559 232799
rect 358329 230997 358363 231031
rect 369921 229025 369955 229059
rect 345909 225421 345943 225455
rect 341953 225149 341987 225183
rect 345909 224741 345943 224775
rect 347933 225081 347967 225115
rect 341953 224673 341987 224707
rect 348025 225081 348059 225115
rect 348025 224741 348059 224775
rect 347933 223041 347967 223075
rect 369185 224129 369219 224163
rect 34857 220457 34891 220491
rect 369921 221341 369955 221375
rect 369185 216445 369219 216479
rect 34857 213861 34891 213895
rect 34857 206857 34891 206891
rect 34857 204681 34891 204715
rect 368725 195229 368759 195263
rect 368725 192373 368759 192407
rect 348025 181697 348059 181731
rect 348025 180813 348059 180847
rect 252253 172585 252287 172619
rect 252253 172381 252287 172415
rect 252345 172585 252379 172619
rect 252345 172245 252379 172279
rect 71657 169389 71691 169423
rect 71657 168845 71691 168879
rect 358605 163337 358639 163371
rect 271297 160753 271331 160787
rect 271297 160617 271331 160651
rect 358605 156401 358639 156435
rect 76073 143957 76107 143991
rect 87113 143957 87147 143991
rect 87113 143821 87147 143855
rect 309385 142257 309419 142291
rect 76073 142053 76107 142087
rect 302485 142189 302519 142223
rect 302485 142053 302519 142087
rect 318953 142257 318987 142291
rect 318953 142121 318987 142155
rect 309385 142053 309419 142087
rect 76073 140149 76107 140183
rect 158781 139877 158815 139911
rect 157401 139673 157435 139707
rect 157401 139537 157435 139571
rect 157585 139605 157619 139639
rect 77545 139469 77579 139503
rect 77545 139333 77579 139367
rect 87113 139469 87147 139503
rect 118485 139469 118519 139503
rect 109285 139401 109319 139435
rect 109193 139333 109227 139367
rect 87113 139265 87147 139299
rect 118485 139129 118519 139163
rect 124465 139333 124499 139367
rect 124465 139129 124499 139163
rect 134125 139333 134159 139367
rect 134125 138993 134159 139027
rect 143693 139129 143727 139163
rect 143693 138993 143727 139027
rect 158781 139537 158815 139571
rect 162737 139673 162771 139707
rect 158045 139401 158079 139435
rect 158045 139129 158079 139163
rect 157585 138789 157619 138823
rect 254093 139469 254127 139503
rect 253357 139401 253391 139435
rect 253357 138993 253391 139027
rect 253449 139333 253483 139367
rect 254001 139061 254035 139095
rect 253449 138925 253483 138959
rect 162737 138789 162771 138823
rect 336801 131105 336835 131139
rect 345265 130833 345299 130867
rect 336801 130697 336835 130731
rect 345357 130629 345391 130663
rect 51601 115125 51635 115159
rect 51601 113697 51635 113731
rect 51693 108257 51727 108291
rect 51693 107441 51727 107475
rect 51693 104041 51727 104075
rect 358329 105333 358363 105367
rect 358329 95813 358363 95847
rect 51509 89013 51543 89047
rect 35961 87517 35995 87551
rect 26485 87449 26519 87483
rect 26485 86973 26519 87007
rect 45713 87517 45747 87551
rect 36145 87449 36179 87483
rect 36145 87109 36179 87143
rect 45897 87449 45931 87483
rect 45713 87109 45747 87143
rect 45805 87381 45839 87415
rect 45805 87109 45839 87143
rect 45897 87041 45931 87075
rect 35961 86973 35995 87007
rect 65033 87449 65067 87483
rect 56109 87381 56143 87415
rect 56109 87109 56143 87143
rect 65033 87041 65067 87075
rect 339929 86905 339963 86939
rect 339929 86701 339963 86735
rect 51509 86089 51543 86123
rect 358421 86021 358455 86055
rect 64481 79153 64515 79187
rect 64481 78949 64515 78983
rect 63929 78881 63963 78915
rect 63929 78541 63963 78575
rect 67057 78745 67091 78779
rect 67057 78473 67091 78507
rect 358421 76433 358455 76467
rect 88217 66709 88251 66743
rect 88217 57121 88251 57155
rect 317573 66709 317607 66743
rect 317573 57121 317607 57155
rect 317481 55013 317515 55047
rect 193465 53313 193499 53347
rect 186749 53177 186783 53211
rect 193465 53177 193499 53211
rect 203033 53313 203067 53347
rect 203033 53109 203067 53143
rect 205793 53313 205827 53347
rect 205793 53109 205827 53143
rect 183713 53041 183747 53075
rect 186749 53041 186783 53075
rect 174145 52973 174179 53007
rect 174145 52837 174179 52871
rect 183713 52837 183747 52871
rect 96773 50933 96807 50967
rect 96773 48485 96807 48519
rect 116185 47805 116219 47839
rect 109377 47669 109411 47703
rect 116185 47669 116219 47703
rect 125753 47805 125787 47839
rect 105053 47601 105087 47635
rect 109193 47601 109227 47635
rect 95485 47533 95519 47567
rect 95485 47397 95519 47431
rect 125845 47805 125879 47839
rect 135413 47805 135447 47839
rect 135413 47669 135447 47703
rect 125845 47601 125879 47635
rect 125753 47533 125787 47567
rect 125845 47465 125879 47499
rect 126029 47465 126063 47499
rect 105053 47397 105087 47431
rect 317481 46105 317515 46139
rect 289973 46037 290007 46071
rect 283165 45561 283199 45595
rect 289973 45561 290007 45595
rect 298253 46037 298287 46071
rect 298345 45833 298379 45867
rect 298345 45629 298379 45663
rect 298253 45561 298287 45595
rect 278565 45493 278599 45527
rect 283073 45493 283107 45527
rect 278565 45289 278599 45323
rect 317113 44813 317147 44847
rect 317113 37809 317147 37843
rect 358421 40597 358455 40631
rect 358421 37809 358455 37843
rect 358237 28085 358271 28119
rect 358237 18497 358271 18531
<< metal1 >>
rect 249018 395180 249024 395192
rect 248979 395152 249024 395180
rect 249018 395140 249024 395152
rect 249076 395140 249082 395192
rect 88570 393780 88576 393832
rect 88628 393820 88634 393832
rect 89582 393820 89588 393832
rect 88628 393792 89588 393820
rect 88628 393780 88634 393792
rect 89582 393780 89588 393792
rect 89640 393780 89646 393832
rect 106510 393780 106516 393832
rect 106568 393820 106574 393832
rect 107246 393820 107252 393832
rect 106568 393792 107252 393820
rect 106568 393780 106574 393792
rect 107246 393780 107252 393792
rect 107304 393780 107310 393832
rect 124450 393780 124456 393832
rect 124508 393820 124514 393832
rect 125002 393820 125008 393832
rect 124508 393792 125008 393820
rect 124508 393780 124514 393792
rect 125002 393780 125008 393792
rect 125060 393780 125066 393832
rect 212770 393780 212776 393832
rect 212828 393820 212834 393832
rect 213506 393820 213512 393832
rect 212828 393792 213512 393820
rect 212828 393780 212834 393792
rect 213506 393780 213512 393792
rect 213564 393780 213570 393832
rect 355186 393780 355192 393832
rect 355244 393820 355250 393832
rect 358590 393820 358596 393832
rect 355244 393792 358596 393820
rect 355244 393780 355250 393792
rect 358590 393780 358596 393792
rect 358648 393780 358654 393832
rect 70630 393644 70636 393696
rect 70688 393684 70694 393696
rect 71826 393684 71832 393696
rect 70688 393656 71832 393684
rect 70688 393644 70694 393656
rect 71826 393644 71832 393656
rect 71884 393644 71890 393696
rect 337522 393372 337528 393424
rect 337580 393412 337586 393424
rect 358498 393412 358504 393424
rect 337580 393384 358504 393412
rect 337580 393372 337586 393384
rect 358498 393372 358504 393384
rect 358556 393372 358562 393424
rect 304586 393304 304592 393356
rect 304644 393344 304650 393356
rect 408362 393344 408368 393356
rect 304644 393316 408368 393344
rect 304644 393304 304650 393316
rect 408362 393304 408368 393316
rect 408420 393304 408426 393356
rect 299434 393236 299440 393288
rect 299492 393276 299498 393288
rect 426026 393276 426032 393288
rect 299492 393248 426032 393276
rect 299492 393236 299498 393248
rect 426026 393236 426032 393248
rect 426084 393236 426090 393288
rect 106326 393168 106332 393220
rect 106384 393208 106390 393220
rect 372942 393208 372948 393220
rect 106384 393180 372948 393208
rect 106384 393168 106390 393180
rect 372942 393168 372948 393180
rect 373000 393168 373006 393220
rect 91330 393100 91336 393152
rect 91388 393140 91394 393152
rect 390606 393140 390612 393152
rect 91388 393112 390612 393140
rect 91388 393100 91394 393112
rect 390606 393100 390612 393112
rect 390664 393100 390670 393152
rect 18190 392760 18196 392812
rect 18248 392800 18254 392812
rect 18742 392800 18748 392812
rect 18248 392772 18748 392800
rect 18248 392760 18254 392772
rect 18742 392760 18748 392772
rect 18800 392760 18806 392812
rect 154813 389811 154871 389817
rect 154813 389777 154825 389811
rect 154859 389808 154871 389811
rect 164381 389811 164439 389817
rect 164381 389808 164393 389811
rect 154859 389780 164393 389808
rect 154859 389777 154871 389780
rect 154813 389771 154871 389777
rect 164381 389777 164393 389780
rect 164427 389777 164439 389811
rect 164381 389771 164439 389777
rect 314614 389700 314620 389752
rect 314672 389740 314678 389752
rect 429430 389740 429436 389752
rect 314672 389712 429436 389740
rect 314672 389700 314678 389712
rect 429430 389700 429436 389712
rect 429488 389700 429494 389752
rect 145153 389675 145211 389681
rect 145153 389641 145165 389675
rect 145199 389672 145211 389675
rect 154813 389675 154871 389681
rect 154813 389672 154825 389675
rect 145199 389644 154825 389672
rect 145199 389641 145211 389644
rect 145153 389635 145211 389641
rect 154813 389641 154825 389644
rect 154859 389641 154871 389675
rect 154813 389635 154871 389641
rect 164381 389607 164439 389613
rect 164381 389573 164393 389607
rect 164427 389604 164439 389607
rect 167233 389607 167291 389613
rect 167233 389604 167245 389607
rect 164427 389576 167245 389604
rect 164427 389573 164439 389576
rect 164381 389567 164439 389573
rect 167233 389573 167245 389576
rect 167279 389573 167291 389607
rect 167233 389567 167291 389573
rect 167325 389607 167383 389613
rect 167325 389573 167337 389607
rect 167371 389604 167383 389607
rect 167371 389576 174084 389604
rect 167371 389573 167383 389576
rect 167325 389567 167383 389573
rect 145153 389539 145211 389545
rect 145153 389536 145165 389539
rect 145076 389508 145165 389536
rect 135493 389471 135551 389477
rect 135493 389437 135505 389471
rect 135539 389468 135551 389471
rect 145076 389468 145104 389508
rect 145153 389505 145165 389508
rect 145199 389505 145211 389539
rect 174056 389536 174084 389576
rect 174056 389508 176844 389536
rect 145153 389499 145211 389505
rect 135539 389440 145104 389468
rect 176816 389468 176844 389508
rect 186461 389471 186519 389477
rect 186461 389468 186473 389471
rect 176816 389440 186473 389468
rect 135539 389437 135551 389440
rect 135493 389431 135551 389437
rect 186461 389437 186473 389440
rect 186507 389437 186519 389471
rect 186461 389431 186519 389437
rect 186553 389471 186611 389477
rect 186553 389437 186565 389471
rect 186599 389468 186611 389471
rect 186599 389440 188528 389468
rect 186599 389437 186611 389440
rect 186553 389431 186611 389437
rect 188500 389400 188528 389440
rect 193453 389403 193511 389409
rect 193453 389400 193465 389403
rect 188500 389372 193465 389400
rect 193453 389369 193465 389372
rect 193499 389369 193511 389403
rect 193453 389363 193511 389369
rect 70630 389292 70636 389344
rect 70688 389332 70694 389344
rect 111294 389332 111300 389344
rect 70688 389304 111300 389332
rect 70688 389292 70694 389304
rect 111294 389292 111300 389304
rect 111352 389292 111358 389344
rect 135493 389335 135551 389341
rect 135493 389332 135505 389335
rect 128608 389304 135505 389332
rect 54070 389224 54076 389276
rect 54128 389264 54134 389276
rect 116262 389264 116268 389276
rect 54128 389236 116268 389264
rect 54128 389224 54134 389236
rect 116262 389224 116268 389236
rect 116320 389224 116326 389276
rect 124450 389224 124456 389276
rect 124508 389264 124514 389276
rect 128608 389264 128636 389304
rect 135493 389301 135505 389304
rect 135539 389301 135551 389335
rect 135493 389295 135551 389301
rect 124508 389236 128636 389264
rect 124508 389224 124514 389236
rect 142666 389224 142672 389276
rect 142724 389264 142730 389276
rect 194830 389264 194836 389276
rect 142724 389236 194836 389264
rect 142724 389224 142730 389236
rect 194830 389224 194836 389236
rect 194888 389224 194894 389276
rect 195842 389224 195848 389276
rect 195900 389264 195906 389276
rect 283978 389264 283984 389276
rect 195900 389236 283984 389264
rect 195900 389224 195906 389236
rect 283978 389224 283984 389236
rect 284036 389224 284042 389276
rect 106510 389156 106516 389208
rect 106568 389196 106574 389208
rect 205318 389196 205324 389208
rect 106568 389168 205324 389196
rect 106568 389156 106574 389168
rect 205318 389156 205324 389168
rect 205376 389156 205382 389208
rect 36130 389088 36136 389140
rect 36188 389128 36194 389140
rect 121322 389128 121328 389140
rect 36188 389100 121328 389128
rect 36188 389088 36194 389100
rect 121322 389088 121328 389100
rect 121380 389088 121386 389140
rect 178086 389088 178092 389140
rect 178144 389128 178150 389140
rect 288946 389128 288952 389140
rect 178144 389100 288952 389128
rect 178144 389088 178150 389100
rect 288946 389088 288952 389100
rect 289004 389088 289010 389140
rect 88570 389020 88576 389072
rect 88628 389060 88634 389072
rect 210286 389060 210292 389072
rect 88628 389032 210292 389060
rect 88628 389020 88634 389032
rect 210286 389020 210292 389032
rect 210344 389020 210350 389072
rect 212770 389020 212776 389072
rect 212828 389060 212834 389072
rect 279010 389060 279016 389072
rect 212828 389032 279016 389060
rect 212828 389020 212834 389032
rect 279010 389020 279016 389032
rect 279068 389020 279074 389072
rect 18190 388952 18196 389004
rect 18248 388992 18254 389004
rect 126290 388992 126296 389004
rect 18248 388964 126296 388992
rect 18248 388952 18254 388964
rect 126290 388952 126296 388964
rect 126348 388952 126354 389004
rect 160422 388952 160428 389004
rect 160480 388992 160486 389004
rect 294190 388992 294196 389004
rect 160480 388964 294196 388992
rect 160480 388952 160486 388964
rect 294190 388952 294196 388964
rect 294248 388952 294254 389004
rect 193453 388927 193511 388933
rect 193453 388893 193465 388927
rect 193499 388924 193511 388927
rect 200350 388924 200356 388936
rect 193499 388896 200356 388924
rect 193499 388893 193511 388896
rect 193453 388887 193511 388893
rect 200350 388884 200356 388896
rect 200408 388884 200414 388936
rect 96298 388544 96304 388596
rect 96356 388584 96362 388596
rect 127854 388584 127860 388596
rect 96356 388556 127860 388584
rect 96356 388544 96362 388556
rect 127854 388544 127860 388556
rect 127912 388544 127918 388596
rect 185354 388544 185360 388596
rect 185412 388584 185418 388596
rect 228594 388584 228600 388596
rect 185412 388556 228600 388584
rect 185412 388544 185418 388556
rect 228594 388544 228600 388556
rect 228652 388544 228658 388596
rect 13406 388476 13412 388528
rect 13464 388516 13470 388528
rect 101266 388516 101272 388528
rect 13464 388488 101272 388516
rect 13464 388476 13470 388488
rect 101266 388476 101272 388488
rect 101324 388476 101330 388528
rect 190322 388476 190328 388528
rect 190380 388516 190386 388528
rect 265854 388516 265860 388528
rect 190380 388488 265860 388516
rect 190380 388476 190386 388488
rect 265854 388476 265860 388488
rect 265912 388476 265918 388528
rect 13498 388408 13504 388460
rect 13556 388448 13562 388460
rect 215346 388448 215352 388460
rect 13556 388420 215352 388448
rect 13556 388408 13562 388420
rect 215346 388408 215352 388420
rect 215404 388408 215410 388460
rect 220314 388408 220320 388460
rect 220372 388448 220378 388460
rect 315626 388448 315632 388460
rect 220372 388420 315632 388448
rect 220372 388408 220378 388420
rect 315626 388408 315632 388420
rect 315684 388408 315690 388460
rect 13590 388340 13596 388392
rect 13648 388380 13654 388392
rect 309002 388380 309008 388392
rect 13648 388352 309008 388380
rect 13648 388340 13654 388352
rect 309002 388340 309008 388352
rect 309060 388340 309066 388392
rect 249021 385595 249079 385601
rect 249021 385561 249033 385595
rect 249067 385592 249079 385595
rect 249110 385592 249116 385604
rect 249067 385564 249116 385592
rect 249067 385561 249079 385564
rect 249021 385555 249079 385561
rect 249110 385552 249116 385564
rect 249168 385552 249174 385604
rect 226478 382764 226484 382816
rect 226536 382804 226542 382816
rect 227214 382804 227220 382816
rect 226536 382776 227220 382804
rect 226536 382764 226542 382776
rect 227214 382764 227220 382776
rect 227272 382804 227278 382816
rect 230894 382804 230900 382816
rect 227272 382776 230900 382804
rect 227272 382764 227278 382776
rect 230894 382764 230900 382776
rect 230952 382764 230958 382816
rect 315810 378616 315816 378668
rect 315868 378656 315874 378668
rect 429430 378656 429436 378668
rect 315868 378628 429436 378656
rect 315868 378616 315874 378628
rect 429430 378616 429436 378628
rect 429488 378616 429494 378668
rect 248926 375896 248932 375948
rect 248984 375936 248990 375948
rect 249018 375936 249024 375948
rect 248984 375908 249024 375936
rect 248984 375896 248990 375908
rect 249018 375896 249024 375908
rect 249076 375896 249082 375948
rect 226478 375148 226484 375200
rect 226536 375188 226542 375200
rect 228778 375188 228784 375200
rect 226536 375160 228784 375188
rect 226536 375148 226542 375160
rect 228778 375148 228784 375160
rect 228836 375188 228842 375200
rect 248926 375188 248932 375200
rect 228836 375160 248932 375188
rect 228836 375148 228842 375160
rect 248926 375148 248932 375160
rect 248984 375148 248990 375200
rect 266590 373176 266596 373228
rect 266648 373216 266654 373228
rect 266774 373216 266780 373228
rect 266648 373188 266780 373216
rect 266648 373176 266654 373188
rect 266774 373176 266780 373188
rect 266832 373176 266838 373228
rect 131810 371748 131816 371800
rect 131868 371788 131874 371800
rect 134754 371788 134760 371800
rect 131868 371760 134760 371788
rect 131868 371748 131874 371760
rect 134754 371748 134760 371760
rect 134812 371748 134818 371800
rect 225834 371748 225840 371800
rect 225892 371788 225898 371800
rect 229974 371788 229980 371800
rect 225892 371760 229980 371788
rect 225892 371748 225898 371760
rect 229974 371748 229980 371760
rect 230032 371748 230038 371800
rect 320318 371748 320324 371800
rect 320376 371788 320382 371800
rect 362454 371788 362460 371800
rect 320376 371760 362460 371788
rect 320376 371748 320382 371760
rect 362454 371748 362460 371760
rect 362512 371748 362518 371800
rect 186274 368620 186280 368672
rect 186332 368660 186338 368672
rect 191518 368660 191524 368672
rect 186332 368632 191524 368660
rect 186332 368620 186338 368632
rect 191518 368620 191524 368632
rect 191576 368620 191582 368672
rect 208998 368552 209004 368604
rect 209056 368592 209062 368604
rect 210010 368592 210016 368604
rect 209056 368564 210016 368592
rect 209056 368552 209062 368564
rect 210010 368552 210016 368564
rect 210068 368552 210074 368604
rect 277538 368280 277544 368332
rect 277596 368320 277602 368332
rect 280390 368320 280396 368332
rect 277596 368292 280396 368320
rect 277596 368280 277602 368292
rect 280390 368280 280396 368292
rect 280448 368280 280454 368332
rect 89858 367668 89864 367720
rect 89916 367708 89922 367720
rect 92526 367708 92532 367720
rect 89916 367680 92532 367708
rect 89916 367668 89922 367680
rect 92526 367668 92532 367680
rect 92584 367668 92590 367720
rect 90042 367600 90048 367652
rect 90100 367640 90106 367652
rect 91422 367640 91428 367652
rect 90100 367612 91428 367640
rect 90100 367600 90106 367612
rect 91422 367600 91428 367612
rect 91480 367600 91486 367652
rect 95010 367600 95016 367652
rect 95068 367640 95074 367652
rect 96850 367640 96856 367652
rect 95068 367612 96856 367640
rect 95068 367600 95074 367612
rect 96850 367600 96856 367612
rect 96908 367600 96914 367652
rect 99978 367600 99984 367652
rect 100036 367640 100042 367652
rect 100898 367640 100904 367652
rect 100036 367612 100904 367640
rect 100036 367600 100042 367612
rect 100898 367600 100904 367612
rect 100956 367600 100962 367652
rect 105038 367600 105044 367652
rect 105096 367640 105102 367652
rect 106602 367640 106608 367652
rect 105096 367612 106608 367640
rect 105096 367600 105102 367612
rect 106602 367600 106608 367612
rect 106660 367600 106666 367652
rect 110006 367600 110012 367652
rect 110064 367640 110070 367652
rect 112030 367640 112036 367652
rect 110064 367612 112036 367640
rect 110064 367600 110070 367612
rect 112030 367600 112036 367612
rect 112088 367600 112094 367652
rect 114974 367600 114980 367652
rect 115032 367640 115038 367652
rect 116170 367640 116176 367652
rect 115032 367612 116176 367640
rect 115032 367600 115038 367612
rect 116170 367600 116176 367612
rect 116228 367600 116234 367652
rect 120034 367600 120040 367652
rect 120092 367640 120098 367652
rect 121690 367640 121696 367652
rect 120092 367612 121696 367640
rect 120092 367600 120098 367612
rect 121690 367600 121696 367612
rect 121748 367600 121754 367652
rect 184066 367600 184072 367652
rect 184124 367640 184130 367652
rect 185170 367640 185176 367652
rect 184124 367612 185176 367640
rect 184124 367600 184130 367612
rect 185170 367600 185176 367612
rect 185228 367600 185234 367652
rect 185262 367600 185268 367652
rect 185320 367640 185326 367652
rect 186550 367640 186556 367652
rect 185320 367612 186556 367640
rect 185320 367600 185326 367612
rect 186550 367600 186556 367612
rect 186608 367600 186614 367652
rect 199062 367600 199068 367652
rect 199120 367640 199126 367652
rect 200258 367640 200264 367652
rect 199120 367612 200264 367640
rect 199120 367600 199126 367612
rect 200258 367600 200264 367612
rect 200316 367600 200322 367652
rect 204030 367600 204036 367652
rect 204088 367640 204094 367652
rect 205870 367640 205876 367652
rect 204088 367612 205876 367640
rect 204088 367600 204094 367612
rect 205870 367600 205876 367612
rect 205928 367600 205934 367652
rect 214058 367600 214064 367652
rect 214116 367640 214122 367652
rect 215530 367640 215536 367652
rect 214116 367612 215536 367640
rect 214116 367600 214122 367612
rect 215530 367600 215536 367612
rect 215588 367600 215594 367652
rect 278366 367600 278372 367652
rect 278424 367640 278430 367652
rect 279654 367640 279660 367652
rect 278424 367612 279660 367640
rect 278424 367600 278430 367612
rect 279654 367600 279660 367612
rect 279712 367600 279718 367652
rect 282966 367600 282972 367652
rect 283024 367640 283030 367652
rect 283794 367640 283800 367652
rect 283024 367612 283800 367640
rect 283024 367600 283030 367612
rect 283794 367600 283800 367612
rect 283852 367600 283858 367652
rect 293362 367600 293368 367652
rect 293420 367640 293426 367652
rect 294282 367640 294288 367652
rect 293420 367612 294288 367640
rect 293420 367600 293426 367612
rect 294282 367600 294288 367612
rect 294340 367600 294346 367652
rect 298238 367600 298244 367652
rect 298296 367640 298302 367652
rect 299710 367640 299716 367652
rect 298296 367612 299716 367640
rect 298296 367600 298302 367612
rect 299710 367600 299716 367612
rect 299768 367600 299774 367652
rect 303298 367600 303304 367652
rect 303356 367640 303362 367652
rect 305230 367640 305236 367652
rect 303356 367612 305236 367640
rect 303356 367600 303362 367612
rect 305230 367600 305236 367612
rect 305288 367600 305294 367652
rect 308358 367600 308364 367652
rect 308416 367640 308422 367652
rect 309278 367640 309284 367652
rect 308416 367612 309284 367640
rect 308416 367600 308422 367612
rect 309278 367600 309284 367612
rect 309336 367600 309342 367652
rect 127854 366172 127860 366224
rect 127912 366212 127918 366224
rect 429430 366212 429436 366224
rect 127912 366184 429436 366212
rect 127912 366172 127918 366184
rect 429430 366172 429436 366184
rect 429488 366172 429494 366224
rect 266590 363520 266596 363572
rect 266648 363560 266654 363572
rect 266774 363560 266780 363572
rect 266648 363532 266780 363560
rect 266648 363520 266654 363532
rect 266774 363520 266780 363532
rect 266832 363520 266838 363572
rect 116170 363452 116176 363504
rect 116228 363492 116234 363504
rect 116998 363492 117004 363504
rect 116228 363464 117004 363492
rect 116228 363452 116234 363464
rect 116998 363452 117004 363464
rect 117056 363452 117062 363504
rect 210010 363452 210016 363504
rect 210068 363492 210074 363504
rect 211022 363492 211028 363504
rect 210068 363464 211028 363492
rect 210068 363452 210074 363464
rect 211022 363452 211028 363464
rect 211080 363452 211086 363504
rect 67686 359848 67692 359900
rect 67744 359888 67750 359900
rect 75966 359888 75972 359900
rect 67744 359860 75972 359888
rect 67744 359848 67750 359860
rect 75966 359848 75972 359860
rect 76024 359848 76030 359900
rect 53702 359780 53708 359832
rect 53760 359820 53766 359832
rect 76978 359820 76984 359832
rect 53760 359792 76984 359820
rect 53760 359780 53766 359792
rect 76978 359780 76984 359792
rect 77036 359780 77042 359832
rect 50206 359712 50212 359764
rect 50264 359752 50270 359764
rect 76794 359752 76800 359764
rect 50264 359724 76800 359752
rect 50264 359712 50270 359724
rect 76794 359712 76800 359724
rect 76852 359712 76858 359764
rect 64190 359644 64196 359696
rect 64248 359684 64254 359696
rect 75690 359684 75696 359696
rect 64248 359656 75696 359684
rect 64248 359644 64254 359656
rect 75690 359644 75696 359656
rect 75748 359644 75754 359696
rect 60694 359576 60700 359628
rect 60752 359616 60758 359628
rect 75782 359616 75788 359628
rect 60752 359588 75788 359616
rect 60752 359576 60758 359588
rect 75782 359576 75788 359588
rect 75840 359576 75846 359628
rect 57198 359508 57204 359560
rect 57256 359548 57262 359560
rect 76058 359548 76064 359560
rect 57256 359520 76064 359548
rect 57256 359508 57262 359520
rect 76058 359508 76064 359520
rect 76116 359508 76122 359560
rect 71182 359372 71188 359424
rect 71240 359412 71246 359424
rect 75874 359412 75880 359424
rect 71240 359384 75880 359412
rect 71240 359372 71246 359384
rect 75874 359372 75880 359384
rect 75932 359372 75938 359424
rect 185170 358624 185176 358676
rect 185228 358664 185234 358676
rect 185998 358664 186004 358676
rect 185228 358636 186004 358664
rect 185228 358624 185234 358636
rect 185998 358624 186004 358636
rect 186056 358624 186062 358676
rect 80198 357876 80204 357928
rect 80256 357916 80262 357928
rect 127210 357916 127216 357928
rect 80256 357888 127216 357916
rect 80256 357876 80262 357888
rect 127210 357876 127216 357888
rect 127268 357916 127274 357928
rect 139630 357916 139636 357928
rect 127268 357888 139636 357916
rect 127268 357876 127274 357888
rect 139630 357876 139636 357888
rect 139688 357876 139694 357928
rect 174038 357876 174044 357928
rect 174096 357916 174102 357928
rect 221050 357916 221056 357928
rect 174096 357888 221056 357916
rect 174096 357876 174102 357888
rect 221050 357876 221056 357888
rect 221108 357916 221114 357928
rect 233470 357916 233476 357928
rect 221108 357888 233476 357916
rect 221108 357876 221114 357888
rect 233470 357876 233476 357888
rect 233528 357876 233534 357928
rect 267326 357876 267332 357928
rect 267384 357916 267390 357928
rect 314890 357916 314896 357928
rect 267384 357888 314896 357916
rect 267384 357876 267390 357888
rect 314890 357876 314896 357888
rect 314948 357916 314954 357928
rect 328414 357916 328420 357928
rect 314948 357888 328420 357916
rect 314948 357876 314954 357888
rect 328414 357876 328420 357888
rect 328472 357876 328478 357928
rect 75690 357536 75696 357588
rect 75748 357576 75754 357588
rect 76426 357576 76432 357588
rect 75748 357548 76432 357576
rect 75748 357536 75754 357548
rect 76426 357536 76432 357548
rect 76484 357536 76490 357588
rect 75782 357468 75788 357520
rect 75840 357508 75846 357520
rect 76150 357508 76156 357520
rect 75840 357480 76156 357508
rect 75840 357468 75846 357480
rect 76150 357468 76156 357480
rect 76208 357468 76214 357520
rect 74770 357400 74776 357452
rect 74828 357440 74834 357452
rect 76886 357440 76892 357452
rect 74828 357412 76892 357440
rect 74828 357400 74834 357412
rect 76886 357400 76892 357412
rect 76944 357400 76950 357452
rect 80198 356516 80204 356568
rect 80256 356556 80262 356568
rect 121782 356556 121788 356568
rect 80256 356528 121788 356556
rect 80256 356516 80262 356528
rect 121782 356516 121788 356528
rect 121840 356556 121846 356568
rect 139630 356556 139636 356568
rect 121840 356528 139636 356556
rect 121840 356516 121846 356528
rect 139630 356516 139636 356528
rect 139688 356516 139694 356568
rect 173486 356516 173492 356568
rect 173544 356556 173550 356568
rect 215622 356556 215628 356568
rect 173544 356528 215628 356556
rect 173544 356516 173550 356528
rect 215622 356516 215628 356528
rect 215680 356556 215686 356568
rect 233470 356556 233476 356568
rect 215680 356528 233476 356556
rect 215680 356516 215686 356528
rect 233470 356516 233476 356528
rect 233528 356516 233534 356568
rect 266590 356516 266596 356568
rect 266648 356556 266654 356568
rect 266774 356556 266780 356568
rect 266648 356528 266780 356556
rect 266648 356516 266654 356528
rect 266774 356516 266780 356528
rect 266832 356516 266838 356568
rect 267878 356516 267884 356568
rect 267936 356556 267942 356568
rect 309370 356556 309376 356568
rect 267936 356528 309376 356556
rect 267936 356516 267942 356528
rect 309370 356516 309376 356528
rect 309428 356556 309434 356568
rect 328322 356556 328328 356568
rect 309428 356528 328328 356556
rect 309428 356516 309434 356528
rect 328322 356516 328328 356528
rect 328380 356516 328386 356568
rect 80198 355156 80204 355208
rect 80256 355196 80262 355208
rect 117550 355196 117556 355208
rect 80256 355168 117556 355196
rect 80256 355156 80262 355168
rect 117550 355156 117556 355168
rect 117608 355196 117614 355208
rect 139630 355196 139636 355208
rect 117608 355168 139636 355196
rect 117608 355156 117614 355168
rect 139630 355156 139636 355168
rect 139688 355156 139694 355208
rect 174038 355156 174044 355208
rect 174096 355196 174102 355208
rect 211390 355196 211396 355208
rect 174096 355168 211396 355196
rect 174096 355156 174102 355168
rect 211390 355156 211396 355168
rect 211448 355196 211454 355208
rect 233470 355196 233476 355208
rect 211448 355168 233476 355196
rect 211448 355156 211454 355168
rect 233470 355156 233476 355168
rect 233528 355156 233534 355208
rect 266774 355156 266780 355208
rect 266832 355196 266838 355208
rect 266866 355196 266872 355208
rect 266832 355168 266872 355196
rect 266832 355156 266838 355168
rect 266866 355156 266872 355168
rect 266924 355156 266930 355208
rect 267878 355156 267884 355208
rect 267936 355196 267942 355208
rect 305322 355196 305328 355208
rect 267936 355168 305328 355196
rect 267936 355156 267942 355168
rect 305322 355156 305328 355168
rect 305380 355196 305386 355208
rect 328414 355196 328420 355208
rect 305380 355168 328420 355196
rect 305380 355156 305386 355168
rect 328414 355156 328420 355168
rect 328472 355156 328478 355208
rect 79278 355088 79284 355140
rect 79336 355128 79342 355140
rect 112122 355128 112128 355140
rect 79336 355100 112128 355128
rect 79336 355088 79342 355100
rect 112122 355088 112128 355100
rect 112180 355128 112186 355140
rect 139722 355128 139728 355140
rect 112180 355100 139728 355128
rect 112180 355088 112186 355100
rect 139722 355088 139728 355100
rect 139780 355088 139786 355140
rect 173762 355088 173768 355140
rect 173820 355128 173826 355140
rect 205962 355128 205968 355140
rect 173820 355100 205968 355128
rect 173820 355088 173826 355100
rect 205962 355088 205968 355100
rect 206020 355128 206026 355140
rect 233562 355128 233568 355140
rect 206020 355100 233568 355128
rect 206020 355088 206026 355100
rect 233562 355088 233568 355100
rect 233620 355088 233626 355140
rect 267418 355088 267424 355140
rect 267476 355128 267482 355140
rect 299802 355128 299808 355140
rect 267476 355100 299808 355128
rect 267476 355088 267482 355100
rect 299802 355088 299808 355100
rect 299860 355128 299866 355140
rect 328506 355128 328512 355140
rect 299860 355100 328512 355128
rect 299860 355088 299866 355100
rect 328506 355088 328512 355100
rect 328564 355088 328570 355140
rect 100898 355020 100904 355072
rect 100956 355060 100962 355072
rect 102370 355060 102376 355072
rect 100956 355032 102376 355060
rect 100956 355020 100962 355032
rect 102370 355020 102376 355032
rect 102428 355020 102434 355072
rect 125738 355020 125744 355072
rect 125796 355060 125802 355072
rect 127210 355060 127216 355072
rect 125796 355032 127216 355060
rect 125796 355020 125802 355032
rect 127210 355020 127216 355032
rect 127268 355020 127274 355072
rect 194738 355020 194744 355072
rect 194796 355060 194802 355072
rect 196302 355060 196308 355072
rect 194796 355032 196308 355060
rect 194796 355020 194802 355032
rect 196302 355020 196308 355032
rect 196360 355020 196366 355072
rect 279654 355020 279660 355072
rect 279712 355060 279718 355072
rect 280390 355060 280396 355072
rect 279712 355032 280396 355060
rect 279712 355020 279718 355032
rect 280390 355020 280396 355032
rect 280448 355020 280454 355072
rect 283794 355020 283800 355072
rect 283852 355060 283858 355072
rect 285358 355060 285364 355072
rect 283852 355032 285364 355060
rect 283852 355020 283858 355032
rect 285358 355020 285364 355032
rect 285416 355020 285422 355072
rect 288578 355020 288584 355072
rect 288636 355060 288642 355072
rect 290326 355060 290332 355072
rect 288636 355032 290332 355060
rect 288636 355020 288642 355032
rect 290326 355020 290332 355032
rect 290384 355020 290390 355072
rect 309278 355020 309284 355072
rect 309336 355060 309342 355072
rect 310382 355060 310388 355072
rect 309336 355032 310388 355060
rect 309336 355020 309342 355032
rect 310382 355020 310388 355032
rect 310440 355020 310446 355072
rect 313418 355020 313424 355072
rect 313476 355060 313482 355072
rect 315350 355060 315356 355072
rect 313476 355032 315356 355060
rect 313476 355020 313482 355032
rect 315350 355020 315356 355032
rect 315408 355020 315414 355072
rect 76058 354000 76064 354052
rect 76116 354040 76122 354052
rect 76116 354012 76288 354040
rect 76116 354000 76122 354012
rect 76260 353916 76288 354012
rect 189218 354000 189224 354052
rect 189276 354040 189282 354052
rect 191334 354040 191340 354052
rect 189276 354012 191340 354040
rect 189276 354000 189282 354012
rect 191334 354000 191340 354012
rect 191392 354000 191398 354052
rect 200258 354000 200264 354052
rect 200316 354040 200322 354052
rect 201362 354040 201368 354052
rect 200316 354012 201368 354040
rect 200316 354000 200322 354012
rect 201362 354000 201368 354012
rect 201420 354000 201426 354052
rect 76242 353864 76248 353916
rect 76300 353864 76306 353916
rect 219578 353864 219584 353916
rect 219636 353904 219642 353916
rect 221326 353904 221332 353916
rect 219636 353876 221332 353904
rect 219636 353864 219642 353876
rect 221326 353864 221332 353876
rect 221384 353864 221390 353916
rect 78910 353796 78916 353848
rect 78968 353836 78974 353848
rect 106510 353836 106516 353848
rect 78968 353808 106516 353836
rect 78968 353796 78974 353808
rect 106510 353796 106516 353808
rect 106568 353836 106574 353848
rect 139630 353836 139636 353848
rect 106568 353808 139636 353836
rect 106568 353796 106574 353808
rect 139630 353796 139636 353808
rect 139688 353796 139694 353848
rect 174038 353796 174044 353848
rect 174096 353836 174102 353848
rect 200350 353836 200356 353848
rect 174096 353808 200356 353836
rect 174096 353796 174102 353808
rect 200350 353796 200356 353808
rect 200408 353836 200414 353848
rect 233470 353836 233476 353848
rect 200408 353808 233476 353836
rect 200408 353796 200414 353808
rect 233470 353796 233476 353808
rect 233528 353796 233534 353848
rect 267878 353796 267884 353848
rect 267936 353836 267942 353848
rect 294190 353836 294196 353848
rect 267936 353808 294196 353836
rect 267936 353796 267942 353808
rect 294190 353796 294196 353808
rect 294248 353836 294254 353848
rect 328046 353836 328052 353848
rect 294248 353808 328052 353836
rect 294248 353796 294254 353808
rect 328046 353796 328052 353808
rect 328104 353796 328110 353848
rect 80198 352368 80204 352420
rect 80256 352408 80262 352420
rect 102646 352408 102652 352420
rect 80256 352380 102652 352408
rect 80256 352368 80262 352380
rect 102646 352368 102652 352380
rect 102704 352408 102710 352420
rect 139630 352408 139636 352420
rect 102704 352380 139636 352408
rect 102704 352368 102710 352380
rect 139630 352368 139636 352380
rect 139688 352368 139694 352420
rect 174038 352368 174044 352420
rect 174096 352408 174102 352420
rect 196210 352408 196216 352420
rect 174096 352380 196216 352408
rect 174096 352368 174102 352380
rect 196210 352368 196216 352380
rect 196268 352408 196274 352420
rect 233470 352408 233476 352420
rect 196268 352380 233476 352408
rect 196268 352368 196274 352380
rect 233470 352368 233476 352380
rect 233528 352368 233534 352420
rect 267878 352368 267884 352420
rect 267936 352408 267942 352420
rect 290050 352408 290056 352420
rect 267936 352380 290056 352408
rect 267936 352368 267942 352380
rect 290050 352368 290056 352380
rect 290108 352408 290114 352420
rect 328506 352408 328512 352420
rect 290108 352380 328512 352408
rect 290108 352368 290114 352380
rect 328506 352368 328512 352380
rect 328564 352368 328570 352420
rect 97310 352000 97316 352012
rect 97271 351972 97316 352000
rect 97310 351960 97316 351972
rect 97368 351960 97374 352012
rect 186274 351864 186280 351876
rect 186235 351836 186280 351864
rect 186274 351824 186280 351836
rect 186332 351824 186338 351876
rect 284990 351592 284996 351604
rect 284951 351564 284996 351592
rect 284990 351552 284996 351564
rect 285048 351552 285054 351604
rect 226294 351280 226300 351332
rect 226352 351320 226358 351332
rect 231630 351320 231636 351332
rect 226352 351292 231636 351320
rect 226352 351280 226358 351292
rect 231630 351280 231636 351292
rect 231688 351280 231694 351332
rect 131810 351076 131816 351128
rect 131868 351116 131874 351128
rect 137422 351116 137428 351128
rect 131868 351088 137428 351116
rect 131868 351076 131874 351088
rect 137422 351076 137428 351088
rect 137480 351076 137486 351128
rect 320594 351076 320600 351128
rect 320652 351116 320658 351128
rect 327218 351116 327224 351128
rect 320652 351088 327224 351116
rect 320652 351076 320658 351088
rect 327218 351076 327224 351088
rect 327276 351076 327282 351128
rect 79094 351008 79100 351060
rect 79152 351048 79158 351060
rect 89858 351048 89864 351060
rect 79152 351020 89864 351048
rect 79152 351008 79158 351020
rect 89858 351008 89864 351020
rect 89916 351048 89922 351060
rect 139630 351048 139636 351060
rect 89916 351020 139636 351048
rect 89916 351008 89922 351020
rect 139630 351008 139636 351020
rect 139688 351008 139694 351060
rect 173762 351008 173768 351060
rect 173820 351048 173826 351060
rect 185262 351048 185268 351060
rect 173820 351020 185268 351048
rect 173820 351008 173826 351020
rect 185262 351008 185268 351020
rect 185320 351048 185326 351060
rect 233562 351048 233568 351060
rect 185320 351020 233568 351048
rect 185320 351008 185326 351020
rect 233562 351008 233568 351020
rect 233620 351008 233626 351060
rect 267510 351008 267516 351060
rect 267568 351048 267574 351060
rect 277538 351048 277544 351060
rect 267568 351020 277544 351048
rect 267568 351008 267574 351020
rect 277538 351008 277544 351020
rect 277596 351048 277602 351060
rect 327862 351048 327868 351060
rect 277596 351020 327868 351048
rect 277596 351008 277602 351020
rect 327862 351008 327868 351020
rect 327920 351008 327926 351060
rect 174038 350940 174044 350992
rect 174096 350980 174102 350992
rect 186277 350983 186335 350989
rect 186277 350980 186289 350983
rect 174096 350952 186289 350980
rect 174096 350940 174102 350952
rect 186277 350949 186289 350952
rect 186323 350980 186335 350983
rect 233470 350980 233476 350992
rect 186323 350952 233476 350980
rect 186323 350949 186335 350952
rect 186277 350943 186335 350949
rect 233470 350940 233476 350952
rect 233528 350940 233534 350992
rect 80198 350328 80204 350380
rect 80256 350368 80262 350380
rect 97313 350371 97371 350377
rect 97313 350368 97325 350371
rect 80256 350340 97325 350368
rect 80256 350328 80262 350340
rect 97313 350337 97325 350340
rect 97359 350368 97371 350371
rect 139722 350368 139728 350380
rect 97359 350340 139728 350368
rect 97359 350337 97371 350340
rect 97313 350331 97371 350337
rect 139722 350328 139728 350340
rect 139780 350328 139786 350380
rect 267694 350328 267700 350380
rect 267752 350368 267758 350380
rect 284993 350371 285051 350377
rect 284993 350368 285005 350371
rect 267752 350340 285005 350368
rect 267752 350328 267758 350340
rect 284993 350337 285005 350340
rect 285039 350368 285051 350371
rect 327494 350368 327500 350380
rect 285039 350340 327500 350368
rect 285039 350337 285051 350340
rect 284993 350331 285051 350337
rect 327494 350328 327500 350340
rect 327552 350328 327558 350380
rect 131810 349716 131816 349768
rect 131868 349756 131874 349768
rect 137514 349756 137520 349768
rect 131868 349728 137520 349756
rect 131868 349716 131874 349728
rect 137514 349716 137520 349728
rect 137572 349716 137578 349768
rect 226386 349716 226392 349768
rect 226444 349756 226450 349768
rect 231170 349756 231176 349768
rect 226444 349728 231176 349756
rect 226444 349716 226450 349728
rect 231170 349716 231176 349728
rect 231228 349716 231234 349768
rect 321606 349716 321612 349768
rect 321664 349756 321670 349768
rect 327126 349756 327132 349768
rect 321664 349728 327132 349756
rect 321664 349716 321670 349728
rect 327126 349716 327132 349728
rect 327184 349716 327190 349768
rect 80198 349648 80204 349700
rect 80256 349688 80262 349700
rect 87190 349688 87196 349700
rect 80256 349660 87196 349688
rect 80256 349648 80262 349660
rect 87190 349648 87196 349660
rect 87248 349648 87254 349700
rect 137422 349648 137428 349700
rect 137480 349688 137486 349700
rect 139630 349688 139636 349700
rect 137480 349660 139636 349688
rect 137480 349648 137486 349660
rect 139630 349648 139636 349660
rect 139688 349648 139694 349700
rect 231630 349648 231636 349700
rect 231688 349688 231694 349700
rect 233470 349688 233476 349700
rect 231688 349660 233476 349688
rect 231688 349648 231694 349660
rect 233470 349648 233476 349660
rect 233528 349648 233534 349700
rect 267878 349648 267884 349700
rect 267936 349688 267942 349700
rect 274778 349688 274784 349700
rect 267936 349660 274784 349688
rect 267936 349648 267942 349660
rect 274778 349648 274784 349660
rect 274836 349648 274842 349700
rect 173026 349036 173032 349088
rect 173084 349076 173090 349088
rect 180846 349076 180852 349088
rect 173084 349048 180852 349076
rect 173084 349036 173090 349048
rect 180846 349036 180852 349048
rect 180904 349036 180910 349088
rect 321606 348424 321612 348476
rect 321664 348464 321670 348476
rect 327034 348464 327040 348476
rect 321664 348436 327040 348464
rect 321664 348424 321670 348436
rect 327034 348424 327040 348436
rect 327092 348424 327098 348476
rect 131902 348356 131908 348408
rect 131960 348396 131966 348408
rect 137422 348396 137428 348408
rect 131960 348368 137428 348396
rect 131960 348356 131966 348368
rect 137422 348356 137428 348368
rect 137480 348356 137486 348408
rect 226386 348356 226392 348408
rect 226444 348396 226450 348408
rect 233286 348396 233292 348408
rect 226444 348368 233292 348396
rect 226444 348356 226450 348368
rect 233286 348356 233292 348368
rect 233344 348356 233350 348408
rect 131810 348288 131816 348340
rect 131868 348328 131874 348340
rect 137606 348328 137612 348340
rect 131868 348300 137612 348328
rect 131868 348288 131874 348300
rect 137606 348288 137612 348300
rect 137664 348288 137670 348340
rect 226478 348288 226484 348340
rect 226536 348328 226542 348340
rect 233378 348328 233384 348340
rect 226536 348300 233384 348328
rect 226536 348288 226542 348300
rect 233378 348288 233384 348300
rect 233436 348288 233442 348340
rect 320686 348288 320692 348340
rect 320744 348328 320750 348340
rect 327218 348328 327224 348340
rect 320744 348300 327224 348328
rect 320744 348288 320750 348300
rect 327218 348288 327224 348300
rect 327276 348288 327282 348340
rect 80198 348220 80204 348272
rect 80256 348260 80262 348272
rect 87466 348260 87472 348272
rect 80256 348232 87472 348260
rect 80256 348220 80262 348232
rect 87466 348220 87472 348232
rect 87524 348220 87530 348272
rect 137514 348220 137520 348272
rect 137572 348260 137578 348272
rect 139630 348260 139636 348272
rect 137572 348232 139636 348260
rect 137572 348220 137578 348232
rect 139630 348220 139636 348232
rect 139688 348220 139694 348272
rect 231170 348220 231176 348272
rect 231228 348260 231234 348272
rect 233470 348260 233476 348272
rect 231228 348232 233476 348260
rect 231228 348220 231234 348232
rect 233470 348220 233476 348232
rect 233528 348220 233534 348272
rect 267878 348220 267884 348272
rect 267936 348260 267942 348272
rect 274962 348260 274968 348272
rect 267936 348232 274968 348260
rect 267936 348220 267942 348232
rect 274962 348220 274968 348232
rect 275020 348220 275026 348272
rect 172934 347948 172940 348000
rect 172992 347988 172998 348000
rect 180938 347988 180944 348000
rect 172992 347960 180944 347988
rect 172992 347948 172998 347960
rect 180938 347948 180944 347960
rect 180996 347948 181002 348000
rect 132178 346928 132184 346980
rect 132236 346968 132242 346980
rect 139814 346968 139820 346980
rect 132236 346940 139820 346968
rect 132236 346928 132242 346940
rect 139814 346928 139820 346940
rect 139872 346928 139878 346980
rect 226386 346928 226392 346980
rect 226444 346968 226450 346980
rect 228410 346968 228416 346980
rect 226444 346940 228416 346968
rect 226444 346928 226450 346940
rect 228410 346928 228416 346940
rect 228468 346928 228474 346980
rect 321054 346928 321060 346980
rect 321112 346968 321118 346980
rect 323170 346968 323176 346980
rect 321112 346940 323176 346968
rect 321112 346928 321118 346940
rect 323170 346928 323176 346940
rect 323228 346928 323234 346980
rect 80198 346860 80204 346912
rect 80256 346900 80262 346912
rect 87282 346900 87288 346912
rect 80256 346872 87288 346900
rect 80256 346860 80262 346872
rect 87282 346860 87288 346872
rect 87340 346860 87346 346912
rect 137422 346860 137428 346912
rect 137480 346900 137486 346912
rect 139630 346900 139636 346912
rect 137480 346872 139636 346900
rect 137480 346860 137486 346872
rect 139630 346860 139636 346872
rect 139688 346860 139694 346912
rect 174038 346860 174044 346912
rect 174096 346900 174102 346912
rect 182318 346900 182324 346912
rect 174096 346872 182324 346900
rect 174096 346860 174102 346872
rect 182318 346860 182324 346872
rect 182376 346860 182382 346912
rect 267878 346860 267884 346912
rect 267936 346900 267942 346912
rect 274870 346900 274876 346912
rect 267936 346872 274876 346900
rect 267936 346860 267942 346872
rect 274870 346860 274876 346872
rect 274928 346860 274934 346912
rect 79278 346792 79284 346844
rect 79336 346832 79342 346844
rect 87374 346832 87380 346844
rect 79336 346804 87380 346832
rect 79336 346792 79342 346804
rect 87374 346792 87380 346804
rect 87432 346792 87438 346844
rect 137606 346792 137612 346844
rect 137664 346832 137670 346844
rect 139722 346832 139728 346844
rect 137664 346804 139728 346832
rect 137664 346792 137670 346804
rect 139722 346792 139728 346804
rect 139780 346792 139786 346844
rect 173762 346792 173768 346844
rect 173820 346832 173826 346844
rect 182134 346832 182140 346844
rect 173820 346804 182140 346832
rect 173820 346792 173826 346804
rect 182134 346792 182140 346804
rect 182192 346792 182198 346844
rect 267418 346792 267424 346844
rect 267476 346832 267482 346844
rect 275054 346832 275060 346844
rect 267476 346804 275060 346832
rect 267476 346792 267482 346804
rect 275054 346792 275060 346804
rect 275112 346792 275118 346844
rect 321606 345704 321612 345756
rect 321664 345744 321670 345756
rect 326942 345744 326948 345756
rect 321664 345716 326948 345744
rect 321664 345704 321670 345716
rect 326942 345704 326948 345716
rect 327000 345704 327006 345756
rect 131810 345636 131816 345688
rect 131868 345676 131874 345688
rect 134110 345676 134116 345688
rect 131868 345648 134116 345676
rect 131868 345636 131874 345648
rect 134110 345636 134116 345648
rect 134168 345636 134174 345688
rect 172842 345636 172848 345688
rect 172900 345676 172906 345688
rect 181582 345676 181588 345688
rect 172900 345648 181588 345676
rect 172900 345636 172906 345648
rect 181582 345636 181588 345648
rect 181640 345636 181646 345688
rect 226294 345636 226300 345688
rect 226352 345676 226358 345688
rect 227950 345676 227956 345688
rect 226352 345648 227956 345676
rect 226352 345636 226358 345648
rect 227950 345636 227956 345648
rect 228008 345636 228014 345688
rect 79646 345568 79652 345620
rect 79704 345608 79710 345620
rect 87190 345608 87196 345620
rect 79704 345580 87196 345608
rect 79704 345568 79710 345580
rect 87190 345568 87196 345580
rect 87248 345568 87254 345620
rect 131902 345568 131908 345620
rect 131960 345608 131966 345620
rect 139630 345608 139636 345620
rect 131960 345580 139636 345608
rect 131960 345568 131966 345580
rect 139630 345568 139636 345580
rect 139688 345568 139694 345620
rect 172934 345568 172940 345620
rect 172992 345608 172998 345620
rect 182318 345608 182324 345620
rect 172992 345580 182324 345608
rect 172992 345568 172998 345580
rect 182318 345568 182324 345580
rect 182376 345568 182382 345620
rect 226386 345568 226392 345620
rect 226444 345608 226450 345620
rect 234574 345608 234580 345620
rect 226444 345580 234580 345608
rect 226444 345568 226450 345580
rect 234574 345568 234580 345580
rect 234632 345568 234638 345620
rect 270730 345568 270736 345620
rect 270788 345608 270794 345620
rect 274870 345608 274876 345620
rect 270788 345580 274876 345608
rect 270788 345568 270794 345580
rect 274870 345568 274876 345580
rect 274928 345568 274934 345620
rect 320502 345568 320508 345620
rect 320560 345608 320566 345620
rect 323262 345608 323268 345620
rect 320560 345580 323268 345608
rect 320560 345568 320566 345580
rect 323262 345568 323268 345580
rect 323320 345568 323326 345620
rect 228410 345500 228416 345552
rect 228468 345540 228474 345552
rect 233470 345540 233476 345552
rect 228468 345512 233476 345540
rect 228468 345500 228474 345512
rect 233470 345500 233476 345512
rect 233528 345500 233534 345552
rect 267878 345500 267884 345552
rect 267936 345540 267942 345552
rect 275146 345540 275152 345552
rect 267936 345512 275152 345540
rect 267936 345500 267942 345512
rect 275146 345500 275152 345512
rect 275204 345500 275210 345552
rect 323170 345500 323176 345552
rect 323228 345540 323234 345552
rect 328046 345540 328052 345552
rect 323228 345512 328052 345540
rect 323228 345500 323234 345512
rect 328046 345500 328052 345512
rect 328104 345500 328110 345552
rect 80198 344752 80204 344804
rect 80256 344792 80262 344804
rect 87098 344792 87104 344804
rect 80256 344764 87104 344792
rect 80256 344752 80262 344764
rect 87098 344752 87104 344764
rect 87156 344752 87162 344804
rect 172750 344752 172756 344804
rect 172808 344792 172814 344804
rect 180938 344792 180944 344804
rect 172808 344764 180944 344792
rect 172808 344752 172814 344764
rect 180938 344752 180944 344764
rect 180996 344752 181002 344804
rect 85810 344616 85816 344668
rect 85868 344656 85874 344668
rect 87374 344656 87380 344668
rect 85868 344628 87380 344656
rect 85868 344616 85874 344628
rect 87374 344616 87380 344628
rect 87432 344616 87438 344668
rect 320962 344480 320968 344532
rect 321020 344520 321026 344532
rect 323262 344520 323268 344532
rect 321020 344492 323268 344520
rect 321020 344480 321026 344492
rect 323262 344480 323268 344492
rect 323320 344480 323326 344532
rect 131810 344208 131816 344260
rect 131868 344248 131874 344260
rect 139814 344248 139820 344260
rect 131868 344220 139820 344248
rect 131868 344208 131874 344220
rect 139814 344208 139820 344220
rect 139872 344208 139878 344260
rect 226478 344208 226484 344260
rect 226536 344248 226542 344260
rect 234482 344248 234488 344260
rect 226536 344220 234488 344248
rect 226536 344208 226542 344220
rect 234482 344208 234488 344220
rect 234540 344208 234546 344260
rect 321606 344208 321612 344260
rect 321664 344248 321670 344260
rect 327402 344248 327408 344260
rect 321664 344220 327408 344248
rect 321664 344208 321670 344220
rect 327402 344208 327408 344220
rect 327460 344208 327466 344260
rect 132362 344140 132368 344192
rect 132420 344180 132426 344192
rect 139722 344180 139728 344192
rect 132420 344152 139728 344180
rect 132420 344140 132426 344152
rect 139722 344140 139728 344152
rect 139780 344140 139786 344192
rect 173118 344140 173124 344192
rect 173176 344180 173182 344192
rect 182318 344180 182324 344192
rect 173176 344152 182324 344180
rect 173176 344140 173182 344152
rect 182318 344140 182324 344152
rect 182376 344140 182382 344192
rect 226386 344140 226392 344192
rect 226444 344180 226450 344192
rect 234390 344180 234396 344192
rect 226444 344152 234396 344180
rect 226444 344140 226450 344152
rect 234390 344140 234396 344152
rect 234448 344140 234454 344192
rect 75969 344115 76027 344121
rect 75969 344081 75981 344115
rect 76015 344112 76027 344115
rect 76058 344112 76064 344124
rect 76015 344084 76064 344112
rect 76015 344081 76027 344084
rect 75969 344075 76027 344081
rect 76058 344072 76064 344084
rect 76116 344072 76122 344124
rect 76150 344072 76156 344124
rect 76208 344072 76214 344124
rect 227950 344072 227956 344124
rect 228008 344112 228014 344124
rect 233470 344112 233476 344124
rect 228008 344084 233476 344112
rect 228008 344072 228014 344084
rect 233470 344072 233476 344084
rect 233528 344072 233534 344124
rect 266682 344072 266688 344124
rect 266740 344112 266746 344124
rect 274962 344112 274968 344124
rect 266740 344084 274968 344112
rect 266740 344072 266746 344084
rect 274962 344072 274968 344084
rect 275020 344072 275026 344124
rect 323170 344072 323176 344124
rect 323228 344112 323234 344124
rect 328506 344112 328512 344124
rect 323228 344084 328512 344112
rect 323228 344072 323234 344084
rect 328506 344072 328512 344084
rect 328564 344072 328570 344124
rect 76168 343784 76196 344072
rect 76150 343732 76156 343784
rect 76208 343732 76214 343784
rect 321606 342848 321612 342900
rect 321664 342888 321670 342900
rect 327218 342888 327224 342900
rect 321664 342860 327224 342888
rect 321664 342848 321670 342860
rect 327218 342848 327224 342860
rect 327276 342848 327282 342900
rect 131810 342780 131816 342832
rect 131868 342820 131874 342832
rect 137514 342820 137520 342832
rect 131868 342792 137520 342820
rect 131868 342780 131874 342792
rect 137514 342780 137520 342792
rect 137572 342780 137578 342832
rect 173946 342780 173952 342832
rect 174004 342820 174010 342832
rect 181398 342820 181404 342832
rect 174004 342792 181404 342820
rect 174004 342780 174010 342792
rect 181398 342780 181404 342792
rect 181456 342780 181462 342832
rect 226386 342780 226392 342832
rect 226444 342820 226450 342832
rect 230526 342820 230532 342832
rect 226444 342792 230532 342820
rect 226444 342780 226450 342792
rect 230526 342780 230532 342792
rect 230584 342780 230590 342832
rect 80198 342712 80204 342764
rect 80256 342752 80262 342764
rect 88110 342752 88116 342764
rect 80256 342724 88116 342752
rect 80256 342712 80262 342724
rect 88110 342712 88116 342724
rect 88168 342712 88174 342764
rect 134110 342712 134116 342764
rect 134168 342752 134174 342764
rect 139630 342752 139636 342764
rect 134168 342724 139636 342752
rect 134168 342712 134174 342724
rect 139630 342712 139636 342724
rect 139688 342712 139694 342764
rect 172750 342712 172756 342764
rect 172808 342752 172814 342764
rect 180938 342752 180944 342764
rect 172808 342724 180944 342752
rect 172808 342712 172814 342724
rect 180938 342712 180944 342724
rect 180996 342712 181002 342764
rect 267602 342712 267608 342764
rect 267660 342752 267666 342764
rect 274870 342752 274876 342764
rect 267660 342724 274876 342752
rect 267660 342712 267666 342724
rect 274870 342712 274876 342724
rect 274928 342712 274934 342764
rect 323262 342712 323268 342764
rect 323320 342752 323326 342764
rect 328046 342752 328052 342764
rect 323320 342724 328052 342752
rect 323320 342712 323326 342724
rect 328046 342712 328052 342724
rect 328104 342712 328110 342764
rect 267878 342644 267884 342696
rect 267936 342684 267942 342696
rect 270730 342684 270736 342696
rect 267936 342656 270736 342684
rect 267936 342644 267942 342656
rect 270730 342644 270736 342656
rect 270788 342644 270794 342696
rect 80198 342100 80204 342152
rect 80256 342140 80262 342152
rect 85810 342140 85816 342152
rect 80256 342112 85816 342140
rect 80256 342100 80262 342112
rect 85810 342100 85816 342112
rect 85868 342100 85874 342152
rect 131902 341488 131908 341540
rect 131960 341528 131966 341540
rect 135398 341528 135404 341540
rect 131960 341500 135404 341528
rect 131960 341488 131966 341500
rect 135398 341488 135404 341500
rect 135456 341488 135462 341540
rect 173762 341488 173768 341540
rect 173820 341528 173826 341540
rect 182318 341528 182324 341540
rect 173820 341500 182324 341528
rect 173820 341488 173826 341500
rect 182318 341488 182324 341500
rect 182376 341488 182382 341540
rect 226478 341488 226484 341540
rect 226536 341528 226542 341540
rect 231998 341528 232004 341540
rect 226536 341500 232004 341528
rect 226536 341488 226542 341500
rect 231998 341488 232004 341500
rect 232056 341488 232062 341540
rect 321054 341488 321060 341540
rect 321112 341528 321118 341540
rect 327126 341528 327132 341540
rect 321112 341500 327132 341528
rect 321112 341488 321118 341500
rect 327126 341488 327132 341500
rect 327184 341488 327190 341540
rect 131810 341420 131816 341472
rect 131868 341460 131874 341472
rect 135306 341460 135312 341472
rect 131868 341432 135312 341460
rect 131868 341420 131874 341432
rect 135306 341420 135312 341432
rect 135364 341420 135370 341472
rect 174038 341420 174044 341472
rect 174096 341460 174102 341472
rect 181398 341460 181404 341472
rect 174096 341432 181404 341460
rect 174096 341420 174102 341432
rect 181398 341420 181404 341432
rect 181456 341420 181462 341472
rect 226386 341420 226392 341472
rect 226444 341460 226450 341472
rect 231814 341460 231820 341472
rect 226444 341432 231820 341460
rect 226444 341420 226450 341432
rect 231814 341420 231820 341432
rect 231872 341420 231878 341472
rect 321606 341420 321612 341472
rect 321664 341460 321670 341472
rect 327034 341460 327040 341472
rect 321664 341432 327040 341460
rect 321664 341420 321670 341432
rect 327034 341420 327040 341432
rect 327092 341420 327098 341472
rect 80198 341352 80204 341404
rect 80256 341392 80262 341404
rect 88478 341392 88484 341404
rect 80256 341364 88484 341392
rect 80256 341352 80262 341364
rect 88478 341352 88484 341364
rect 88536 341352 88542 341404
rect 267878 341352 267884 341404
rect 267936 341392 267942 341404
rect 275054 341392 275060 341404
rect 267936 341364 275060 341392
rect 267936 341352 267942 341364
rect 275054 341352 275060 341364
rect 275112 341352 275118 341404
rect 131810 340060 131816 340112
rect 131868 340100 131874 340112
rect 139538 340100 139544 340112
rect 131868 340072 139544 340100
rect 131868 340060 131874 340072
rect 139538 340060 139544 340072
rect 139596 340060 139602 340112
rect 173854 340060 173860 340112
rect 173912 340100 173918 340112
rect 181398 340100 181404 340112
rect 173912 340072 181404 340100
rect 173912 340060 173918 340072
rect 181398 340060 181404 340072
rect 181456 340060 181462 340112
rect 226386 340060 226392 340112
rect 226444 340100 226450 340112
rect 233562 340100 233568 340112
rect 226444 340072 233568 340100
rect 226444 340060 226450 340072
rect 233562 340060 233568 340072
rect 233620 340060 233626 340112
rect 272018 340060 272024 340112
rect 272076 340100 272082 340112
rect 274870 340100 274876 340112
rect 272076 340072 274876 340100
rect 272076 340060 272082 340072
rect 274870 340060 274876 340072
rect 274928 340060 274934 340112
rect 320594 340060 320600 340112
rect 320652 340100 320658 340112
rect 327862 340100 327868 340112
rect 320652 340072 327868 340100
rect 320652 340060 320658 340072
rect 327862 340060 327868 340072
rect 327920 340060 327926 340112
rect 374138 340060 374144 340112
rect 374196 340100 374202 340112
rect 429430 340100 429436 340112
rect 374196 340072 429436 340100
rect 374196 340060 374202 340072
rect 429430 340060 429436 340072
rect 429488 340060 429494 340112
rect 80198 339992 80204 340044
rect 80256 340032 80262 340044
rect 87282 340032 87288 340044
rect 80256 340004 87288 340032
rect 80256 339992 80262 340004
rect 87282 339992 87288 340004
rect 87340 339992 87346 340044
rect 137514 339992 137520 340044
rect 137572 340032 137578 340044
rect 139630 340032 139636 340044
rect 137572 340004 139636 340032
rect 137572 339992 137578 340004
rect 139630 339992 139636 340004
rect 139688 339992 139694 340044
rect 230526 339992 230532 340044
rect 230584 340032 230590 340044
rect 233470 340032 233476 340044
rect 230584 340004 233476 340032
rect 230584 339992 230590 340004
rect 233470 339992 233476 340004
rect 233528 339992 233534 340044
rect 267878 339992 267884 340044
rect 267936 340032 267942 340044
rect 275146 340032 275152 340044
rect 267936 340004 275152 340032
rect 267936 339992 267942 340004
rect 275146 339992 275152 340004
rect 275204 339992 275210 340044
rect 266961 339355 267019 339361
rect 266961 339321 266973 339355
rect 267007 339352 267019 339355
rect 267142 339352 267148 339364
rect 267007 339324 267148 339352
rect 267007 339321 267019 339324
rect 266961 339315 267019 339321
rect 267142 339312 267148 339324
rect 267200 339312 267206 339364
rect 320410 338768 320416 338820
rect 320468 338808 320474 338820
rect 326574 338808 326580 338820
rect 320468 338780 326580 338808
rect 320468 338768 320474 338780
rect 326574 338768 326580 338780
rect 326632 338768 326638 338820
rect 131810 338700 131816 338752
rect 131868 338740 131874 338752
rect 136134 338740 136140 338752
rect 131868 338712 136140 338740
rect 131868 338700 131874 338712
rect 136134 338700 136140 338712
rect 136192 338700 136198 338752
rect 226478 338700 226484 338752
rect 226536 338740 226542 338752
rect 231906 338740 231912 338752
rect 226536 338712 231912 338740
rect 226536 338700 226542 338712
rect 231906 338700 231912 338712
rect 231964 338700 231970 338752
rect 85074 338632 85080 338684
rect 85132 338672 85138 338684
rect 87466 338672 87472 338684
rect 85132 338644 87472 338672
rect 85132 338632 85138 338644
rect 87466 338632 87472 338644
rect 87524 338632 87530 338684
rect 131902 338632 131908 338684
rect 131960 338672 131966 338684
rect 139630 338672 139636 338684
rect 131960 338644 139636 338672
rect 131960 338632 131966 338644
rect 139630 338632 139636 338644
rect 139688 338632 139694 338684
rect 173486 338632 173492 338684
rect 173544 338672 173550 338684
rect 181582 338672 181588 338684
rect 173544 338644 181588 338672
rect 173544 338632 173550 338644
rect 181582 338632 181588 338644
rect 181640 338632 181646 338684
rect 226386 338632 226392 338684
rect 226444 338672 226450 338684
rect 234114 338672 234120 338684
rect 226444 338644 234120 338672
rect 226444 338632 226450 338644
rect 234114 338632 234120 338644
rect 234172 338632 234178 338684
rect 267786 338632 267792 338684
rect 267844 338672 267850 338684
rect 274870 338672 274876 338684
rect 267844 338644 274876 338672
rect 267844 338632 267850 338644
rect 274870 338632 274876 338644
rect 274928 338632 274934 338684
rect 320502 338632 320508 338684
rect 320560 338672 320566 338684
rect 327218 338672 327224 338684
rect 320560 338644 327224 338672
rect 320560 338632 320566 338644
rect 327218 338632 327224 338644
rect 327276 338632 327282 338684
rect 80198 338564 80204 338616
rect 80256 338604 80262 338616
rect 87558 338604 87564 338616
rect 80256 338576 87564 338604
rect 80256 338564 80262 338576
rect 87558 338564 87564 338576
rect 87616 338564 87622 338616
rect 135398 338564 135404 338616
rect 135456 338604 135462 338616
rect 139722 338604 139728 338616
rect 135456 338576 139728 338604
rect 135456 338564 135462 338576
rect 139722 338564 139728 338576
rect 139780 338564 139786 338616
rect 231998 338564 232004 338616
rect 232056 338604 232062 338616
rect 233470 338604 233476 338616
rect 232056 338576 233476 338604
rect 232056 338564 232062 338576
rect 233470 338564 233476 338576
rect 233528 338564 233534 338616
rect 267510 338564 267516 338616
rect 267568 338604 267574 338616
rect 274962 338604 274968 338616
rect 267568 338576 274968 338604
rect 267568 338564 267574 338576
rect 274962 338564 274968 338576
rect 275020 338564 275026 338616
rect 80106 338496 80112 338548
rect 80164 338536 80170 338548
rect 87190 338536 87196 338548
rect 80164 338508 87196 338536
rect 80164 338496 80170 338508
rect 87190 338496 87196 338508
rect 87248 338496 87254 338548
rect 135306 338496 135312 338548
rect 135364 338536 135370 338548
rect 139814 338536 139820 338548
rect 135364 338508 139820 338536
rect 135364 338496 135370 338508
rect 139814 338496 139820 338508
rect 139872 338496 139878 338548
rect 231814 338496 231820 338548
rect 231872 338536 231878 338548
rect 233654 338536 233660 338548
rect 231872 338508 233660 338536
rect 231872 338496 231878 338508
rect 233654 338496 233660 338508
rect 233712 338496 233718 338548
rect 267878 338496 267884 338548
rect 267936 338536 267942 338548
rect 275238 338536 275244 338548
rect 267936 338508 275244 338536
rect 267936 338496 267942 338508
rect 275238 338496 275244 338508
rect 275296 338496 275302 338548
rect 226386 337612 226392 337664
rect 226444 337652 226450 337664
rect 231538 337652 231544 337664
rect 226444 337624 231544 337652
rect 226444 337612 226450 337624
rect 231538 337612 231544 337624
rect 231596 337612 231602 337664
rect 85166 337272 85172 337324
rect 85224 337312 85230 337324
rect 87190 337312 87196 337324
rect 85224 337284 87196 337312
rect 85224 337272 85230 337284
rect 87190 337272 87196 337284
rect 87248 337272 87254 337324
rect 131810 337272 131816 337324
rect 131868 337312 131874 337324
rect 136226 337312 136232 337324
rect 131868 337284 136232 337312
rect 131868 337272 131874 337284
rect 136226 337272 136232 337284
rect 136284 337272 136290 337324
rect 173670 337272 173676 337324
rect 173728 337312 173734 337324
rect 181766 337312 181772 337324
rect 173728 337284 181772 337312
rect 173728 337272 173734 337284
rect 181766 337272 181772 337284
rect 181824 337272 181830 337324
rect 270822 337272 270828 337324
rect 270880 337312 270886 337324
rect 274870 337312 274876 337324
rect 270880 337284 274876 337312
rect 270880 337272 270886 337284
rect 274870 337272 274876 337284
rect 274928 337272 274934 337324
rect 320410 337272 320416 337324
rect 320468 337312 320474 337324
rect 326758 337312 326764 337324
rect 320468 337284 326764 337312
rect 320468 337272 320474 337284
rect 326758 337272 326764 337284
rect 326816 337272 326822 337324
rect 79830 337204 79836 337256
rect 79888 337244 79894 337256
rect 87374 337244 87380 337256
rect 79888 337216 87380 337244
rect 79888 337204 79894 337216
rect 87374 337204 87380 337216
rect 87432 337204 87438 337256
rect 267326 337204 267332 337256
rect 267384 337244 267390 337256
rect 272018 337244 272024 337256
rect 267384 337216 272024 337244
rect 267384 337204 267390 337216
rect 272018 337204 272024 337216
rect 272076 337204 272082 337256
rect 320410 336048 320416 336100
rect 320468 336088 320474 336100
rect 327310 336088 327316 336100
rect 320468 336060 327316 336088
rect 320468 336048 320474 336060
rect 327310 336048 327316 336060
rect 327368 336048 327374 336100
rect 131902 335980 131908 336032
rect 131960 336020 131966 336032
rect 137606 336020 137612 336032
rect 131960 335992 137612 336020
rect 131960 335980 131966 335992
rect 137606 335980 137612 335992
rect 137664 335980 137670 336032
rect 172842 335980 172848 336032
rect 172900 336020 172906 336032
rect 181582 336020 181588 336032
rect 172900 335992 181588 336020
rect 172900 335980 172906 335992
rect 181582 335980 181588 335992
rect 181640 335980 181646 336032
rect 270730 335980 270736 336032
rect 270788 336020 270794 336032
rect 274962 336020 274968 336032
rect 270788 335992 274968 336020
rect 270788 335980 270794 335992
rect 274962 335980 274968 335992
rect 275020 335980 275026 336032
rect 85810 335912 85816 335964
rect 85868 335952 85874 335964
rect 87190 335952 87196 335964
rect 85868 335924 87196 335952
rect 85868 335912 85874 335924
rect 87190 335912 87196 335924
rect 87248 335912 87254 335964
rect 131810 335912 131816 335964
rect 131868 335952 131874 335964
rect 139814 335952 139820 335964
rect 131868 335924 139820 335952
rect 131868 335912 131874 335924
rect 139814 335912 139820 335924
rect 139872 335912 139878 335964
rect 172934 335912 172940 335964
rect 172992 335952 172998 335964
rect 181766 335952 181772 335964
rect 172992 335924 181772 335952
rect 172992 335912 172998 335924
rect 181766 335912 181772 335924
rect 181824 335912 181830 335964
rect 226386 335912 226392 335964
rect 226444 335952 226450 335964
rect 230710 335952 230716 335964
rect 226444 335924 230716 335952
rect 226444 335912 226450 335924
rect 230710 335912 230716 335924
rect 230768 335912 230774 335964
rect 266774 335912 266780 335964
rect 266832 335952 266838 335964
rect 274870 335952 274876 335964
rect 266832 335924 274876 335952
rect 266832 335912 266838 335924
rect 274870 335912 274876 335924
rect 274928 335912 274934 335964
rect 80198 335844 80204 335896
rect 80256 335884 80262 335896
rect 87282 335884 87288 335896
rect 80256 335856 87288 335884
rect 80256 335844 80262 335856
rect 87282 335844 87288 335856
rect 87340 335844 87346 335896
rect 231906 335844 231912 335896
rect 231964 335884 231970 335896
rect 233470 335884 233476 335896
rect 231964 335856 233476 335884
rect 231964 335844 231970 335856
rect 233470 335844 233476 335856
rect 233528 335844 233534 335896
rect 267878 335844 267884 335896
rect 267936 335884 267942 335896
rect 275054 335884 275060 335896
rect 267936 335856 275060 335884
rect 267936 335844 267942 335856
rect 275054 335844 275060 335856
rect 275112 335844 275118 335896
rect 75417 334799 75475 334805
rect 75417 334765 75429 334799
rect 75463 334796 75475 334799
rect 75966 334796 75972 334808
rect 75463 334768 75972 334796
rect 75463 334765 75475 334768
rect 75417 334759 75475 334765
rect 75966 334756 75972 334768
rect 76024 334756 76030 334808
rect 75509 334731 75567 334737
rect 75509 334697 75521 334731
rect 75555 334728 75567 334731
rect 75874 334728 75880 334740
rect 75555 334700 75880 334728
rect 75555 334697 75567 334700
rect 75509 334691 75567 334697
rect 75874 334688 75880 334700
rect 75932 334688 75938 334740
rect 76058 334688 76064 334740
rect 76116 334688 76122 334740
rect 76076 334536 76104 334688
rect 75966 334524 75972 334536
rect 75927 334496 75972 334524
rect 75966 334484 75972 334496
rect 76024 334484 76030 334536
rect 76058 334484 76064 334536
rect 76116 334484 76122 334536
rect 108258 334456 108264 334468
rect 75800 334428 108264 334456
rect 75800 334320 75828 334428
rect 108258 334416 108264 334428
rect 108316 334456 108322 334468
rect 131626 334456 131632 334468
rect 108316 334428 131632 334456
rect 108316 334416 108322 334428
rect 131626 334416 131632 334428
rect 131684 334416 131690 334468
rect 136134 334416 136140 334468
rect 136192 334456 136198 334468
rect 139630 334456 139636 334468
rect 136192 334428 139636 334456
rect 136192 334416 136198 334428
rect 139630 334416 139636 334428
rect 139688 334416 139694 334468
rect 202466 334416 202472 334468
rect 202524 334456 202530 334468
rect 225374 334456 225380 334468
rect 202524 334428 225380 334456
rect 202524 334416 202530 334428
rect 225374 334416 225380 334428
rect 225432 334416 225438 334468
rect 267326 334416 267332 334468
rect 267384 334456 267390 334468
rect 270822 334456 270828 334468
rect 267384 334428 270828 334456
rect 267384 334416 267390 334428
rect 270822 334416 270828 334428
rect 270880 334416 270886 334468
rect 306242 334416 306248 334468
rect 306300 334456 306306 334468
rect 319122 334456 319128 334468
rect 306300 334428 319128 334456
rect 306300 334416 306306 334428
rect 319122 334416 319128 334428
rect 319180 334456 319186 334468
rect 319674 334456 319680 334468
rect 319180 334428 319680 334456
rect 319180 334416 319186 334428
rect 319674 334416 319680 334428
rect 319732 334416 319738 334468
rect 75874 334348 75880 334400
rect 75932 334388 75938 334400
rect 104854 334388 104860 334400
rect 75932 334360 104860 334388
rect 75932 334348 75938 334360
rect 104854 334348 104860 334360
rect 104912 334388 104918 334400
rect 131718 334388 131724 334400
rect 104912 334360 131724 334388
rect 104912 334348 104918 334360
rect 131718 334348 131724 334360
rect 131776 334348 131782 334400
rect 174038 334348 174044 334400
rect 174096 334388 174102 334400
rect 180294 334388 180300 334400
rect 174096 334360 180300 334388
rect 174096 334348 174102 334360
rect 180294 334348 180300 334360
rect 180352 334348 180358 334400
rect 212310 334348 212316 334400
rect 212368 334388 212374 334400
rect 225190 334388 225196 334400
rect 212368 334360 225196 334388
rect 212368 334348 212374 334360
rect 225190 334348 225196 334360
rect 225248 334348 225254 334400
rect 75966 334320 75972 334332
rect 75800 334292 75972 334320
rect 75966 334280 75972 334292
rect 76024 334280 76030 334332
rect 76978 334280 76984 334332
rect 77036 334320 77042 334332
rect 98230 334320 98236 334332
rect 77036 334292 98236 334320
rect 77036 334280 77042 334292
rect 98230 334280 98236 334292
rect 98288 334280 98294 334332
rect 111386 334280 111392 334332
rect 111444 334320 111450 334332
rect 131534 334320 131540 334332
rect 111444 334292 131540 334320
rect 111444 334280 111450 334292
rect 131534 334280 131540 334292
rect 131592 334280 131598 334332
rect 114790 334212 114796 334264
rect 114848 334252 114854 334264
rect 131442 334252 131448 334264
rect 114848 334224 131448 334252
rect 114848 334212 114854 334224
rect 131442 334212 131448 334224
rect 131500 334212 131506 334264
rect 136226 334212 136232 334264
rect 136284 334252 136290 334264
rect 139630 334252 139636 334264
rect 136284 334224 139636 334252
rect 136284 334212 136290 334224
rect 139630 334212 139636 334224
rect 139688 334212 139694 334264
rect 118194 334144 118200 334196
rect 118252 334184 118258 334196
rect 131350 334184 131356 334196
rect 118252 334156 131356 334184
rect 118252 334144 118258 334156
rect 131350 334144 131356 334156
rect 131408 334144 131414 334196
rect 131718 334144 131724 334196
rect 131776 334184 131782 334196
rect 136870 334184 136876 334196
rect 131776 334156 136876 334184
rect 131776 334144 131782 334156
rect 136870 334144 136876 334156
rect 136928 334144 136934 334196
rect 131534 334076 131540 334128
rect 131592 334116 131598 334128
rect 137054 334116 137060 334128
rect 131592 334088 137060 334116
rect 131592 334076 131598 334088
rect 137054 334076 137060 334088
rect 137112 334076 137118 334128
rect 231538 334076 231544 334128
rect 231596 334116 231602 334128
rect 234298 334116 234304 334128
rect 231596 334088 234304 334116
rect 231596 334076 231602 334088
rect 234298 334076 234304 334088
rect 234356 334076 234362 334128
rect 80198 334008 80204 334060
rect 80256 334048 80262 334060
rect 85166 334048 85172 334060
rect 80256 334020 85172 334048
rect 80256 334008 80262 334020
rect 85166 334008 85172 334020
rect 85224 334008 85230 334060
rect 116078 334008 116084 334060
rect 116136 334048 116142 334060
rect 127854 334048 127860 334060
rect 116136 334020 127860 334048
rect 116136 334008 116142 334020
rect 127854 334008 127860 334020
rect 127912 334008 127918 334060
rect 131626 334008 131632 334060
rect 131684 334048 131690 334060
rect 137330 334048 137336 334060
rect 131684 334020 137336 334048
rect 131684 334008 131690 334020
rect 137330 334008 137336 334020
rect 137388 334008 137394 334060
rect 103658 333940 103664 333992
rect 103716 333980 103722 333992
rect 124542 333980 124548 333992
rect 103716 333952 124548 333980
rect 103716 333940 103722 333952
rect 124542 333940 124548 333952
rect 124600 333940 124606 333992
rect 131442 333940 131448 333992
rect 131500 333980 131506 333992
rect 137514 333980 137520 333992
rect 131500 333952 137520 333980
rect 131500 333940 131506 333952
rect 137514 333940 137520 333952
rect 137572 333940 137578 333992
rect 211298 333940 211304 333992
rect 211356 333980 211362 333992
rect 221878 333980 221884 333992
rect 211356 333952 221884 333980
rect 211356 333940 211362 333952
rect 221878 333940 221884 333952
rect 221936 333940 221942 333992
rect 305138 333940 305144 333992
rect 305196 333980 305202 333992
rect 316178 333980 316184 333992
rect 305196 333952 316184 333980
rect 305196 333940 305202 333952
rect 316178 333940 316184 333952
rect 316236 333940 316242 333992
rect 80106 333872 80112 333924
rect 80164 333912 80170 333924
rect 85074 333912 85080 333924
rect 80164 333884 85080 333912
rect 80164 333872 80170 333884
rect 85074 333872 85080 333884
rect 85132 333872 85138 333924
rect 91238 333872 91244 333924
rect 91296 333912 91302 333924
rect 121230 333912 121236 333924
rect 91296 333884 121236 333912
rect 91296 333872 91302 333884
rect 121230 333872 121236 333884
rect 121288 333872 121294 333924
rect 131350 333872 131356 333924
rect 131408 333912 131414 333924
rect 137698 333912 137704 333924
rect 131408 333884 137704 333912
rect 131408 333872 131414 333884
rect 137698 333872 137704 333884
rect 137756 333872 137762 333924
rect 197498 333872 197504 333924
rect 197556 333912 197562 333924
rect 218566 333912 218572 333924
rect 197556 333884 218572 333912
rect 197556 333872 197562 333884
rect 218566 333872 218572 333884
rect 218624 333872 218630 333924
rect 292718 333872 292724 333924
rect 292776 333912 292782 333924
rect 312866 333912 312872 333924
rect 292776 333884 312872 333912
rect 292776 333872 292782 333884
rect 312866 333872 312872 333884
rect 312924 333872 312930 333924
rect 98230 333804 98236 333856
rect 98288 333844 98294 333856
rect 137790 333844 137796 333856
rect 98288 333816 137796 333844
rect 98288 333804 98294 333816
rect 137790 333804 137796 333816
rect 137848 333804 137854 333856
rect 185078 333804 185084 333856
rect 185136 333844 185142 333856
rect 215622 333844 215628 333856
rect 185136 333816 215628 333844
rect 185136 333804 185142 333816
rect 215622 333804 215628 333816
rect 215680 333804 215686 333856
rect 280298 333804 280304 333856
rect 280356 333844 280362 333856
rect 309554 333844 309560 333856
rect 280356 333816 309560 333844
rect 280356 333804 280362 333816
rect 309554 333804 309560 333816
rect 309612 333804 309618 333856
rect 91882 333736 91888 333788
rect 91940 333776 91946 333788
rect 134846 333776 134852 333788
rect 91940 333748 134852 333776
rect 91940 333736 91946 333748
rect 134846 333736 134852 333748
rect 134904 333736 134910 333788
rect 185906 333736 185912 333788
rect 185964 333776 185970 333788
rect 228686 333776 228692 333788
rect 185964 333748 228692 333776
rect 185964 333736 185970 333748
rect 228686 333736 228692 333748
rect 228744 333736 228750 333788
rect 279562 333736 279568 333788
rect 279620 333776 279626 333788
rect 323814 333776 323820 333788
rect 279620 333748 323820 333776
rect 279620 333736 279626 333748
rect 323814 333736 323820 333748
rect 323872 333736 323878 333788
rect 225190 333532 225196 333584
rect 225248 333572 225254 333584
rect 230986 333572 230992 333584
rect 225248 333544 230992 333572
rect 225248 333532 225254 333544
rect 230986 333532 230992 333544
rect 231044 333572 231050 333584
rect 231814 333572 231820 333584
rect 231044 333544 231820 333572
rect 231044 333532 231050 333544
rect 231814 333532 231820 333544
rect 231872 333532 231878 333584
rect 225374 333124 225380 333176
rect 225432 333164 225438 333176
rect 231354 333164 231360 333176
rect 225432 333136 231360 333164
rect 225432 333124 225438 333136
rect 231354 333124 231360 333136
rect 231412 333124 231418 333176
rect 319674 333124 319680 333176
rect 319732 333164 319738 333176
rect 325378 333164 325384 333176
rect 319732 333136 325384 333164
rect 319732 333124 319738 333136
rect 325378 333124 325384 333136
rect 325436 333124 325442 333176
rect 80198 333056 80204 333108
rect 80256 333096 80262 333108
rect 87558 333096 87564 333108
rect 80256 333068 87564 333096
rect 80256 333056 80262 333068
rect 87558 333056 87564 333068
rect 87616 333056 87622 333108
rect 137606 333056 137612 333108
rect 137664 333096 137670 333108
rect 139630 333096 139636 333108
rect 137664 333068 139636 333096
rect 137664 333056 137670 333068
rect 139630 333056 139636 333068
rect 139688 333056 139694 333108
rect 230710 333056 230716 333108
rect 230768 333096 230774 333108
rect 233930 333096 233936 333108
rect 230768 333068 233936 333096
rect 230768 333056 230774 333068
rect 233930 333056 233936 333068
rect 233988 333056 233994 333108
rect 267142 333056 267148 333108
rect 267200 333096 267206 333108
rect 270730 333096 270736 333108
rect 267200 333068 270736 333096
rect 267200 333056 267206 333068
rect 270730 333056 270736 333068
rect 270788 333056 270794 333108
rect 198786 332920 198792 332972
rect 198844 332960 198850 332972
rect 228778 332960 228784 332972
rect 198844 332932 228784 332960
rect 198844 332920 198850 332932
rect 228778 332920 228784 332932
rect 228836 332960 228842 332972
rect 231446 332960 231452 332972
rect 228836 332932 231452 332960
rect 228836 332920 228842 332932
rect 231446 332920 231452 332932
rect 231504 332920 231510 332972
rect 319858 331764 319864 331816
rect 319916 331804 319922 331816
rect 325194 331804 325200 331816
rect 319916 331776 325200 331804
rect 319916 331764 319922 331776
rect 325194 331764 325200 331776
rect 325252 331764 325258 331816
rect 76886 331696 76892 331748
rect 76944 331736 76950 331748
rect 118194 331736 118200 331748
rect 76944 331708 118200 331736
rect 76944 331696 76950 331708
rect 118194 331696 118200 331708
rect 118252 331696 118258 331748
rect 226570 331696 226576 331748
rect 226628 331736 226634 331748
rect 233470 331736 233476 331748
rect 226628 331708 233476 331736
rect 226628 331696 226634 331708
rect 233470 331696 233476 331708
rect 233528 331696 233534 331748
rect 319122 331736 319128 331748
rect 312056 331708 319128 331736
rect 75509 331671 75567 331677
rect 75509 331637 75521 331671
rect 75555 331668 75567 331671
rect 114790 331668 114796 331680
rect 75555 331640 114796 331668
rect 75555 331637 75567 331640
rect 75509 331631 75567 331637
rect 114790 331628 114796 331640
rect 114848 331628 114854 331680
rect 75417 331603 75475 331609
rect 75417 331569 75429 331603
rect 75463 331600 75475 331603
rect 111386 331600 111392 331612
rect 75463 331572 111392 331600
rect 75463 331569 75475 331572
rect 75417 331563 75475 331569
rect 111386 331560 111392 331572
rect 111444 331560 111450 331612
rect 309281 331603 309339 331609
rect 309281 331569 309293 331603
rect 309327 331600 309339 331603
rect 312056 331600 312084 331708
rect 319122 331696 319128 331708
rect 319180 331696 319186 331748
rect 320502 331696 320508 331748
rect 320560 331736 320566 331748
rect 328506 331736 328512 331748
rect 320560 331708 328512 331736
rect 320560 331696 320566 331708
rect 328506 331696 328512 331708
rect 328564 331696 328570 331748
rect 309327 331572 312084 331600
rect 309327 331569 309339 331572
rect 309281 331563 309339 331569
rect 299526 331492 299532 331544
rect 299584 331532 299590 331544
rect 299713 331535 299771 331541
rect 299713 331532 299725 331535
rect 299584 331504 299725 331532
rect 299584 331492 299590 331504
rect 299713 331501 299725 331504
rect 299759 331501 299771 331535
rect 299713 331495 299771 331501
rect 299713 331399 299771 331405
rect 299713 331365 299725 331399
rect 299759 331396 299771 331399
rect 309281 331399 309339 331405
rect 309281 331396 309293 331399
rect 299759 331368 309293 331396
rect 299759 331365 299771 331368
rect 299713 331359 299771 331365
rect 309281 331365 309293 331368
rect 309327 331365 309339 331399
rect 309281 331359 309339 331365
rect 80198 330744 80204 330796
rect 80256 330784 80262 330796
rect 85810 330784 85816 330796
rect 80256 330756 85816 330784
rect 80256 330744 80262 330756
rect 85810 330744 85816 330756
rect 85868 330744 85874 330796
rect 225282 330608 225288 330660
rect 225340 330648 225346 330660
rect 231722 330648 231728 330660
rect 225340 330620 231728 330648
rect 225340 330608 225346 330620
rect 231722 330608 231728 330620
rect 231780 330608 231786 330660
rect 319674 330472 319680 330524
rect 319732 330512 319738 330524
rect 325746 330512 325752 330524
rect 319732 330484 325752 330512
rect 319732 330472 319738 330484
rect 325746 330472 325752 330484
rect 325804 330472 325810 330524
rect 319122 330404 319128 330456
rect 319180 330444 319186 330456
rect 325286 330444 325292 330456
rect 319180 330416 325292 330444
rect 319180 330404 319186 330416
rect 325286 330404 325292 330416
rect 325344 330404 325350 330456
rect 75506 330172 75512 330184
rect 75467 330144 75512 330172
rect 75506 330132 75512 330144
rect 75564 330132 75570 330184
rect 75414 330104 75420 330116
rect 75375 330076 75420 330104
rect 75414 330064 75420 330076
rect 75472 330064 75478 330116
rect 290053 329359 290111 329365
rect 290053 329325 290065 329359
rect 290099 329356 290111 329359
rect 299621 329359 299679 329365
rect 299621 329356 299633 329359
rect 290099 329328 299633 329356
rect 290099 329325 290111 329328
rect 290053 329319 290111 329325
rect 299621 329325 299633 329328
rect 299667 329325 299679 329359
rect 299621 329319 299679 329325
rect 96853 329291 96911 329297
rect 96853 329257 96865 329291
rect 96899 329288 96911 329291
rect 106421 329291 106479 329297
rect 106421 329288 106433 329291
rect 96899 329260 106433 329288
rect 96899 329257 96911 329260
rect 96853 329251 96911 329257
rect 106421 329257 106433 329260
rect 106467 329257 106479 329291
rect 106421 329251 106479 329257
rect 128498 329220 128504 329232
rect 128332 329192 128504 329220
rect 87193 329155 87251 329161
rect 87193 329121 87205 329155
rect 87239 329152 87251 329155
rect 96853 329155 96911 329161
rect 96853 329152 96865 329155
rect 87239 329124 96865 329152
rect 87239 329121 87251 329124
rect 87193 329115 87251 329121
rect 96853 329121 96865 329124
rect 96899 329121 96911 329155
rect 96853 329115 96911 329121
rect 106421 329087 106479 329093
rect 106421 329053 106433 329087
rect 106467 329084 106479 329087
rect 106467 329056 109132 329084
rect 106467 329053 106479 329056
rect 106421 329047 106479 329053
rect 82314 328976 82320 329028
rect 82372 329016 82378 329028
rect 87193 329019 87251 329025
rect 87193 329016 87205 329019
rect 82372 328988 87205 329016
rect 82372 328976 82378 328988
rect 87193 328985 87205 328988
rect 87239 328985 87251 329019
rect 109104 329016 109132 329056
rect 109181 329019 109239 329025
rect 109181 329016 109193 329019
rect 109104 328988 109193 329016
rect 87193 328979 87251 328985
rect 109181 328985 109193 328988
rect 109227 328985 109239 329019
rect 109181 328979 109239 328985
rect 109365 329019 109423 329025
rect 109365 328985 109377 329019
rect 109411 329016 109423 329019
rect 116173 329019 116231 329025
rect 116173 329016 116185 329019
rect 109411 328988 116185 329016
rect 109411 328985 109423 328988
rect 109365 328979 109423 328985
rect 116173 328985 116185 328988
rect 116219 328985 116231 329019
rect 116173 328979 116231 328985
rect 119393 329019 119451 329025
rect 119393 328985 119405 329019
rect 119439 329016 119451 329019
rect 128332 329016 128360 329192
rect 128498 329180 128504 329192
rect 128556 329220 128562 329232
rect 140550 329220 140556 329232
rect 128556 329192 140556 329220
rect 128556 329180 128562 329192
rect 140550 329180 140556 329192
rect 140608 329180 140614 329232
rect 219673 329223 219731 329229
rect 219673 329189 219685 329223
rect 219719 329220 219731 329223
rect 222522 329220 222528 329232
rect 219719 329192 222528 329220
rect 219719 329189 219731 329192
rect 219673 329183 219731 329189
rect 222522 329180 222528 329192
rect 222580 329220 222586 329232
rect 233470 329220 233476 329232
rect 222580 329192 233476 329220
rect 222580 329180 222586 329192
rect 233470 329180 233476 329192
rect 233528 329180 233534 329232
rect 283061 329223 283119 329229
rect 283061 329220 283073 329223
rect 280408 329192 283073 329220
rect 267878 329112 267884 329164
rect 267936 329152 267942 329164
rect 280408 329152 280436 329192
rect 283061 329189 283073 329192
rect 283107 329189 283119 329223
rect 283061 329183 283119 329189
rect 283245 329223 283303 329229
rect 283245 329189 283257 329223
rect 283291 329220 283303 329223
rect 290053 329223 290111 329229
rect 290053 329220 290065 329223
rect 283291 329192 290065 329220
rect 283291 329189 283303 329192
rect 283245 329183 283303 329189
rect 290053 329189 290065 329192
rect 290099 329189 290111 329223
rect 290053 329183 290111 329189
rect 319033 329223 319091 329229
rect 319033 329189 319045 329223
rect 319079 329220 319091 329223
rect 319582 329220 319588 329232
rect 319079 329192 319588 329220
rect 319079 329189 319091 329192
rect 319033 329183 319091 329189
rect 319582 329180 319588 329192
rect 319640 329180 319646 329232
rect 267936 329124 280436 329152
rect 267936 329112 267942 329124
rect 173394 329044 173400 329096
rect 173452 329084 173458 329096
rect 186369 329087 186427 329093
rect 186369 329084 186381 329087
rect 173452 329056 186381 329084
rect 173452 329044 173458 329056
rect 186369 329053 186381 329056
rect 186415 329053 186427 329087
rect 186369 329047 186427 329053
rect 186553 329087 186611 329093
rect 186553 329053 186565 329087
rect 186599 329084 186611 329087
rect 203021 329087 203079 329093
rect 186599 329056 186780 329084
rect 186599 329053 186611 329056
rect 186553 329047 186611 329053
rect 119439 328988 128360 329016
rect 119439 328985 119451 328988
rect 119393 328979 119451 328985
rect 137698 328976 137704 329028
rect 137756 329016 137762 329028
rect 137882 329016 137888 329028
rect 137756 328988 137888 329016
rect 137756 328976 137762 328988
rect 137882 328976 137888 328988
rect 137940 329016 137946 329028
rect 161710 329016 161716 329028
rect 137940 328988 161716 329016
rect 137940 328976 137946 328988
rect 161710 328976 161716 328988
rect 161768 328976 161774 329028
rect 186752 329016 186780 329056
rect 203021 329053 203033 329087
rect 203067 329084 203079 329087
rect 205689 329087 205747 329093
rect 205689 329084 205701 329087
rect 203067 329056 205701 329084
rect 203067 329053 203079 329056
rect 203021 329047 203079 329053
rect 205689 329053 205701 329056
rect 205735 329053 205747 329087
rect 205689 329047 205747 329053
rect 205965 329087 206023 329093
rect 205965 329053 205977 329087
rect 206011 329084 206023 329087
rect 316546 329084 316552 329096
rect 206011 329056 215484 329084
rect 206011 329053 206023 329056
rect 205965 329047 206023 329053
rect 193453 329019 193511 329025
rect 193453 329016 193465 329019
rect 186752 328988 193465 329016
rect 193453 328985 193465 328988
rect 193499 328985 193511 329019
rect 215456 329016 215484 329056
rect 302488 329056 316552 329084
rect 219673 329019 219731 329025
rect 219673 329016 219685 329019
rect 215456 328988 219685 329016
rect 193453 328979 193511 328985
rect 219673 328985 219685 328988
rect 219719 328985 219731 329019
rect 219673 328979 219731 328985
rect 231354 328976 231360 329028
rect 231412 329016 231418 329028
rect 231722 329016 231728 329028
rect 231412 328988 231728 329016
rect 231412 328976 231418 328988
rect 231722 328976 231728 328988
rect 231780 329016 231786 329028
rect 253710 329016 253716 329028
rect 231780 328988 253716 329016
rect 231780 328976 231786 328988
rect 253710 328976 253716 328988
rect 253768 329016 253774 329028
rect 299526 329016 299532 329028
rect 253768 328988 299532 329016
rect 253768 328976 253774 328988
rect 299526 328976 299532 328988
rect 299584 328976 299590 329028
rect 299621 329019 299679 329025
rect 299621 328985 299633 329019
rect 299667 329016 299679 329019
rect 302488 329016 302516 329056
rect 316546 329044 316552 329056
rect 316604 329084 316610 329096
rect 319033 329087 319091 329093
rect 319033 329084 319045 329087
rect 316604 329056 319045 329084
rect 316604 329044 316610 329056
rect 319033 329053 319045 329056
rect 319079 329053 319091 329087
rect 319033 329047 319091 329053
rect 299667 328988 302516 329016
rect 299667 328985 299679 328988
rect 299621 328979 299679 328985
rect 209274 328908 209280 328960
rect 209332 328948 209338 328960
rect 227214 328948 227220 328960
rect 209332 328920 227220 328948
rect 209332 328908 209338 328920
rect 227214 328908 227220 328920
rect 227272 328948 227278 328960
rect 231446 328948 231452 328960
rect 227272 328920 231452 328948
rect 227272 328908 227278 328920
rect 231446 328908 231452 328920
rect 231504 328908 231510 328960
rect 265305 328951 265363 328957
rect 265305 328917 265317 328951
rect 265351 328948 265363 328951
rect 266961 328951 267019 328957
rect 266961 328948 266973 328951
rect 265351 328920 266973 328948
rect 265351 328917 265363 328920
rect 265305 328911 265363 328917
rect 266961 328917 266973 328920
rect 267007 328948 267019 328951
rect 285910 328948 285916 328960
rect 267007 328920 285916 328948
rect 267007 328917 267019 328920
rect 266961 328911 267019 328917
rect 285910 328908 285916 328920
rect 285968 328908 285974 328960
rect 303114 328908 303120 328960
rect 303172 328948 303178 328960
rect 319030 328948 319036 328960
rect 303172 328920 319036 328948
rect 303172 328908 303178 328920
rect 319030 328908 319036 328920
rect 319088 328948 319094 328960
rect 324734 328948 324740 328960
rect 319088 328920 324740 328948
rect 319088 328908 319094 328920
rect 324734 328908 324740 328920
rect 324792 328908 324798 328960
rect 116173 328883 116231 328889
rect 116173 328849 116185 328883
rect 116219 328880 116231 328883
rect 119393 328883 119451 328889
rect 119393 328880 119405 328883
rect 116219 328852 119405 328880
rect 116219 328849 116231 328852
rect 116173 328843 116231 328849
rect 119393 328849 119405 328852
rect 119439 328849 119451 328883
rect 119393 328843 119451 328849
rect 193453 328883 193511 328889
rect 193453 328849 193465 328883
rect 193499 328880 193511 328883
rect 203021 328883 203079 328889
rect 203021 328880 203033 328883
rect 193499 328852 203033 328880
rect 193499 328849 193511 328852
rect 193453 328843 193511 328849
rect 203021 328849 203033 328852
rect 203067 328849 203079 328883
rect 203021 328843 203079 328849
rect 285910 328228 285916 328280
rect 285968 328268 285974 328280
rect 325654 328268 325660 328280
rect 285968 328240 325660 328268
rect 285968 328228 285974 328240
rect 325654 328228 325660 328240
rect 325712 328228 325718 328280
rect 345250 327616 345256 327668
rect 345308 327656 345314 327668
rect 346078 327656 346084 327668
rect 345308 327628 346084 327656
rect 345308 327616 345314 327628
rect 346078 327616 346084 327628
rect 346136 327616 346142 327668
rect 76058 327548 76064 327600
rect 76116 327588 76122 327600
rect 100990 327588 100996 327600
rect 76116 327560 100996 327588
rect 76116 327548 76122 327560
rect 100990 327548 100996 327560
rect 101048 327588 101054 327600
rect 102278 327588 102284 327600
rect 101048 327560 102284 327588
rect 101048 327548 101054 327560
rect 102278 327548 102284 327560
rect 102336 327548 102342 327600
rect 137330 327548 137336 327600
rect 137388 327588 137394 327600
rect 137514 327588 137520 327600
rect 137388 327560 137520 327588
rect 137388 327548 137394 327560
rect 137514 327548 137520 327560
rect 137572 327548 137578 327600
rect 137698 327548 137704 327600
rect 137756 327588 137762 327600
rect 160974 327588 160980 327600
rect 137756 327560 160980 327588
rect 137756 327548 137762 327560
rect 160974 327548 160980 327560
rect 161032 327588 161038 327600
rect 209274 327588 209280 327600
rect 161032 327560 209280 327588
rect 161032 327548 161038 327560
rect 209274 327548 209280 327560
rect 209332 327548 209338 327600
rect 231446 327548 231452 327600
rect 231504 327588 231510 327600
rect 254354 327588 254360 327600
rect 231504 327560 254360 327588
rect 231504 327548 231510 327560
rect 254354 327548 254360 327560
rect 254412 327588 254418 327600
rect 303114 327588 303120 327600
rect 254412 327560 303120 327588
rect 254412 327548 254418 327560
rect 303114 327548 303120 327560
rect 303172 327548 303178 327600
rect 337154 327548 337160 327600
rect 337212 327588 337218 327600
rect 352794 327588 352800 327600
rect 337212 327560 352800 327588
rect 337212 327548 337218 327560
rect 352794 327548 352800 327560
rect 352852 327548 352858 327600
rect 137532 327520 137560 327548
rect 158398 327520 158404 327532
rect 137532 327492 158404 327520
rect 158398 327480 158404 327492
rect 158456 327480 158462 327532
rect 239542 327480 239548 327532
rect 239600 327520 239606 327532
rect 248834 327520 248840 327532
rect 239600 327492 248840 327520
rect 239600 327480 239606 327492
rect 248834 327480 248840 327492
rect 248892 327480 248898 327532
rect 249570 327480 249576 327532
rect 249628 327520 249634 327532
rect 250401 327523 250459 327529
rect 250401 327520 250413 327523
rect 249628 327492 250413 327520
rect 249628 327480 249634 327492
rect 250401 327489 250413 327492
rect 250447 327489 250459 327523
rect 250401 327483 250459 327489
rect 250490 327480 250496 327532
rect 250548 327520 250554 327532
rect 288670 327520 288676 327532
rect 250548 327492 288676 327520
rect 250548 327480 250554 327492
rect 288670 327480 288676 327492
rect 288728 327480 288734 327532
rect 341294 327480 341300 327532
rect 341352 327520 341358 327532
rect 357578 327520 357584 327532
rect 341352 327492 357584 327520
rect 341352 327480 341358 327492
rect 357578 327480 357584 327492
rect 357636 327480 357642 327532
rect 137790 327412 137796 327464
rect 137848 327452 137854 327464
rect 155914 327452 155920 327464
rect 137848 327424 155920 327452
rect 137848 327412 137854 327424
rect 155914 327412 155920 327424
rect 155972 327452 155978 327464
rect 192070 327452 192076 327464
rect 155972 327424 192076 327452
rect 155972 327412 155978 327424
rect 192070 327412 192076 327424
rect 192128 327412 192134 327464
rect 231998 327412 232004 327464
rect 232056 327452 232062 327464
rect 249110 327452 249116 327464
rect 232056 327424 249116 327452
rect 232056 327412 232062 327424
rect 249110 327412 249116 327424
rect 249168 327452 249174 327464
rect 281770 327452 281776 327464
rect 249168 327424 281776 327452
rect 249168 327412 249174 327424
rect 281770 327412 281776 327424
rect 281828 327412 281834 327464
rect 341018 327412 341024 327464
rect 341076 327452 341082 327464
rect 356014 327452 356020 327464
rect 341076 327424 356020 327452
rect 341076 327412 341082 327424
rect 356014 327412 356020 327424
rect 356072 327412 356078 327464
rect 58302 327344 58308 327396
rect 58360 327384 58366 327396
rect 59222 327384 59228 327396
rect 58360 327356 59228 327384
rect 58360 327344 58366 327356
rect 59222 327344 59228 327356
rect 59280 327344 59286 327396
rect 62350 327344 62356 327396
rect 62408 327384 62414 327396
rect 63362 327384 63368 327396
rect 62408 327356 63368 327384
rect 62408 327344 62414 327356
rect 63362 327344 63368 327356
rect 63420 327344 63426 327396
rect 65202 327344 65208 327396
rect 65260 327384 65266 327396
rect 68514 327384 68520 327396
rect 65260 327356 68520 327384
rect 65260 327344 65266 327356
rect 68514 327344 68520 327356
rect 68572 327344 68578 327396
rect 154810 327344 154816 327396
rect 154868 327384 154874 327396
rect 187930 327384 187936 327396
rect 154868 327356 187936 327384
rect 154868 327344 154874 327356
rect 187930 327344 187936 327356
rect 187988 327384 187994 327396
rect 189218 327384 189224 327396
rect 187988 327356 189224 327384
rect 187988 327344 187994 327356
rect 189218 327344 189224 327356
rect 189276 327344 189282 327396
rect 241750 327344 241756 327396
rect 241808 327384 241814 327396
rect 242762 327384 242768 327396
rect 241808 327356 242768 327384
rect 241808 327344 241814 327356
rect 242762 327344 242768 327356
rect 242820 327344 242826 327396
rect 248926 327344 248932 327396
rect 248984 327384 248990 327396
rect 256286 327384 256292 327396
rect 248984 327356 256292 327384
rect 248984 327344 248990 327356
rect 256286 327344 256292 327356
rect 256344 327344 256350 327396
rect 256381 327387 256439 327393
rect 256381 327353 256393 327387
rect 256427 327384 256439 327387
rect 265305 327387 265363 327393
rect 265305 327384 265317 327387
rect 256427 327356 265317 327384
rect 256427 327353 256439 327356
rect 256381 327347 256439 327353
rect 265305 327353 265317 327356
rect 265351 327353 265363 327387
rect 265305 327347 265363 327353
rect 339638 327344 339644 327396
rect 339696 327384 339702 327396
rect 353622 327384 353628 327396
rect 339696 327356 353628 327384
rect 339696 327344 339702 327356
rect 353622 327344 353628 327356
rect 353680 327344 353686 327396
rect 150854 327276 150860 327328
rect 150912 327316 150918 327328
rect 165206 327316 165212 327328
rect 150912 327288 165212 327316
rect 150912 327276 150918 327288
rect 165206 327276 165212 327288
rect 165264 327276 165270 327328
rect 342398 327276 342404 327328
rect 342456 327316 342462 327328
rect 355554 327316 355560 327328
rect 342456 327288 355560 327316
rect 342456 327276 342462 327288
rect 355554 327276 355560 327288
rect 355612 327276 355618 327328
rect 149382 327208 149388 327260
rect 149440 327248 149446 327260
rect 163274 327248 163280 327260
rect 149440 327220 163280 327248
rect 149440 327208 149446 327220
rect 163274 327208 163280 327220
rect 163332 327208 163338 327260
rect 243777 327251 243835 327257
rect 243777 327217 243789 327251
rect 243823 327248 243835 327251
rect 250490 327248 250496 327260
rect 243823 327220 250496 327248
rect 243823 327217 243835 327220
rect 243777 327211 243835 327217
rect 250490 327208 250496 327220
rect 250548 327208 250554 327260
rect 250585 327251 250643 327257
rect 250585 327217 250597 327251
rect 250631 327248 250643 327251
rect 256381 327251 256439 327257
rect 256381 327248 256393 327251
rect 250631 327220 256393 327248
rect 250631 327217 250643 327220
rect 250585 327211 250643 327217
rect 256381 327217 256393 327220
rect 256427 327217 256439 327251
rect 256381 327211 256439 327217
rect 256473 327251 256531 327257
rect 256473 327217 256485 327251
rect 256519 327248 256531 327251
rect 258402 327248 258408 327260
rect 256519 327220 258408 327248
rect 256519 327217 256531 327220
rect 256473 327211 256531 327217
rect 258402 327208 258408 327220
rect 258460 327208 258466 327260
rect 345618 327208 345624 327260
rect 345676 327248 345682 327260
rect 359694 327248 359700 327260
rect 345676 327220 359700 327248
rect 345676 327208 345682 327220
rect 359694 327208 359700 327220
rect 359752 327208 359758 327260
rect 152234 327140 152240 327192
rect 152292 327180 152298 327192
rect 166126 327180 166132 327192
rect 152292 327152 166132 327180
rect 152292 327140 152298 327152
rect 166126 327140 166132 327152
rect 166184 327140 166190 327192
rect 238622 327140 238628 327192
rect 238680 327180 238686 327192
rect 244418 327180 244424 327192
rect 238680 327152 244424 327180
rect 238680 327140 238686 327152
rect 244418 327140 244424 327152
rect 244476 327140 244482 327192
rect 247178 327140 247184 327192
rect 247236 327180 247242 327192
rect 258954 327180 258960 327192
rect 247236 327152 258960 327180
rect 247236 327140 247242 327152
rect 258954 327140 258960 327152
rect 259012 327140 259018 327192
rect 344790 327140 344796 327192
rect 344848 327180 344854 327192
rect 358314 327180 358320 327192
rect 344848 327152 358320 327180
rect 344848 327140 344854 327152
rect 358314 327140 358320 327152
rect 358372 327140 358378 327192
rect 154074 327072 154080 327124
rect 154132 327112 154138 327124
rect 168058 327112 168064 327124
rect 154132 327084 168064 327112
rect 154132 327072 154138 327084
rect 168058 327072 168064 327084
rect 168116 327072 168122 327124
rect 194830 327072 194836 327124
rect 194888 327112 194894 327124
rect 232090 327112 232096 327124
rect 194888 327084 232096 327112
rect 194888 327072 194894 327084
rect 232090 327072 232096 327084
rect 232148 327112 232154 327124
rect 243777 327115 243835 327121
rect 243777 327112 243789 327115
rect 232148 327084 243789 327112
rect 232148 327072 232154 327084
rect 243777 327081 243789 327084
rect 243823 327081 243835 327115
rect 243777 327075 243835 327081
rect 244234 327072 244240 327124
rect 244292 327112 244298 327124
rect 257298 327112 257304 327124
rect 244292 327084 257304 327112
rect 244292 327072 244298 327084
rect 257298 327072 257304 327084
rect 257356 327072 257362 327124
rect 288670 327072 288676 327124
rect 288728 327112 288734 327124
rect 325102 327112 325108 327124
rect 288728 327084 325108 327112
rect 288728 327072 288734 327084
rect 325102 327072 325108 327084
rect 325160 327072 325166 327124
rect 341202 327072 341208 327124
rect 341260 327112 341266 327124
rect 358406 327112 358412 327124
rect 341260 327084 358412 327112
rect 341260 327072 341266 327084
rect 358406 327072 358412 327084
rect 358464 327072 358470 327124
rect 150762 327004 150768 327056
rect 150820 327044 150826 327056
rect 164562 327044 164568 327056
rect 150820 327016 164568 327044
rect 150820 327004 150826 327016
rect 164562 327004 164568 327016
rect 164620 327004 164626 327056
rect 192070 327004 192076 327056
rect 192128 327044 192134 327056
rect 233470 327044 233476 327056
rect 192128 327016 233476 327044
rect 192128 327004 192134 327016
rect 233470 327004 233476 327016
rect 233528 327044 233534 327056
rect 249570 327044 249576 327056
rect 233528 327016 249576 327044
rect 233528 327004 233534 327016
rect 249570 327004 249576 327016
rect 249628 327004 249634 327056
rect 250030 327004 250036 327056
rect 250088 327044 250094 327056
rect 264106 327044 264112 327056
rect 250088 327016 264112 327044
rect 250088 327004 250094 327016
rect 264106 327004 264112 327016
rect 264164 327004 264170 327056
rect 281770 327004 281776 327056
rect 281828 327044 281834 327056
rect 282874 327044 282880 327056
rect 281828 327016 282880 327044
rect 281828 327004 281834 327016
rect 282874 327004 282880 327016
rect 282932 327044 282938 327056
rect 325562 327044 325568 327056
rect 282932 327016 325568 327044
rect 282932 327004 282938 327016
rect 325562 327004 325568 327016
rect 325620 327004 325626 327056
rect 339914 327004 339920 327056
rect 339972 327044 339978 327056
rect 356750 327044 356756 327056
rect 339972 327016 356756 327044
rect 339972 327004 339978 327016
rect 356750 327004 356756 327016
rect 356808 327004 356814 327056
rect 137606 326936 137612 326988
rect 137664 326976 137670 326988
rect 154810 326976 154816 326988
rect 137664 326948 154816 326976
rect 137664 326936 137670 326948
rect 154810 326936 154816 326948
rect 154868 326936 154874 326988
rect 156282 326936 156288 326988
rect 156340 326976 156346 326988
rect 169990 326976 169996 326988
rect 156340 326948 169996 326976
rect 156340 326936 156346 326948
rect 169990 326936 169996 326948
rect 170048 326936 170054 326988
rect 189218 326936 189224 326988
rect 189276 326976 189282 326988
rect 230710 326976 230716 326988
rect 189276 326948 230716 326976
rect 189276 326936 189282 326948
rect 230710 326936 230716 326948
rect 230768 326976 230774 326988
rect 231998 326976 232004 326988
rect 230768 326948 232004 326976
rect 230768 326936 230774 326948
rect 231998 326936 232004 326948
rect 232056 326936 232062 326988
rect 248282 326936 248288 326988
rect 248340 326976 248346 326988
rect 365214 326976 365220 326988
rect 248340 326948 365220 326976
rect 248340 326936 248346 326948
rect 365214 326936 365220 326948
rect 365272 326936 365278 326988
rect 102278 326868 102284 326920
rect 102336 326908 102342 326920
rect 136962 326908 136968 326920
rect 102336 326880 136968 326908
rect 102336 326868 102342 326880
rect 136962 326868 136968 326880
rect 137020 326868 137026 326920
rect 154258 326868 154264 326920
rect 154316 326908 154322 326920
rect 326574 326908 326580 326920
rect 154316 326880 326580 326908
rect 154316 326868 154322 326880
rect 326574 326868 326580 326880
rect 326632 326868 326638 326920
rect 335682 326868 335688 326920
rect 335740 326908 335746 326920
rect 336786 326908 336792 326920
rect 335740 326880 336792 326908
rect 335740 326868 335746 326880
rect 336786 326868 336792 326880
rect 336844 326868 336850 326920
rect 338534 326868 338540 326920
rect 338592 326908 338598 326920
rect 355186 326908 355192 326920
rect 338592 326880 355192 326908
rect 338592 326868 338598 326880
rect 355186 326868 355192 326880
rect 355244 326868 355250 326920
rect 154902 326800 154908 326852
rect 154960 326840 154966 326852
rect 169070 326840 169076 326852
rect 154960 326812 169076 326840
rect 154960 326800 154966 326812
rect 169070 326800 169076 326812
rect 169128 326800 169134 326852
rect 238990 326800 238996 326852
rect 239048 326840 239054 326852
rect 239910 326840 239916 326852
rect 239048 326812 239916 326840
rect 239048 326800 239054 326812
rect 239910 326800 239916 326812
rect 239968 326800 239974 326852
rect 245890 326800 245896 326852
rect 245948 326840 245954 326852
rect 260150 326840 260156 326852
rect 245948 326812 260156 326840
rect 245948 326800 245954 326812
rect 260150 326800 260156 326812
rect 260208 326800 260214 326852
rect 334210 326800 334216 326852
rect 334268 326840 334274 326852
rect 335222 326840 335228 326852
rect 334268 326812 335228 326840
rect 334268 326800 334274 326812
rect 335222 326800 335228 326812
rect 335280 326800 335286 326852
rect 339362 326800 339368 326852
rect 339420 326840 339426 326852
rect 354358 326840 354364 326852
rect 339420 326812 354364 326840
rect 339420 326800 339426 326812
rect 354358 326800 354364 326812
rect 354416 326800 354422 326852
rect 153522 326732 153528 326784
rect 153580 326772 153586 326784
rect 167322 326772 167328 326784
rect 153580 326744 167328 326772
rect 153580 326732 153586 326744
rect 167322 326732 167328 326744
rect 167380 326732 167386 326784
rect 247270 326732 247276 326784
rect 247328 326772 247334 326784
rect 261162 326772 261168 326784
rect 247328 326744 261168 326772
rect 247328 326732 247334 326744
rect 261162 326732 261168 326744
rect 261220 326732 261226 326784
rect 343226 326732 343232 326784
rect 343284 326772 343290 326784
rect 355646 326772 355652 326784
rect 343284 326744 355652 326772
rect 343284 326732 343290 326744
rect 355646 326732 355652 326744
rect 355704 326732 355710 326784
rect 144598 326664 144604 326716
rect 144656 326704 144662 326716
rect 156190 326704 156196 326716
rect 144656 326676 156196 326704
rect 144656 326664 144662 326676
rect 156190 326664 156196 326676
rect 156248 326664 156254 326716
rect 157573 326707 157631 326713
rect 157573 326673 157585 326707
rect 157619 326704 157631 326707
rect 164473 326707 164531 326713
rect 164473 326704 164485 326707
rect 157619 326676 164485 326704
rect 157619 326673 157631 326676
rect 157573 326667 157631 326673
rect 164473 326673 164485 326676
rect 164519 326673 164531 326707
rect 164473 326667 164531 326673
rect 248650 326664 248656 326716
rect 248708 326704 248714 326716
rect 263094 326704 263100 326716
rect 248708 326676 263100 326704
rect 248708 326664 248714 326676
rect 263094 326664 263100 326676
rect 263152 326664 263158 326716
rect 340834 326664 340840 326716
rect 340892 326704 340898 326716
rect 352794 326704 352800 326716
rect 340892 326676 352800 326704
rect 340892 326664 340898 326676
rect 352794 326664 352800 326676
rect 352852 326664 352858 326716
rect 65110 326596 65116 326648
rect 65168 326636 65174 326648
rect 69618 326636 69624 326648
rect 65168 326608 69624 326636
rect 65168 326596 65174 326608
rect 69618 326596 69624 326608
rect 69676 326596 69682 326648
rect 147450 326596 147456 326648
rect 147508 326636 147514 326648
rect 159042 326636 159048 326648
rect 147508 326608 159048 326636
rect 147508 326596 147514 326608
rect 159042 326596 159048 326608
rect 159100 326596 159106 326648
rect 241474 326596 241480 326648
rect 241532 326636 241538 326648
rect 252882 326636 252888 326648
rect 241532 326608 252888 326636
rect 241532 326596 241538 326608
rect 252882 326596 252888 326608
rect 252940 326596 252946 326648
rect 259690 326596 259696 326648
rect 259748 326636 259754 326648
rect 262082 326636 262088 326648
rect 259748 326608 262088 326636
rect 259748 326596 259754 326608
rect 262082 326596 262088 326608
rect 262140 326596 262146 326648
rect 341570 326596 341576 326648
rect 341628 326636 341634 326648
rect 354174 326636 354180 326648
rect 341628 326608 354180 326636
rect 341628 326596 341634 326608
rect 354174 326596 354180 326608
rect 354232 326596 354238 326648
rect 148462 326528 148468 326580
rect 148520 326568 148526 326580
rect 160238 326568 160244 326580
rect 148520 326540 160244 326568
rect 148520 326528 148526 326540
rect 160238 326528 160244 326540
rect 160296 326528 160302 326580
rect 246350 326528 246356 326580
rect 246408 326568 246414 326580
rect 258310 326568 258316 326580
rect 246408 326540 258316 326568
rect 246408 326528 246414 326540
rect 258310 326528 258316 326540
rect 258368 326528 258374 326580
rect 332922 326528 332928 326580
rect 332980 326568 332986 326580
rect 333658 326568 333664 326580
rect 332980 326540 333664 326568
rect 332980 326528 332986 326540
rect 333658 326528 333664 326540
rect 333716 326528 333722 326580
rect 343962 326528 343968 326580
rect 344020 326568 344026 326580
rect 356934 326568 356940 326580
rect 344020 326540 356940 326568
rect 344020 326528 344026 326540
rect 356934 326528 356940 326540
rect 356992 326528 356998 326580
rect 136962 326460 136968 326512
rect 137020 326500 137026 326512
rect 137020 326472 138296 326500
rect 137020 326460 137026 326472
rect 138268 326432 138296 326472
rect 150394 326460 150400 326512
rect 150452 326500 150458 326512
rect 158950 326500 158956 326512
rect 150452 326472 158956 326500
rect 150452 326460 150458 326472
rect 158950 326460 158956 326472
rect 159008 326460 159014 326512
rect 242486 326460 242492 326512
rect 242544 326500 242550 326512
rect 254078 326500 254084 326512
rect 242544 326472 254084 326500
rect 242544 326460 242550 326472
rect 254078 326460 254084 326472
rect 254136 326460 254142 326512
rect 337062 326460 337068 326512
rect 337120 326500 337126 326512
rect 351966 326500 351972 326512
rect 337120 326472 351972 326500
rect 337120 326460 337126 326472
rect 351966 326460 351972 326472
rect 352024 326460 352030 326512
rect 152053 326435 152111 326441
rect 152053 326432 152065 326435
rect 138268 326404 152065 326432
rect 152053 326401 152065 326404
rect 152099 326401 152111 326435
rect 152053 326395 152111 326401
rect 152142 326392 152148 326444
rect 152200 326432 152206 326444
rect 162998 326432 163004 326444
rect 152200 326404 163004 326432
rect 152200 326392 152206 326404
rect 162998 326392 163004 326404
rect 163056 326392 163062 326444
rect 244326 326392 244332 326444
rect 244384 326432 244390 326444
rect 253526 326432 253532 326444
rect 244384 326404 253532 326432
rect 244384 326392 244390 326404
rect 253526 326392 253532 326404
rect 253584 326392 253590 326444
rect 74034 326324 74040 326376
rect 74092 326364 74098 326376
rect 76058 326364 76064 326376
rect 74092 326336 76064 326364
rect 74092 326324 74098 326336
rect 76058 326324 76064 326336
rect 76116 326324 76122 326376
rect 145518 326324 145524 326376
rect 145576 326364 145582 326376
rect 152326 326364 152332 326376
rect 145576 326336 152332 326364
rect 145576 326324 145582 326336
rect 152326 326324 152332 326336
rect 152384 326324 152390 326376
rect 152421 326367 152479 326373
rect 152421 326333 152433 326367
rect 152467 326364 152479 326367
rect 156834 326364 156840 326376
rect 152467 326336 156840 326364
rect 152467 326333 152479 326336
rect 152421 326327 152479 326333
rect 156834 326324 156840 326336
rect 156892 326364 156898 326376
rect 157573 326367 157631 326373
rect 157573 326364 157585 326367
rect 156892 326336 157585 326364
rect 156892 326324 156898 326336
rect 157573 326333 157585 326336
rect 157619 326333 157631 326367
rect 157573 326327 157631 326333
rect 244510 326324 244516 326376
rect 244568 326364 244574 326376
rect 256473 326367 256531 326373
rect 256473 326364 256485 326367
rect 244568 326336 256485 326364
rect 244568 326324 244574 326336
rect 256473 326333 256485 326336
rect 256519 326333 256531 326367
rect 256473 326327 256531 326333
rect 75782 326256 75788 326308
rect 75840 326296 75846 326308
rect 76978 326296 76984 326308
rect 75840 326268 76984 326296
rect 75840 326256 75846 326268
rect 76978 326256 76984 326268
rect 77036 326256 77042 326308
rect 145334 326256 145340 326308
rect 145392 326296 145398 326308
rect 145886 326296 145892 326308
rect 145392 326268 145892 326296
rect 145392 326256 145398 326268
rect 145886 326256 145892 326268
rect 145944 326256 145950 326308
rect 147910 326256 147916 326308
rect 147968 326296 147974 326308
rect 148738 326296 148744 326308
rect 147968 326268 148744 326296
rect 147968 326256 147974 326268
rect 148738 326256 148744 326268
rect 148796 326256 148802 326308
rect 151314 326256 151320 326308
rect 151372 326296 151378 326308
rect 154810 326296 154816 326308
rect 151372 326268 154816 326296
rect 151372 326256 151378 326268
rect 154810 326256 154816 326268
rect 154868 326256 154874 326308
rect 155638 326256 155644 326308
rect 155696 326296 155702 326308
rect 162262 326296 162268 326308
rect 155696 326268 162268 326296
rect 155696 326256 155702 326268
rect 162262 326256 162268 326268
rect 162320 326256 162326 326308
rect 164473 326299 164531 326305
rect 164473 326265 164485 326299
rect 164519 326296 164531 326299
rect 194830 326296 194836 326308
rect 164519 326268 194836 326296
rect 164519 326265 164531 326268
rect 164473 326259 164531 326265
rect 194830 326256 194836 326268
rect 194888 326256 194894 326308
rect 243222 326256 243228 326308
rect 243280 326296 243286 326308
rect 244234 326296 244240 326308
rect 243280 326268 244240 326296
rect 243280 326256 243286 326268
rect 244234 326256 244240 326268
rect 244292 326256 244298 326308
rect 245338 326256 245344 326308
rect 245396 326296 245402 326308
rect 248742 326296 248748 326308
rect 245396 326268 248748 326296
rect 245396 326256 245402 326268
rect 248742 326256 248748 326268
rect 248800 326256 248806 326308
rect 254538 326256 254544 326308
rect 254596 326296 254602 326308
rect 259230 326296 259236 326308
rect 254596 326268 259236 326296
rect 254596 326256 254602 326268
rect 259230 326256 259236 326268
rect 259288 326256 259294 326308
rect 70630 325236 70636 325288
rect 70688 325276 70694 325288
rect 71366 325276 71372 325288
rect 70688 325248 71372 325276
rect 70688 325236 70694 325248
rect 71366 325236 71372 325248
rect 71424 325236 71430 325288
rect 348010 325168 348016 325220
rect 348068 325208 348074 325220
rect 348470 325208 348476 325220
rect 348068 325180 348476 325208
rect 348068 325168 348074 325180
rect 348470 325168 348476 325180
rect 348528 325168 348534 325220
rect 54070 324828 54076 324880
rect 54128 324868 54134 324880
rect 54806 324868 54812 324880
rect 54128 324840 54812 324868
rect 54128 324828 54134 324840
rect 54806 324828 54812 324840
rect 54864 324828 54870 324880
rect 325102 324828 325108 324880
rect 325160 324868 325166 324880
rect 343962 324868 343968 324880
rect 325160 324840 343968 324868
rect 325160 324828 325166 324840
rect 343962 324828 343968 324840
rect 344020 324868 344026 324880
rect 347182 324868 347188 324880
rect 344020 324840 347188 324868
rect 344020 324828 344026 324840
rect 347182 324828 347188 324840
rect 347240 324828 347246 324880
rect 279102 324760 279108 324812
rect 279160 324800 279166 324812
rect 280298 324800 280304 324812
rect 279160 324772 280304 324800
rect 279160 324760 279166 324772
rect 280298 324760 280304 324772
rect 280356 324760 280362 324812
rect 291522 324760 291528 324812
rect 291580 324800 291586 324812
rect 292718 324800 292724 324812
rect 291580 324772 292724 324800
rect 291580 324760 291586 324772
rect 292718 324760 292724 324772
rect 292776 324760 292782 324812
rect 210010 324148 210016 324200
rect 210068 324188 210074 324200
rect 211298 324188 211304 324200
rect 210068 324160 211304 324188
rect 210068 324148 210074 324160
rect 211298 324148 211304 324160
rect 211356 324148 211362 324200
rect 344790 324080 344796 324132
rect 344848 324120 344854 324132
rect 348102 324120 348108 324132
rect 344848 324092 348108 324120
rect 344848 324080 344854 324092
rect 348102 324080 348108 324092
rect 348160 324080 348166 324132
rect 304034 324012 304040 324064
rect 304092 324052 304098 324064
rect 305138 324052 305144 324064
rect 304092 324024 305144 324052
rect 304092 324012 304098 324024
rect 305138 324012 305144 324024
rect 305196 324012 305202 324064
rect 325746 323468 325752 323520
rect 325804 323508 325810 323520
rect 344790 323508 344796 323520
rect 325804 323480 344796 323508
rect 325804 323468 325810 323480
rect 344790 323468 344796 323480
rect 344848 323468 344854 323520
rect 343870 322788 343876 322840
rect 343928 322828 343934 322840
rect 345158 322828 345164 322840
rect 343928 322800 345164 322828
rect 343928 322788 343934 322800
rect 345158 322788 345164 322800
rect 345216 322828 345222 322840
rect 348010 322828 348016 322840
rect 345216 322800 348016 322828
rect 345216 322788 345222 322800
rect 348010 322788 348016 322800
rect 348068 322788 348074 322840
rect 324550 322720 324556 322772
rect 324608 322760 324614 322772
rect 325378 322760 325384 322772
rect 324608 322732 325384 322760
rect 324608 322720 324614 322732
rect 325378 322720 325384 322732
rect 325436 322720 325442 322772
rect 325194 322176 325200 322228
rect 325252 322216 325258 322228
rect 343870 322216 343876 322228
rect 325252 322188 343876 322216
rect 325252 322176 325258 322188
rect 343870 322176 343876 322188
rect 343928 322176 343934 322228
rect 13958 322108 13964 322160
rect 14016 322148 14022 322160
rect 16350 322148 16356 322160
rect 14016 322120 16356 322148
rect 14016 322108 14022 322120
rect 16350 322108 16356 322120
rect 16408 322108 16414 322160
rect 325378 322108 325384 322160
rect 325436 322148 325442 322160
rect 346998 322148 347004 322160
rect 325436 322120 347004 322148
rect 325436 322108 325442 322120
rect 346998 322108 347004 322120
rect 347056 322148 347062 322160
rect 351230 322148 351236 322160
rect 347056 322120 351236 322148
rect 347056 322108 347062 322120
rect 351230 322108 351236 322120
rect 351288 322108 351294 322160
rect 342490 322040 342496 322092
rect 342548 322080 342554 322092
rect 345250 322080 345256 322092
rect 342548 322052 345256 322080
rect 342548 322040 342554 322052
rect 345250 322040 345256 322052
rect 345308 322040 345314 322092
rect 325654 320748 325660 320800
rect 325712 320788 325718 320800
rect 342490 320788 342496 320800
rect 325712 320760 342496 320788
rect 325712 320748 325718 320760
rect 342490 320748 342496 320760
rect 342548 320788 342554 320800
rect 342950 320788 342956 320800
rect 342548 320760 342956 320788
rect 342548 320748 342554 320760
rect 342950 320748 342956 320760
rect 343008 320748 343014 320800
rect 324734 320680 324740 320732
rect 324792 320720 324798 320732
rect 346446 320720 346452 320732
rect 324792 320692 346452 320720
rect 324792 320680 324798 320692
rect 346446 320680 346452 320692
rect 346504 320720 346510 320732
rect 349482 320720 349488 320732
rect 346504 320692 349488 320720
rect 346504 320680 346510 320692
rect 349482 320680 349488 320692
rect 349540 320680 349546 320732
rect 62442 320612 62448 320664
rect 62500 320652 62506 320664
rect 67686 320652 67692 320664
rect 62500 320624 67692 320652
rect 62500 320612 62506 320624
rect 67686 320612 67692 320624
rect 67744 320612 67750 320664
rect 150854 320612 150860 320664
rect 150912 320652 150918 320664
rect 151958 320652 151964 320664
rect 150912 320624 151964 320652
rect 150912 320612 150918 320624
rect 151958 320612 151964 320624
rect 152016 320612 152022 320664
rect 156190 320612 156196 320664
rect 156248 320652 156254 320664
rect 156926 320652 156932 320664
rect 156248 320624 156932 320652
rect 156248 320612 156254 320624
rect 156926 320612 156932 320624
rect 156984 320612 156990 320664
rect 158950 320612 158956 320664
rect 159008 320652 159014 320664
rect 162630 320652 162636 320664
rect 159008 320624 162636 320652
rect 159008 320612 159014 320624
rect 162630 320612 162636 320624
rect 162688 320612 162694 320664
rect 243222 320612 243228 320664
rect 243280 320652 243286 320664
rect 243774 320652 243780 320664
rect 243280 320624 243780 320652
rect 243280 320612 243286 320624
rect 243774 320612 243780 320624
rect 243832 320612 243838 320664
rect 245890 320612 245896 320664
rect 245948 320652 245954 320664
rect 246442 320652 246448 320664
rect 245948 320624 246448 320652
rect 245948 320612 245954 320624
rect 246442 320612 246448 320624
rect 246500 320612 246506 320664
rect 250950 320652 250956 320664
rect 246552 320624 250956 320652
rect 63730 320544 63736 320596
rect 63788 320584 63794 320596
rect 69434 320584 69440 320596
rect 63788 320556 69440 320584
rect 63788 320544 63794 320556
rect 69434 320544 69440 320556
rect 69492 320544 69498 320596
rect 154810 320544 154816 320596
rect 154868 320584 154874 320596
rect 163458 320584 163464 320596
rect 154868 320556 163464 320584
rect 154868 320544 154874 320556
rect 163458 320544 163464 320556
rect 163516 320544 163522 320596
rect 244418 320544 244424 320596
rect 244476 320584 244482 320596
rect 246552 320584 246580 320624
rect 250950 320612 250956 320624
rect 251008 320612 251014 320664
rect 337154 320612 337160 320664
rect 337212 320652 337218 320664
rect 337522 320652 337528 320664
rect 337212 320624 337528 320652
rect 337212 320612 337218 320624
rect 337522 320612 337528 320624
rect 337580 320612 337586 320664
rect 339914 320612 339920 320664
rect 339972 320652 339978 320664
rect 340558 320652 340564 320664
rect 339972 320624 340564 320652
rect 339972 320612 339978 320624
rect 340558 320612 340564 320624
rect 340616 320612 340622 320664
rect 248926 320584 248932 320596
rect 244476 320556 246580 320584
rect 246644 320556 248932 320584
rect 244476 320544 244482 320556
rect 58210 320476 58216 320528
rect 58268 320516 58274 320528
rect 64098 320516 64104 320528
rect 58268 320488 64104 320516
rect 58268 320476 58274 320488
rect 64098 320476 64104 320488
rect 64156 320476 64162 320528
rect 65110 320516 65116 320528
rect 64208 320488 65116 320516
rect 57934 320408 57940 320460
rect 57992 320448 57998 320460
rect 64208 320448 64236 320488
rect 65110 320476 65116 320488
rect 65168 320476 65174 320528
rect 243590 320476 243596 320528
rect 243648 320516 243654 320528
rect 246644 320516 246672 320556
rect 248926 320544 248932 320556
rect 248984 320544 248990 320596
rect 332922 320544 332928 320596
rect 332980 320584 332986 320596
rect 348562 320584 348568 320596
rect 332980 320556 348568 320584
rect 332980 320544 332986 320556
rect 348562 320544 348568 320556
rect 348620 320544 348626 320596
rect 352794 320544 352800 320596
rect 352852 320544 352858 320596
rect 243648 320488 246672 320516
rect 243648 320476 243654 320488
rect 248650 320476 248656 320528
rect 248708 320516 248714 320528
rect 249110 320516 249116 320528
rect 248708 320488 249116 320516
rect 248708 320476 248714 320488
rect 249110 320476 249116 320488
rect 249168 320476 249174 320528
rect 331450 320476 331456 320528
rect 331508 320516 331514 320528
rect 340377 320519 340435 320525
rect 340377 320516 340389 320519
rect 331508 320488 340389 320516
rect 331508 320476 331514 320488
rect 340377 320485 340389 320488
rect 340423 320485 340435 320519
rect 340377 320479 340435 320485
rect 340466 320476 340472 320528
rect 340524 320516 340530 320528
rect 341018 320516 341024 320528
rect 340524 320488 341024 320516
rect 340524 320476 340530 320488
rect 341018 320476 341024 320488
rect 341076 320476 341082 320528
rect 352242 320516 352248 320528
rect 341128 320488 352248 320516
rect 57992 320420 64236 320448
rect 64285 320451 64343 320457
rect 57992 320408 57998 320420
rect 64285 320417 64297 320451
rect 64331 320448 64343 320451
rect 65202 320448 65208 320460
rect 64331 320420 65208 320448
rect 64331 320417 64343 320420
rect 64285 320411 64343 320417
rect 65202 320408 65208 320420
rect 65260 320408 65266 320460
rect 338442 320408 338448 320460
rect 338500 320448 338506 320460
rect 341128 320448 341156 320488
rect 352242 320476 352248 320488
rect 352300 320476 352306 320528
rect 352812 320516 352840 320544
rect 352886 320516 352892 320528
rect 352812 320488 352892 320516
rect 352886 320476 352892 320488
rect 352944 320476 352950 320528
rect 351598 320448 351604 320460
rect 338500 320420 341156 320448
rect 341220 320420 351604 320448
rect 338500 320408 338506 320420
rect 59682 320340 59688 320392
rect 59740 320380 59746 320392
rect 70630 320380 70636 320392
rect 59740 320352 70636 320380
rect 59740 320340 59746 320352
rect 70630 320340 70636 320352
rect 70688 320340 70694 320392
rect 336970 320340 336976 320392
rect 337028 320380 337034 320392
rect 341220 320380 341248 320420
rect 351598 320408 351604 320420
rect 351656 320408 351662 320460
rect 350402 320380 350408 320392
rect 337028 320352 341248 320380
rect 341312 320352 350408 320380
rect 337028 320340 337034 320352
rect 56094 320272 56100 320324
rect 56152 320312 56158 320324
rect 66582 320312 66588 320324
rect 56152 320284 66588 320312
rect 56152 320272 56158 320284
rect 66582 320272 66588 320284
rect 66640 320272 66646 320324
rect 248742 320272 248748 320324
rect 248800 320312 248806 320324
rect 257114 320312 257120 320324
rect 248800 320284 257120 320312
rect 248800 320272 248806 320284
rect 257114 320272 257120 320284
rect 257172 320272 257178 320324
rect 335590 320272 335596 320324
rect 335648 320312 335654 320324
rect 341312 320312 341340 320352
rect 350402 320340 350408 320352
rect 350460 320340 350466 320392
rect 335648 320284 341340 320312
rect 341389 320315 341447 320321
rect 335648 320272 335654 320284
rect 341389 320281 341401 320315
rect 341435 320312 341447 320315
rect 350954 320312 350960 320324
rect 341435 320284 350960 320312
rect 341435 320281 341447 320284
rect 341389 320275 341447 320281
rect 350954 320272 350960 320284
rect 351012 320272 351018 320324
rect 60602 320204 60608 320256
rect 60660 320244 60666 320256
rect 71918 320244 71924 320256
rect 60660 320216 71924 320244
rect 60660 320204 60666 320216
rect 71918 320204 71924 320216
rect 71976 320204 71982 320256
rect 332830 320204 332836 320256
rect 332888 320244 332894 320256
rect 348010 320244 348016 320256
rect 332888 320216 348016 320244
rect 332888 320204 332894 320216
rect 348010 320204 348016 320216
rect 348068 320204 348074 320256
rect 55266 320136 55272 320188
rect 55324 320176 55330 320188
rect 60237 320179 60295 320185
rect 60237 320176 60249 320179
rect 55324 320148 60249 320176
rect 55324 320136 55330 320148
rect 60237 320145 60249 320148
rect 60283 320145 60295 320179
rect 60237 320139 60295 320145
rect 62350 320136 62356 320188
rect 62408 320176 62414 320188
rect 74770 320176 74776 320188
rect 62408 320148 74776 320176
rect 62408 320136 62414 320148
rect 74770 320136 74776 320148
rect 74828 320136 74834 320188
rect 246258 320136 246264 320188
rect 246316 320176 246322 320188
rect 254538 320176 254544 320188
rect 246316 320148 254544 320176
rect 246316 320136 246322 320148
rect 254538 320136 254544 320148
rect 254596 320136 254602 320188
rect 325562 320136 325568 320188
rect 325620 320176 325626 320188
rect 325838 320176 325844 320188
rect 325620 320148 325844 320176
rect 325620 320136 325626 320148
rect 325838 320136 325844 320148
rect 325896 320136 325902 320188
rect 340377 320179 340435 320185
rect 340377 320145 340389 320179
rect 340423 320176 340435 320179
rect 347274 320176 347280 320188
rect 340423 320148 347280 320176
rect 340423 320145 340435 320148
rect 340377 320139 340435 320145
rect 347274 320136 347280 320148
rect 347332 320136 347338 320188
rect 59590 320068 59596 320120
rect 59648 320108 59654 320120
rect 65938 320108 65944 320120
rect 59648 320080 65944 320108
rect 59648 320068 59654 320080
rect 65938 320068 65944 320080
rect 65996 320068 66002 320120
rect 149290 320068 149296 320120
rect 149348 320108 149354 320120
rect 155638 320108 155644 320120
rect 149348 320080 155644 320108
rect 149348 320068 149354 320080
rect 155638 320068 155644 320080
rect 155696 320068 155702 320120
rect 248926 320068 248932 320120
rect 248984 320108 248990 320120
rect 259690 320108 259696 320120
rect 248984 320080 259696 320108
rect 248984 320068 248990 320080
rect 259690 320068 259696 320080
rect 259748 320068 259754 320120
rect 334302 320068 334308 320120
rect 334360 320108 334366 320120
rect 349390 320108 349396 320120
rect 334360 320080 349396 320108
rect 334360 320068 334366 320080
rect 349390 320068 349396 320080
rect 349448 320068 349454 320120
rect 61430 320000 61436 320052
rect 61488 320040 61494 320052
rect 73390 320040 73396 320052
rect 61488 320012 73396 320040
rect 61488 320000 61494 320012
rect 73390 320000 73396 320012
rect 73448 320000 73454 320052
rect 147910 320000 147916 320052
rect 147968 320040 147974 320052
rect 161710 320040 161716 320052
rect 147968 320012 161716 320040
rect 147968 320000 147974 320012
rect 161710 320000 161716 320012
rect 161768 320000 161774 320052
rect 241750 320000 241756 320052
rect 241808 320040 241814 320052
rect 255550 320040 255556 320052
rect 241808 320012 255556 320040
rect 241808 320000 241814 320012
rect 255550 320000 255556 320012
rect 255608 320000 255614 320052
rect 325102 320000 325108 320052
rect 325160 320040 325166 320052
rect 325562 320040 325568 320052
rect 325160 320012 325568 320040
rect 325160 320000 325166 320012
rect 325562 320000 325568 320012
rect 325620 320000 325626 320052
rect 334210 320000 334216 320052
rect 334268 320040 334274 320052
rect 349758 320040 349764 320052
rect 334268 320012 349764 320040
rect 334268 320000 334274 320012
rect 349758 320000 349764 320012
rect 349816 320000 349822 320052
rect 58762 319932 58768 319984
rect 58820 319972 58826 319984
rect 70722 319972 70728 319984
rect 58820 319944 70728 319972
rect 58820 319932 58826 319944
rect 70722 319932 70728 319944
rect 70780 319932 70786 319984
rect 145334 319932 145340 319984
rect 145392 319972 145398 319984
rect 159042 319972 159048 319984
rect 145392 319944 159048 319972
rect 145392 319932 145398 319944
rect 159042 319932 159048 319944
rect 159100 319932 159106 319984
rect 162998 319932 163004 319984
rect 163056 319972 163062 319984
rect 164378 319972 164384 319984
rect 163056 319944 164384 319972
rect 163056 319932 163062 319944
rect 164378 319932 164384 319944
rect 164436 319932 164442 319984
rect 238990 319932 238996 319984
rect 239048 319972 239054 319984
rect 252790 319972 252796 319984
rect 239048 319944 252796 319972
rect 239048 319932 239054 319944
rect 252790 319932 252796 319944
rect 252848 319932 252854 319984
rect 335682 319932 335688 319984
rect 335740 319972 335746 319984
rect 341389 319975 341447 319981
rect 341389 319972 341401 319975
rect 335740 319944 341401 319972
rect 335740 319932 335746 319944
rect 341389 319941 341401 319944
rect 341435 319941 341447 319975
rect 341389 319935 341447 319941
rect 349482 319932 349488 319984
rect 349540 319972 349546 319984
rect 429430 319972 429436 319984
rect 349540 319944 429436 319972
rect 349540 319932 349546 319944
rect 429430 319932 429436 319944
rect 429488 319932 429494 319984
rect 65021 319907 65079 319913
rect 65021 319873 65033 319907
rect 65067 319904 65079 319907
rect 66490 319904 66496 319916
rect 65067 319876 66496 319904
rect 65067 319873 65079 319876
rect 65021 319867 65079 319873
rect 66490 319864 66496 319876
rect 66548 319864 66554 319916
rect 60970 319796 60976 319848
rect 61028 319836 61034 319848
rect 66766 319836 66772 319848
rect 61028 319808 66772 319836
rect 61028 319796 61034 319808
rect 66766 319796 66772 319808
rect 66824 319796 66830 319848
rect 62442 319728 62448 319780
rect 62500 319768 62506 319780
rect 68606 319768 68612 319780
rect 62500 319740 68612 319768
rect 62500 319728 62506 319740
rect 68606 319728 68612 319740
rect 68664 319728 68670 319780
rect 338534 319728 338540 319780
rect 338592 319768 338598 319780
rect 339454 319768 339460 319780
rect 338592 319740 339460 319768
rect 338592 319728 338598 319740
rect 339454 319728 339460 319740
rect 339512 319728 339518 319780
rect 56830 319660 56836 319712
rect 56888 319700 56894 319712
rect 63270 319700 63276 319712
rect 56888 319672 63276 319700
rect 56888 319660 56894 319672
rect 63270 319660 63276 319672
rect 63328 319660 63334 319712
rect 248834 319660 248840 319712
rect 248892 319700 248898 319712
rect 251778 319700 251784 319712
rect 248892 319672 251784 319700
rect 248892 319660 248898 319672
rect 251778 319660 251784 319672
rect 251836 319660 251842 319712
rect 57014 319592 57020 319644
rect 57072 319632 57078 319644
rect 64285 319635 64343 319641
rect 64285 319632 64297 319635
rect 57072 319604 64297 319632
rect 57072 319592 57078 319604
rect 64285 319601 64297 319604
rect 64331 319601 64343 319635
rect 64285 319595 64343 319601
rect 338718 319592 338724 319644
rect 338776 319632 338782 319644
rect 339638 319632 339644 319644
rect 338776 319604 339644 319632
rect 338776 319592 338782 319604
rect 339638 319592 339644 319604
rect 339696 319592 339702 319644
rect 58302 319524 58308 319576
rect 58360 319564 58366 319576
rect 65018 319564 65024 319576
rect 58360 319536 65024 319564
rect 58360 319524 58366 319536
rect 65018 319524 65024 319536
rect 65076 319524 65082 319576
rect 253526 319524 253532 319576
rect 253584 319564 253590 319576
rect 256286 319564 256292 319576
rect 253584 319536 256292 319564
rect 253584 319524 253590 319536
rect 256286 319524 256292 319536
rect 256344 319524 256350 319576
rect 152326 319456 152332 319508
rect 152384 319496 152390 319508
rect 158122 319496 158128 319508
rect 152384 319468 158128 319496
rect 152384 319456 152390 319468
rect 158122 319456 158128 319468
rect 158180 319456 158186 319508
rect 341202 319456 341208 319508
rect 341260 319496 341266 319508
rect 341754 319496 341760 319508
rect 341260 319468 341760 319496
rect 341260 319456 341266 319468
rect 341754 319456 341760 319468
rect 341812 319456 341818 319508
rect 60237 319431 60295 319437
rect 60237 319397 60249 319431
rect 60283 319428 60295 319431
rect 65021 319431 65079 319437
rect 65021 319428 65033 319431
rect 60283 319400 65033 319428
rect 60283 319397 60295 319400
rect 60237 319391 60295 319397
rect 65021 319397 65033 319400
rect 65067 319397 65079 319431
rect 65021 319391 65079 319397
rect 65294 319388 65300 319440
rect 65352 319428 65358 319440
rect 70354 319428 70360 319440
rect 65352 319400 70360 319428
rect 65352 319388 65358 319400
rect 70354 319388 70360 319400
rect 70412 319388 70418 319440
rect 325470 319388 325476 319440
rect 325528 319428 325534 319440
rect 325838 319428 325844 319440
rect 325528 319400 325844 319428
rect 325528 319388 325534 319400
rect 325838 319388 325844 319400
rect 325896 319428 325902 319440
rect 342490 319428 342496 319440
rect 325896 319400 342496 319428
rect 325896 319388 325902 319400
rect 342490 319388 342496 319400
rect 342548 319388 342554 319440
rect 325286 319320 325292 319372
rect 325344 319360 325350 319372
rect 345710 319360 345716 319372
rect 325344 319332 345716 319360
rect 325344 319320 325350 319332
rect 325856 319304 325884 319332
rect 345710 319320 345716 319332
rect 345768 319360 345774 319372
rect 349482 319360 349488 319372
rect 345768 319332 349488 319360
rect 345768 319320 345774 319332
rect 349482 319320 349488 319332
rect 349540 319320 349546 319372
rect 325838 319252 325844 319304
rect 325896 319252 325902 319304
rect 352886 316572 352892 316584
rect 352847 316544 352892 316572
rect 352886 316532 352892 316544
rect 352944 316532 352950 316584
rect 38798 315852 38804 315904
rect 38856 315892 38862 315904
rect 52690 315892 52696 315904
rect 38856 315864 52696 315892
rect 38856 315852 38862 315864
rect 52690 315852 52696 315864
rect 52748 315852 52754 315904
rect 357670 315852 357676 315904
rect 357728 315892 357734 315904
rect 358314 315892 358320 315904
rect 357728 315864 358320 315892
rect 357728 315852 357734 315864
rect 358314 315852 358320 315864
rect 358372 315892 358378 315904
rect 405970 315892 405976 315904
rect 358372 315864 405976 315892
rect 358372 315852 358378 315864
rect 405970 315852 405976 315864
rect 406028 315852 406034 315904
rect 325286 314424 325292 314476
rect 325344 314464 325350 314476
rect 430166 314464 430172 314476
rect 325344 314436 430172 314464
rect 325344 314424 325350 314436
rect 430166 314424 430172 314436
rect 430224 314424 430230 314476
rect 38430 313744 38436 313796
rect 38488 313784 38494 313796
rect 51218 313784 51224 313796
rect 38488 313756 51224 313784
rect 38488 313744 38494 313756
rect 51218 313744 51224 313756
rect 51276 313744 51282 313796
rect 356198 313744 356204 313796
rect 356256 313784 356262 313796
rect 405970 313784 405976 313796
rect 356256 313756 405976 313784
rect 356256 313744 356262 313756
rect 405970 313744 405976 313756
rect 406028 313744 406034 313796
rect 76978 313540 76984 313592
rect 77036 313580 77042 313592
rect 81670 313580 81676 313592
rect 77036 313552 81676 313580
rect 77036 313540 77042 313552
rect 81670 313540 81676 313552
rect 81728 313540 81734 313592
rect 165114 313064 165120 313116
rect 165172 313104 165178 313116
rect 175510 313104 175516 313116
rect 165172 313076 175516 313104
rect 165172 313064 165178 313076
rect 175510 313064 175516 313076
rect 175568 313064 175574 313116
rect 258954 313064 258960 313116
rect 259012 313104 259018 313116
rect 270270 313104 270276 313116
rect 259012 313076 270276 313104
rect 259012 313064 259018 313076
rect 270270 313064 270276 313076
rect 270328 313064 270334 313116
rect 76150 312452 76156 312504
rect 76208 312492 76214 312504
rect 76978 312492 76984 312504
rect 76208 312464 76984 312492
rect 76208 312452 76214 312464
rect 76978 312452 76984 312464
rect 77036 312452 77042 312504
rect 38798 310276 38804 310328
rect 38856 310316 38862 310328
rect 54070 310316 54076 310328
rect 38856 310288 54076 310316
rect 38856 310276 38862 310288
rect 54070 310276 54076 310288
rect 54128 310276 54134 310328
rect 356934 310276 356940 310328
rect 356992 310316 356998 310328
rect 405970 310316 405976 310328
rect 356992 310288 405976 310316
rect 356992 310276 356998 310288
rect 405970 310276 405976 310288
rect 406028 310276 406034 310328
rect 13958 309664 13964 309716
rect 14016 309704 14022 309716
rect 16534 309704 16540 309716
rect 14016 309676 16540 309704
rect 14016 309664 14022 309676
rect 16534 309664 16540 309676
rect 16592 309664 16598 309716
rect 137698 309664 137704 309716
rect 137756 309704 137762 309716
rect 145518 309704 145524 309716
rect 137756 309676 145524 309704
rect 137756 309664 137762 309676
rect 145518 309664 145524 309676
rect 145576 309664 145582 309716
rect 231446 309664 231452 309716
rect 231504 309704 231510 309716
rect 240646 309704 240652 309716
rect 231504 309676 240652 309704
rect 231504 309664 231510 309676
rect 240646 309664 240652 309676
rect 240704 309664 240710 309716
rect 325378 309664 325384 309716
rect 325436 309704 325442 309716
rect 334210 309704 334216 309716
rect 325436 309676 334216 309704
rect 325436 309664 325442 309676
rect 334210 309664 334216 309676
rect 334268 309664 334274 309716
rect 356290 309664 356296 309716
rect 356348 309704 356354 309716
rect 356934 309704 356940 309716
rect 356348 309676 356940 309704
rect 356348 309664 356354 309676
rect 356934 309664 356940 309676
rect 356992 309664 356998 309716
rect 38798 308236 38804 308288
rect 38856 308276 38862 308288
rect 51218 308276 51224 308288
rect 38856 308248 51224 308276
rect 38856 308236 38862 308248
rect 51218 308236 51224 308248
rect 51276 308236 51282 308288
rect 356198 308236 356204 308288
rect 356256 308276 356262 308288
rect 405970 308276 405976 308288
rect 356256 308248 405976 308276
rect 356256 308236 356262 308248
rect 405970 308236 405976 308248
rect 406028 308236 406034 308288
rect 352886 306984 352892 306996
rect 352847 306956 352892 306984
rect 352886 306944 352892 306956
rect 352944 306944 352950 306996
rect 38798 306196 38804 306248
rect 38856 306236 38862 306248
rect 54438 306236 54444 306248
rect 38856 306208 54444 306236
rect 38856 306196 38862 306208
rect 54438 306196 54444 306208
rect 54496 306196 54502 306248
rect 354910 306196 354916 306248
rect 354968 306236 354974 306248
rect 355646 306236 355652 306248
rect 354968 306208 355652 306236
rect 354968 306196 354974 306208
rect 355646 306196 355652 306208
rect 355704 306236 355710 306248
rect 406062 306236 406068 306248
rect 355704 306208 406068 306236
rect 355704 306196 355710 306208
rect 406062 306196 406068 306208
rect 406120 306196 406126 306248
rect 232090 304156 232096 304208
rect 232148 304196 232154 304208
rect 232734 304196 232740 304208
rect 232148 304168 232740 304196
rect 232148 304156 232154 304168
rect 232734 304156 232740 304168
rect 232792 304156 232798 304208
rect 38614 304088 38620 304140
rect 38672 304128 38678 304140
rect 51402 304128 51408 304140
rect 38672 304100 51408 304128
rect 38672 304088 38678 304100
rect 51402 304088 51408 304100
rect 51460 304088 51466 304140
rect 356198 304088 356204 304140
rect 356256 304128 356262 304140
rect 405970 304128 405976 304140
rect 356256 304100 405976 304128
rect 356256 304088 356262 304100
rect 405970 304088 405976 304100
rect 406028 304088 406034 304140
rect 352886 301476 352892 301488
rect 352812 301448 352892 301476
rect 231998 301368 232004 301420
rect 232056 301408 232062 301420
rect 233470 301408 233476 301420
rect 232056 301380 233476 301408
rect 232056 301368 232062 301380
rect 233470 301368 233476 301380
rect 233528 301408 233534 301420
rect 234114 301408 234120 301420
rect 233528 301380 234120 301408
rect 233528 301368 233534 301380
rect 234114 301368 234120 301380
rect 234172 301368 234178 301420
rect 352812 301352 352840 301448
rect 352886 301436 352892 301448
rect 352944 301436 352950 301488
rect 352794 301300 352800 301352
rect 352852 301300 352858 301352
rect 38798 300620 38804 300672
rect 38856 300660 38862 300672
rect 50298 300660 50304 300672
rect 38856 300632 50304 300660
rect 38856 300620 38862 300632
rect 50298 300620 50304 300632
rect 50356 300620 50362 300672
rect 355554 300620 355560 300672
rect 355612 300660 355618 300672
rect 405970 300660 405976 300672
rect 355612 300632 405976 300660
rect 355612 300620 355618 300632
rect 405970 300620 405976 300632
rect 406028 300620 406034 300672
rect 355002 300008 355008 300060
rect 355060 300048 355066 300060
rect 355554 300048 355560 300060
rect 355060 300020 355560 300048
rect 355060 300008 355066 300020
rect 355554 300008 355560 300020
rect 355612 300008 355618 300060
rect 38246 298580 38252 298632
rect 38304 298620 38310 298632
rect 51402 298620 51408 298632
rect 38304 298592 51408 298620
rect 38304 298580 38310 298592
rect 51402 298580 51408 298592
rect 51460 298580 51466 298632
rect 356198 298580 356204 298632
rect 356256 298620 356262 298632
rect 405970 298620 405976 298632
rect 356256 298592 405976 298620
rect 356256 298580 356262 298592
rect 405970 298580 405976 298592
rect 406028 298580 406034 298632
rect 74218 297152 74224 297204
rect 74276 297192 74282 297204
rect 81670 297192 81676 297204
rect 74276 297164 81676 297192
rect 74276 297152 74282 297164
rect 81670 297152 81676 297164
rect 81728 297152 81734 297204
rect 167874 297152 167880 297204
rect 167932 297192 167938 297204
rect 175510 297192 175516 297204
rect 167932 297164 175516 297192
rect 167932 297152 167938 297164
rect 175510 297152 175516 297164
rect 175568 297152 175574 297204
rect 261714 297152 261720 297204
rect 261772 297192 261778 297204
rect 270362 297192 270368 297204
rect 261772 297164 270368 297192
rect 261772 297152 261778 297164
rect 270362 297152 270368 297164
rect 270420 297152 270426 297204
rect 13682 296132 13688 296184
rect 13740 296172 13746 296184
rect 16718 296172 16724 296184
rect 13740 296144 16724 296172
rect 13740 296132 13746 296144
rect 16718 296132 16724 296144
rect 16776 296132 16782 296184
rect 137790 295860 137796 295912
rect 137848 295900 137854 295912
rect 145426 295900 145432 295912
rect 137848 295872 145432 295900
rect 137848 295860 137854 295872
rect 145426 295860 145432 295872
rect 145484 295860 145490 295912
rect 231538 295860 231544 295912
rect 231596 295900 231602 295912
rect 240922 295900 240928 295912
rect 231596 295872 240928 295900
rect 231596 295860 231602 295872
rect 240922 295860 240928 295872
rect 240980 295860 240986 295912
rect 325470 295860 325476 295912
rect 325528 295900 325534 295912
rect 334210 295900 334216 295912
rect 325528 295872 334216 295900
rect 325528 295860 325534 295872
rect 334210 295860 334216 295872
rect 334268 295860 334274 295912
rect 353530 295792 353536 295844
rect 353588 295832 353594 295844
rect 354174 295832 354180 295844
rect 353588 295804 354180 295832
rect 353588 295792 353594 295804
rect 354174 295792 354180 295804
rect 354232 295792 354238 295844
rect 38798 295112 38804 295164
rect 38856 295152 38862 295164
rect 51310 295152 51316 295164
rect 38856 295124 51316 295152
rect 38856 295112 38862 295124
rect 51310 295112 51316 295124
rect 51368 295112 51374 295164
rect 353530 295112 353536 295164
rect 353588 295152 353594 295164
rect 405970 295152 405976 295164
rect 353588 295124 405976 295152
rect 353588 295112 353594 295124
rect 405970 295112 405976 295124
rect 406028 295112 406034 295164
rect 38430 293752 38436 293804
rect 38488 293792 38494 293804
rect 51310 293792 51316 293804
rect 38488 293764 51316 293792
rect 38488 293752 38494 293764
rect 51310 293752 51316 293764
rect 51368 293752 51374 293804
rect 356198 293752 356204 293804
rect 356256 293792 356262 293804
rect 405970 293792 405976 293804
rect 356256 293764 405976 293792
rect 356256 293752 356262 293764
rect 405970 293752 405976 293764
rect 406028 293752 406034 293804
rect 14694 293140 14700 293192
rect 14752 293180 14758 293192
rect 17454 293180 17460 293192
rect 14752 293152 17460 293180
rect 14752 293140 14758 293152
rect 17454 293140 17460 293152
rect 17512 293140 17518 293192
rect 38614 291644 38620 291696
rect 38672 291684 38678 291696
rect 50022 291684 50028 291696
rect 38672 291656 50028 291684
rect 38672 291644 38678 291656
rect 50022 291644 50028 291656
rect 50080 291644 50086 291696
rect 50022 291236 50028 291288
rect 50080 291276 50086 291288
rect 51678 291276 51684 291288
rect 50080 291248 51684 291276
rect 50080 291236 50086 291248
rect 51678 291236 51684 291248
rect 51736 291236 51742 291288
rect 352981 291007 353039 291013
rect 352981 290973 352993 291007
rect 353027 291004 353039 291007
rect 353990 291004 353996 291016
rect 353027 290976 353996 291004
rect 353027 290973 353039 290976
rect 352981 290967 353039 290973
rect 353990 290964 353996 290976
rect 354048 291004 354054 291016
rect 405970 291004 405976 291016
rect 354048 290976 405976 291004
rect 354048 290964 354054 290976
rect 405970 290964 405976 290976
rect 406028 290964 406034 291016
rect 427682 290352 427688 290404
rect 427740 290392 427746 290404
rect 429430 290392 429436 290404
rect 427740 290364 429436 290392
rect 427740 290352 427746 290364
rect 429430 290352 429436 290364
rect 429488 290352 429494 290404
rect 427222 288992 427228 289044
rect 427280 289032 427286 289044
rect 430258 289032 430264 289044
rect 427280 289004 430264 289032
rect 427280 288992 427286 289004
rect 430258 288992 430264 289004
rect 430316 288992 430322 289044
rect 38798 288924 38804 288976
rect 38856 288964 38862 288976
rect 51310 288964 51316 288976
rect 38856 288936 51316 288964
rect 38856 288924 38862 288936
rect 51310 288924 51316 288936
rect 51368 288924 51374 288976
rect 356198 288924 356204 288976
rect 356256 288964 356262 288976
rect 406062 288964 406068 288976
rect 356256 288936 406068 288964
rect 356256 288924 356262 288936
rect 406062 288924 406068 288936
rect 406120 288924 406126 288976
rect 51402 288720 51408 288772
rect 51460 288760 51466 288772
rect 51678 288760 51684 288772
rect 51460 288732 51684 288760
rect 51460 288720 51466 288732
rect 51678 288720 51684 288732
rect 51736 288720 51742 288772
rect 261254 286272 261260 286324
rect 261312 286312 261318 286324
rect 269258 286312 269264 286324
rect 261312 286284 269264 286312
rect 261312 286272 261318 286284
rect 269258 286272 269264 286284
rect 269316 286272 269322 286324
rect 168058 286204 168064 286256
rect 168116 286244 168122 286256
rect 175418 286244 175424 286256
rect 168116 286216 175424 286244
rect 168116 286204 168122 286216
rect 175418 286204 175424 286216
rect 175476 286204 175482 286256
rect 38798 285456 38804 285508
rect 38856 285496 38862 285508
rect 49930 285496 49936 285508
rect 38856 285468 49936 285496
rect 38856 285456 38862 285468
rect 49930 285456 49936 285468
rect 49988 285456 49994 285508
rect 354266 285456 354272 285508
rect 354324 285496 354330 285508
rect 405970 285496 405976 285508
rect 354324 285468 405976 285496
rect 354324 285456 354330 285468
rect 405970 285456 405976 285468
rect 406028 285456 406034 285508
rect 51494 283524 51500 283536
rect 48476 283496 51500 283524
rect 38062 283416 38068 283468
rect 38120 283456 38126 283468
rect 48476 283456 48504 283496
rect 51494 283484 51500 283496
rect 51552 283484 51558 283536
rect 137882 283484 137888 283536
rect 137940 283524 137946 283536
rect 145150 283524 145156 283536
rect 137940 283496 145156 283524
rect 137940 283484 137946 283496
rect 145150 283484 145156 283496
rect 145208 283484 145214 283536
rect 231814 283484 231820 283536
rect 231872 283524 231878 283536
rect 240370 283524 240376 283536
rect 231872 283496 240376 283524
rect 231872 283484 231878 283496
rect 240370 283484 240376 283496
rect 240428 283484 240434 283536
rect 325562 283484 325568 283536
rect 325620 283524 325626 283536
rect 334210 283524 334216 283536
rect 325620 283496 334216 283524
rect 325620 283484 325626 283496
rect 334210 283484 334216 283496
rect 334268 283484 334274 283536
rect 38120 283428 48504 283456
rect 38120 283416 38126 283428
rect 356198 283416 356204 283468
rect 356256 283456 356262 283468
rect 405970 283456 405976 283468
rect 356256 283428 405976 283456
rect 356256 283416 356262 283428
rect 405970 283416 405976 283428
rect 406028 283416 406034 283468
rect 12670 283348 12676 283400
rect 12728 283388 12734 283400
rect 14694 283388 14700 283400
rect 12728 283360 14700 283388
rect 12728 283348 12734 283360
rect 14694 283348 14700 283360
rect 14752 283348 14758 283400
rect 142390 283348 142396 283400
rect 142448 283388 142454 283400
rect 143034 283388 143040 283400
rect 142448 283360 143040 283388
rect 142448 283348 142454 283360
rect 143034 283348 143040 283360
rect 143092 283348 143098 283400
rect 236230 283008 236236 283060
rect 236288 283048 236294 283060
rect 236874 283048 236880 283060
rect 236288 283020 236880 283048
rect 236288 283008 236294 283020
rect 236874 283008 236880 283020
rect 236932 283008 236938 283060
rect 325838 282804 325844 282856
rect 325896 282844 325902 282856
rect 330070 282844 330076 282856
rect 325896 282816 330076 282844
rect 325896 282804 325902 282816
rect 330070 282804 330076 282816
rect 330128 282804 330134 282856
rect 231630 282736 231636 282788
rect 231688 282776 231694 282788
rect 236230 282776 236236 282788
rect 231688 282748 236236 282776
rect 231688 282736 231694 282748
rect 236230 282736 236236 282748
rect 236288 282736 236294 282788
rect 138158 282328 138164 282380
rect 138216 282368 138222 282380
rect 143034 282368 143040 282380
rect 138216 282340 143040 282368
rect 138216 282328 138222 282340
rect 143034 282328 143040 282340
rect 143092 282328 143098 282380
rect 16350 280628 16356 280680
rect 16408 280668 16414 280680
rect 16718 280668 16724 280680
rect 16408 280640 16724 280668
rect 16408 280628 16414 280640
rect 16718 280628 16724 280640
rect 16776 280628 16782 280680
rect 74126 280628 74132 280680
rect 74184 280668 74190 280680
rect 81670 280668 81676 280680
rect 74184 280640 81676 280668
rect 74184 280628 74190 280640
rect 81670 280628 81676 280640
rect 81728 280628 81734 280680
rect 427866 280628 427872 280680
rect 427924 280668 427930 280680
rect 430166 280668 430172 280680
rect 427924 280640 430172 280668
rect 427924 280628 427930 280640
rect 430166 280628 430172 280640
rect 430224 280628 430230 280680
rect 38062 279948 38068 280000
rect 38120 279988 38126 280000
rect 48550 279988 48556 280000
rect 38120 279960 48556 279988
rect 38120 279948 38126 279960
rect 48550 279948 48556 279960
rect 48608 279948 48614 280000
rect 352978 279376 352984 279388
rect 352939 279348 352984 279376
rect 352978 279336 352984 279348
rect 353036 279336 353042 279388
rect 38614 279268 38620 279320
rect 38672 279308 38678 279320
rect 51494 279308 51500 279320
rect 38672 279280 51500 279308
rect 38672 279268 38678 279280
rect 51494 279268 51500 279280
rect 51552 279268 51558 279320
rect 356198 279268 356204 279320
rect 356256 279308 356262 279320
rect 405970 279308 405976 279320
rect 356256 279280 405976 279308
rect 356256 279268 356262 279280
rect 405970 279268 405976 279280
rect 406028 279268 406034 279320
rect 64190 276548 64196 276600
rect 64248 276588 64254 276600
rect 64742 276588 64748 276600
rect 64248 276560 64748 276588
rect 64248 276548 64254 276560
rect 64742 276548 64748 276560
rect 64800 276548 64806 276600
rect 137514 275120 137520 275172
rect 137572 275160 137578 275172
rect 155914 275160 155920 275172
rect 137572 275132 155920 275160
rect 137572 275120 137578 275132
rect 155914 275120 155920 275132
rect 155972 275120 155978 275172
rect 343321 275163 343379 275169
rect 343321 275129 343333 275163
rect 343367 275160 343379 275163
rect 348746 275160 348752 275172
rect 343367 275132 348752 275160
rect 343367 275129 343379 275132
rect 343321 275123 343379 275129
rect 348746 275120 348752 275132
rect 348804 275120 348810 275172
rect 138434 275052 138440 275104
rect 138492 275092 138498 275104
rect 155270 275092 155276 275104
rect 138492 275064 155276 275092
rect 138492 275052 138498 275064
rect 155270 275052 155276 275064
rect 155328 275052 155334 275104
rect 234114 275052 234120 275104
rect 234172 275092 234178 275104
rect 249110 275092 249116 275104
rect 234172 275064 249116 275092
rect 234172 275052 234178 275064
rect 249110 275052 249116 275064
rect 249168 275052 249174 275104
rect 342309 275095 342367 275101
rect 342309 275061 342321 275095
rect 342355 275092 342367 275095
rect 346998 275092 347004 275104
rect 342355 275064 347004 275092
rect 342355 275061 342367 275064
rect 342309 275055 342367 275061
rect 346998 275052 347004 275064
rect 347056 275052 347062 275104
rect 149198 274984 149204 275036
rect 149256 275024 149262 275036
rect 158214 275024 158220 275036
rect 149256 274996 158220 275024
rect 149256 274984 149262 274996
rect 158214 274984 158220 274996
rect 158272 274984 158278 275036
rect 338258 274984 338264 275036
rect 338316 275024 338322 275036
rect 349574 275024 349580 275036
rect 338316 274996 349580 275024
rect 338316 274984 338322 274996
rect 349574 274984 349580 274996
rect 349632 274984 349638 275036
rect 149750 274916 149756 274968
rect 149808 274956 149814 274968
rect 160514 274956 160520 274968
rect 149808 274928 160520 274956
rect 149808 274916 149814 274928
rect 160514 274916 160520 274928
rect 160572 274916 160578 274968
rect 339638 274916 339644 274968
rect 339696 274956 339702 274968
rect 351230 274956 351236 274968
rect 339696 274928 351236 274956
rect 339696 274916 339702 274928
rect 351230 274916 351236 274928
rect 351288 274916 351294 274968
rect 150578 274848 150584 274900
rect 150636 274888 150642 274900
rect 162722 274888 162728 274900
rect 150636 274860 162728 274888
rect 150636 274848 150642 274860
rect 162722 274848 162728 274860
rect 162780 274848 162786 274900
rect 243498 274848 243504 274900
rect 243556 274888 243562 274900
rect 252974 274888 252980 274900
rect 243556 274860 252980 274888
rect 243556 274848 243562 274860
rect 252974 274848 252980 274860
rect 253032 274848 253038 274900
rect 341018 274848 341024 274900
rect 341076 274888 341082 274900
rect 352150 274888 352156 274900
rect 341076 274860 352156 274888
rect 341076 274848 341082 274860
rect 352150 274848 352156 274860
rect 352208 274848 352214 274900
rect 59682 274780 59688 274832
rect 59740 274820 59746 274832
rect 60786 274820 60792 274832
rect 59740 274792 60792 274820
rect 59740 274780 59746 274792
rect 60786 274780 60792 274792
rect 60844 274780 60850 274832
rect 151866 274780 151872 274832
rect 151924 274820 151930 274832
rect 163274 274820 163280 274832
rect 151924 274792 163280 274820
rect 151924 274780 151930 274792
rect 163274 274780 163280 274792
rect 163332 274780 163338 274832
rect 244050 274780 244056 274832
rect 244108 274820 244114 274832
rect 254446 274820 254452 274832
rect 244108 274792 254452 274820
rect 244108 274780 244114 274792
rect 254446 274780 254452 274792
rect 254504 274780 254510 274832
rect 336878 274780 336884 274832
rect 336936 274820 336942 274832
rect 343321 274823 343379 274829
rect 343321 274820 343333 274823
rect 336936 274792 343333 274820
rect 336936 274780 336942 274792
rect 343321 274789 343333 274792
rect 343367 274789 343379 274823
rect 346170 274820 346176 274832
rect 343321 274783 343379 274789
rect 343428 274792 346176 274820
rect 34566 274712 34572 274764
rect 34624 274752 34630 274764
rect 46986 274752 46992 274764
rect 34624 274724 46992 274752
rect 34624 274712 34630 274724
rect 46986 274712 46992 274724
rect 47044 274712 47050 274764
rect 149198 274712 149204 274764
rect 149256 274752 149262 274764
rect 162078 274752 162084 274764
rect 149256 274724 162084 274752
rect 149256 274712 149262 274724
rect 162078 274712 162084 274724
rect 162136 274712 162142 274764
rect 243038 274712 243044 274764
rect 243096 274752 243102 274764
rect 255734 274752 255740 274764
rect 243096 274724 255740 274752
rect 243096 274712 243102 274724
rect 255734 274712 255740 274724
rect 255792 274712 255798 274764
rect 334118 274712 334124 274764
rect 334176 274752 334182 274764
rect 343428 274752 343456 274792
rect 346170 274780 346176 274792
rect 346228 274780 346234 274832
rect 334176 274724 343456 274752
rect 334176 274712 334182 274724
rect 343502 274712 343508 274764
rect 343560 274752 343566 274764
rect 348194 274752 348200 274764
rect 343560 274724 348200 274752
rect 343560 274712 343566 274724
rect 348194 274712 348200 274724
rect 348252 274712 348258 274764
rect 31898 274644 31904 274696
rect 31956 274684 31962 274696
rect 46618 274684 46624 274696
rect 31956 274656 46624 274684
rect 31956 274644 31962 274656
rect 46618 274644 46624 274656
rect 46676 274644 46682 274696
rect 147818 274644 147824 274696
rect 147876 274684 147882 274696
rect 161434 274684 161440 274696
rect 147876 274656 161440 274684
rect 147876 274644 147882 274656
rect 161434 274644 161440 274656
rect 161492 274644 161498 274696
rect 241658 274644 241664 274696
rect 241716 274684 241722 274696
rect 255090 274684 255096 274696
rect 241716 274656 255096 274684
rect 241716 274644 241722 274656
rect 255090 274644 255096 274656
rect 255148 274644 255154 274696
rect 335406 274644 335412 274696
rect 335464 274684 335470 274696
rect 342309 274687 342367 274693
rect 342309 274684 342321 274687
rect 335464 274656 342321 274684
rect 335464 274644 335470 274656
rect 342309 274653 342321 274656
rect 342355 274653 342367 274687
rect 342309 274647 342367 274653
rect 342398 274644 342404 274696
rect 342456 274684 342462 274696
rect 345894 274684 345900 274696
rect 342456 274656 345900 274684
rect 342456 274644 342462 274656
rect 345894 274644 345900 274656
rect 345952 274644 345958 274696
rect 29230 274576 29236 274628
rect 29288 274616 29294 274628
rect 46526 274616 46532 274628
rect 29288 274588 46532 274616
rect 29288 274576 29294 274588
rect 46526 274576 46532 274588
rect 46584 274576 46590 274628
rect 145058 274576 145064 274628
rect 145116 274616 145122 274628
rect 160238 274616 160244 274628
rect 145116 274588 160244 274616
rect 145116 274576 145122 274588
rect 160238 274576 160244 274588
rect 160296 274576 160302 274628
rect 240278 274576 240284 274628
rect 240336 274616 240342 274628
rect 254538 274616 254544 274628
rect 240336 274588 254544 274616
rect 240336 274576 240342 274588
rect 254538 274576 254544 274588
rect 254596 274576 254602 274628
rect 332738 274576 332744 274628
rect 332796 274616 332802 274628
rect 332796 274588 341708 274616
rect 332796 274576 332802 274588
rect 26562 274508 26568 274560
rect 26620 274548 26626 274560
rect 47078 274548 47084 274560
rect 26620 274520 47084 274548
rect 26620 274508 26626 274520
rect 47078 274508 47084 274520
rect 47136 274508 47142 274560
rect 146438 274508 146444 274560
rect 146496 274548 146502 274560
rect 160882 274548 160888 274560
rect 146496 274520 160888 274548
rect 146496 274508 146502 274520
rect 160882 274508 160888 274520
rect 160940 274508 160946 274560
rect 238898 274508 238904 274560
rect 238956 274548 238962 274560
rect 254170 274548 254176 274560
rect 238956 274520 254176 274548
rect 238956 274508 238962 274520
rect 254170 274508 254176 274520
rect 254228 274508 254234 274560
rect 335498 274508 335504 274560
rect 335556 274548 335562 274560
rect 335556 274520 341156 274548
rect 335556 274508 335562 274520
rect 23894 274440 23900 274492
rect 23952 274480 23958 274492
rect 46434 274480 46440 274492
rect 23952 274452 46440 274480
rect 23952 274440 23958 274452
rect 46434 274440 46440 274452
rect 46492 274440 46498 274492
rect 57014 274440 57020 274492
rect 57072 274480 57078 274492
rect 68054 274480 68060 274492
rect 57072 274452 68060 274480
rect 57072 274440 57078 274452
rect 68054 274440 68060 274452
rect 68112 274440 68118 274492
rect 143678 274440 143684 274492
rect 143736 274480 143742 274492
rect 159594 274480 159600 274492
rect 143736 274452 159600 274480
rect 143736 274440 143742 274452
rect 159594 274440 159600 274452
rect 159652 274440 159658 274492
rect 237518 274440 237524 274492
rect 237576 274480 237582 274492
rect 253250 274480 253256 274492
rect 237576 274452 253256 274480
rect 237576 274440 237582 274452
rect 253250 274440 253256 274452
rect 253308 274440 253314 274492
rect 246534 274236 246540 274288
rect 246592 274276 246598 274288
rect 247178 274276 247184 274288
rect 246592 274248 247184 274276
rect 246592 274236 246598 274248
rect 247178 274236 247184 274248
rect 247236 274236 247242 274288
rect 341128 274276 341156 274520
rect 341680 274412 341708 274588
rect 344330 274576 344336 274628
rect 344388 274616 344394 274628
rect 349574 274616 349580 274628
rect 344388 274588 349580 274616
rect 344388 274576 344394 274588
rect 349574 274576 349580 274588
rect 349632 274576 349638 274628
rect 341754 274508 341760 274560
rect 341812 274548 341818 274560
rect 345986 274548 345992 274560
rect 341812 274520 345992 274548
rect 341812 274508 341818 274520
rect 345986 274508 345992 274520
rect 346044 274508 346050 274560
rect 345158 274440 345164 274492
rect 345216 274480 345222 274492
rect 367974 274480 367980 274492
rect 345216 274452 367980 274480
rect 345216 274440 345222 274452
rect 367974 274440 367980 274452
rect 368032 274440 368038 274492
rect 369906 274440 369912 274492
rect 369964 274480 369970 274492
rect 410202 274480 410208 274492
rect 369964 274452 410208 274480
rect 369964 274440 369970 274452
rect 410202 274440 410208 274452
rect 410260 274440 410266 274492
rect 345342 274412 345348 274424
rect 341680 274384 345348 274412
rect 345342 274372 345348 274384
rect 345400 274372 345406 274424
rect 348010 274276 348016 274288
rect 341128 274248 348016 274276
rect 348010 274236 348016 274248
rect 348068 274236 348074 274288
rect 338166 274032 338172 274084
rect 338224 274072 338230 274084
rect 342582 274072 342588 274084
rect 338224 274044 342588 274072
rect 338224 274032 338230 274044
rect 342582 274032 342588 274044
rect 342640 274032 342646 274084
rect 62350 273964 62356 274016
rect 62408 274004 62414 274016
rect 63638 274004 63644 274016
rect 62408 273976 63644 274004
rect 62408 273964 62414 273976
rect 63638 273964 63644 273976
rect 63696 273964 63702 274016
rect 247270 273964 247276 274016
rect 247328 274004 247334 274016
rect 247822 274004 247828 274016
rect 247328 273976 247828 274004
rect 247328 273964 247334 273976
rect 247822 273964 247828 273976
rect 247880 274004 247886 274016
rect 249570 274004 249576 274016
rect 247880 273976 249576 274004
rect 247880 273964 247886 273976
rect 249570 273964 249576 273976
rect 249628 273964 249634 274016
rect 339270 273964 339276 274016
rect 339328 274004 339334 274016
rect 341938 274004 341944 274016
rect 339328 273976 341944 274004
rect 339328 273964 339334 273976
rect 341938 273964 341944 273976
rect 341996 273964 342002 274016
rect 254814 273896 254820 273948
rect 254872 273936 254878 273948
rect 257574 273936 257580 273948
rect 254872 273908 257580 273936
rect 254872 273896 254878 273908
rect 257574 273896 257580 273908
rect 257632 273896 257638 273948
rect 337614 273896 337620 273948
rect 337672 273936 337678 273948
rect 341110 273936 341116 273948
rect 337672 273908 341116 273936
rect 337672 273896 337678 273908
rect 341110 273896 341116 273908
rect 341168 273896 341174 273948
rect 61614 273828 61620 273880
rect 61672 273868 61678 273880
rect 63270 273868 63276 273880
rect 61672 273840 63276 273868
rect 61672 273828 61678 273840
rect 63270 273828 63276 273840
rect 63328 273828 63334 273880
rect 64374 273828 64380 273880
rect 64432 273868 64438 273880
rect 65938 273868 65944 273880
rect 64432 273840 65944 273868
rect 64432 273828 64438 273840
rect 65938 273828 65944 273840
rect 65996 273828 66002 273880
rect 151038 273828 151044 273880
rect 151096 273868 151102 273880
rect 151958 273868 151964 273880
rect 151096 273840 151964 273868
rect 151096 273828 151102 273840
rect 151958 273828 151964 273840
rect 152016 273828 152022 273880
rect 234114 273828 234120 273880
rect 234172 273868 234178 273880
rect 234758 273868 234764 273880
rect 234172 273840 234764 273868
rect 234172 273828 234178 273840
rect 234758 273828 234764 273840
rect 234816 273828 234822 273880
rect 256194 273828 256200 273880
rect 256252 273868 256258 273880
rect 258310 273868 258316 273880
rect 256252 273840 258316 273868
rect 256252 273828 256258 273840
rect 258310 273828 258316 273840
rect 258368 273828 258374 273880
rect 340098 273828 340104 273880
rect 340156 273868 340162 273880
rect 341846 273868 341852 273880
rect 340156 273840 341852 273868
rect 340156 273828 340162 273840
rect 341846 273828 341852 273840
rect 341904 273828 341910 273880
rect 21226 273760 21232 273812
rect 21284 273800 21290 273812
rect 22238 273800 22244 273812
rect 21284 273772 22244 273800
rect 21284 273760 21290 273772
rect 22238 273760 22244 273772
rect 22296 273760 22302 273812
rect 61430 273760 61436 273812
rect 61488 273800 61494 273812
rect 62258 273800 62264 273812
rect 61488 273772 62264 273800
rect 61488 273760 61494 273772
rect 62258 273760 62264 273772
rect 62316 273760 62322 273812
rect 62994 273760 63000 273812
rect 63052 273800 63058 273812
rect 64098 273800 64104 273812
rect 63052 273772 64104 273800
rect 63052 273760 63058 273772
rect 64098 273760 64104 273772
rect 64156 273760 64162 273812
rect 65754 273760 65760 273812
rect 65812 273800 65818 273812
rect 66766 273800 66772 273812
rect 65812 273772 66772 273800
rect 65812 273760 65818 273772
rect 66766 273760 66772 273772
rect 66824 273760 66830 273812
rect 68514 273760 68520 273812
rect 68572 273800 68578 273812
rect 69434 273800 69440 273812
rect 68572 273772 69440 273800
rect 68572 273760 68578 273772
rect 69434 273760 69440 273772
rect 69492 273760 69498 273812
rect 152234 273760 152240 273812
rect 152292 273800 152298 273812
rect 153246 273800 153252 273812
rect 152292 273772 153252 273800
rect 152292 273760 152298 273772
rect 153246 273760 153252 273772
rect 153304 273760 153310 273812
rect 153430 273760 153436 273812
rect 153488 273800 153494 273812
rect 153488 273772 154764 273800
rect 153488 273760 153494 273772
rect 154736 273744 154764 273772
rect 162354 273760 162360 273812
rect 162412 273800 162418 273812
rect 163918 273800 163924 273812
rect 162412 273772 163924 273800
rect 162412 273760 162418 273772
rect 163918 273760 163924 273772
rect 163976 273760 163982 273812
rect 245338 273760 245344 273812
rect 245396 273800 245402 273812
rect 245798 273800 245804 273812
rect 245396 273772 245804 273800
rect 245396 273760 245402 273772
rect 245798 273760 245804 273772
rect 245856 273760 245862 273812
rect 247730 273760 247736 273812
rect 247788 273800 247794 273812
rect 248466 273800 248472 273812
rect 247788 273772 248472 273800
rect 247788 273760 247794 273772
rect 248466 273760 248472 273772
rect 248524 273760 248530 273812
rect 249018 273760 249024 273812
rect 249076 273800 249082 273812
rect 249938 273800 249944 273812
rect 249076 273772 249944 273800
rect 249076 273760 249082 273772
rect 249938 273760 249944 273772
rect 249996 273760 250002 273812
rect 256286 273760 256292 273812
rect 256344 273800 256350 273812
rect 256930 273800 256936 273812
rect 256344 273772 256936 273800
rect 256344 273760 256350 273772
rect 256930 273760 256936 273772
rect 256988 273760 256994 273812
rect 340926 273760 340932 273812
rect 340984 273800 340990 273812
rect 341754 273800 341760 273812
rect 340984 273772 341760 273800
rect 340984 273760 340990 273772
rect 341754 273760 341760 273772
rect 341812 273760 341818 273812
rect 154718 273692 154724 273744
rect 154776 273692 154782 273744
rect 352794 272400 352800 272452
rect 352852 272440 352858 272452
rect 352978 272440 352984 272452
rect 352852 272412 352984 272440
rect 352852 272400 352858 272412
rect 352978 272400 352984 272412
rect 353036 272400 353042 272452
rect 349482 271720 349488 271772
rect 349540 271760 349546 271772
rect 350402 271760 350408 271772
rect 349540 271732 350408 271760
rect 349540 271720 349546 271732
rect 350402 271720 350408 271732
rect 350460 271720 350466 271772
rect 12854 270020 12860 270072
rect 12912 270060 12918 270072
rect 16442 270060 16448 270072
rect 12912 270032 16448 270060
rect 12912 270020 12918 270032
rect 16442 270020 16448 270032
rect 16500 270020 16506 270072
rect 88386 269612 88392 269664
rect 88444 269652 88450 269664
rect 182410 269652 182416 269664
rect 88444 269624 182416 269652
rect 88444 269612 88450 269624
rect 182410 269612 182416 269624
rect 182468 269652 182474 269664
rect 182962 269652 182968 269664
rect 182468 269624 182968 269652
rect 182468 269612 182474 269624
rect 182962 269612 182968 269624
rect 183020 269652 183026 269664
rect 276434 269652 276440 269664
rect 183020 269624 276440 269652
rect 183020 269612 183026 269624
rect 276434 269612 276440 269624
rect 276492 269612 276498 269664
rect 290694 269612 290700 269664
rect 290752 269652 290758 269664
rect 430074 269652 430080 269664
rect 290752 269624 430080 269652
rect 290752 269612 290758 269624
rect 430074 269612 430080 269624
rect 430132 269612 430138 269664
rect 13314 269544 13320 269596
rect 13372 269584 13378 269596
rect 95470 269584 95476 269596
rect 13372 269556 95476 269584
rect 13372 269544 13378 269556
rect 95470 269544 95476 269556
rect 95528 269584 95534 269596
rect 96758 269584 96764 269596
rect 95528 269556 96764 269584
rect 95528 269544 95534 269556
rect 96758 269544 96764 269556
rect 96816 269544 96822 269596
rect 102646 269544 102652 269596
rect 102704 269584 102710 269596
rect 196670 269584 196676 269596
rect 102704 269556 196676 269584
rect 102704 269544 102710 269556
rect 196670 269544 196676 269556
rect 196728 269544 196734 269596
rect 189402 269476 189408 269528
rect 189460 269516 189466 269528
rect 283518 269516 283524 269528
rect 189460 269488 283524 269516
rect 189460 269476 189466 269488
rect 283518 269476 283524 269488
rect 283576 269476 283582 269528
rect 127762 269340 127768 269392
rect 127820 269380 127826 269392
rect 131166 269380 131172 269392
rect 127820 269352 131172 269380
rect 127820 269340 127826 269352
rect 131166 269340 131172 269352
rect 131224 269340 131230 269392
rect 303758 269340 303764 269392
rect 303816 269380 303822 269392
rect 304954 269380 304960 269392
rect 303816 269352 304960 269380
rect 303816 269340 303822 269352
rect 304954 269340 304960 269352
rect 305012 269340 305018 269392
rect 310750 269340 310756 269392
rect 310808 269380 310814 269392
rect 312038 269380 312044 269392
rect 310808 269352 312044 269380
rect 310808 269340 310814 269352
rect 312038 269340 312044 269352
rect 312096 269340 312102 269392
rect 95562 269000 95568 269052
rect 95620 269040 95626 269052
rect 109730 269040 109736 269052
rect 95620 269012 109736 269040
rect 95620 269000 95626 269012
rect 109730 269000 109736 269012
rect 109788 269000 109794 269052
rect 189310 269000 189316 269052
rect 189368 269040 189374 269052
rect 203754 269040 203760 269052
rect 189368 269012 203760 269040
rect 189368 269000 189374 269012
rect 203754 269000 203760 269012
rect 203812 269000 203818 269052
rect 284530 269000 284536 269052
rect 284588 269040 284594 269052
rect 297778 269040 297784 269052
rect 284588 269012 297784 269040
rect 284588 269000 284594 269012
rect 297778 269000 297784 269012
rect 297836 269000 297842 269052
rect 96758 268932 96764 268984
rect 96816 268972 96822 268984
rect 170634 268972 170640 268984
rect 96816 268944 170640 268972
rect 96816 268932 96822 268944
rect 170634 268932 170640 268944
rect 170692 268972 170698 268984
rect 189402 268972 189408 268984
rect 170692 268944 189408 268972
rect 170692 268932 170698 268944
rect 189402 268932 189408 268944
rect 189460 268932 189466 268984
rect 196670 268932 196676 268984
rect 196728 268972 196734 268984
rect 268614 268972 268620 268984
rect 196728 268944 268620 268972
rect 196728 268932 196734 268944
rect 268614 268932 268620 268944
rect 268672 268972 268678 268984
rect 290694 268972 290700 268984
rect 268672 268944 290700 268972
rect 268672 268932 268678 268944
rect 290694 268932 290700 268944
rect 290752 268932 290758 268984
rect 210010 268864 210016 268916
rect 210068 268904 210074 268916
rect 210930 268904 210936 268916
rect 210068 268876 210936 268904
rect 210068 268864 210074 268876
rect 210930 268864 210936 268876
rect 210988 268864 210994 268916
rect 114790 268524 114796 268576
rect 114848 268564 114854 268576
rect 116906 268564 116912 268576
rect 114848 268536 116912 268564
rect 114848 268524 114854 268536
rect 116906 268524 116912 268536
rect 116964 268524 116970 268576
rect 354910 267844 354916 267896
rect 354968 267884 354974 267896
rect 355830 267884 355836 267896
rect 354968 267856 355836 267884
rect 354968 267844 354974 267856
rect 355830 267844 355836 267856
rect 355888 267844 355894 267896
rect 64834 266824 64840 266876
rect 64892 266864 64898 266876
rect 68514 266864 68520 266876
rect 64892 266836 68520 266864
rect 64892 266824 64898 266836
rect 68514 266824 68520 266836
rect 68572 266824 68578 266876
rect 158214 266824 158220 266876
rect 158272 266864 158278 266876
rect 158950 266864 158956 266876
rect 158272 266836 158956 266864
rect 158272 266824 158278 266836
rect 158950 266824 158956 266836
rect 159008 266824 159014 266876
rect 247638 266824 247644 266876
rect 247696 266864 247702 266876
rect 254814 266864 254820 266876
rect 247696 266836 254820 266864
rect 247696 266824 247702 266836
rect 254814 266824 254820 266836
rect 254872 266824 254878 266876
rect 153154 266756 153160 266808
rect 153212 266796 153218 266808
rect 162354 266796 162360 266808
rect 153212 266768 162360 266796
rect 153212 266756 153218 266768
rect 162354 266756 162360 266768
rect 162412 266756 162418 266808
rect 246258 266756 246264 266808
rect 246316 266796 246322 266808
rect 256286 266796 256292 266808
rect 246316 266768 256292 266796
rect 246316 266756 246322 266768
rect 256286 266756 256292 266768
rect 256344 266756 256350 266808
rect 59682 266688 59688 266740
rect 59740 266728 59746 266740
rect 63822 266728 63828 266740
rect 59740 266700 63828 266728
rect 59740 266688 59746 266700
rect 63822 266688 63828 266700
rect 63880 266688 63886 266740
rect 154718 266688 154724 266740
rect 154776 266728 154782 266740
rect 164470 266728 164476 266740
rect 154776 266700 164476 266728
rect 154776 266688 154782 266700
rect 164470 266688 164476 266700
rect 164528 266688 164534 266740
rect 244878 266688 244884 266740
rect 244936 266728 244942 266740
rect 255642 266728 255648 266740
rect 244936 266700 255648 266728
rect 244936 266688 244942 266700
rect 255642 266688 255648 266700
rect 255700 266688 255706 266740
rect 63638 266620 63644 266672
rect 63696 266660 63702 266672
rect 75230 266660 75236 266672
rect 63696 266632 75236 266660
rect 63696 266620 63702 266632
rect 75230 266620 75236 266632
rect 75288 266620 75294 266672
rect 151958 266620 151964 266672
rect 152016 266660 152022 266672
rect 156837 266663 156895 266669
rect 156837 266660 156849 266663
rect 152016 266632 156849 266660
rect 152016 266620 152022 266632
rect 156837 266629 156849 266632
rect 156883 266629 156895 266663
rect 161710 266660 161716 266672
rect 156837 266623 156895 266629
rect 156944 266632 161716 266660
rect 62258 266552 62264 266604
rect 62316 266592 62322 266604
rect 74218 266592 74224 266604
rect 62316 266564 74224 266592
rect 62316 266552 62322 266564
rect 74218 266552 74224 266564
rect 74276 266552 74282 266604
rect 150486 266552 150492 266604
rect 150544 266592 150550 266604
rect 156944 266592 156972 266632
rect 161710 266620 161716 266632
rect 161768 266620 161774 266672
rect 245798 266620 245804 266672
rect 245856 266660 245862 266672
rect 256930 266660 256936 266672
rect 245856 266632 256936 266660
rect 245856 266620 245862 266632
rect 256930 266620 256936 266632
rect 256988 266620 256994 266672
rect 150544 266564 156972 266592
rect 150544 266552 150550 266564
rect 244418 266552 244424 266604
rect 244476 266592 244482 266604
rect 255550 266592 255556 266604
rect 244476 266564 255556 266592
rect 244476 266552 244482 266564
rect 255550 266552 255556 266564
rect 255608 266552 255614 266604
rect 60878 266484 60884 266536
rect 60936 266524 60942 266536
rect 73114 266524 73120 266536
rect 60936 266496 73120 266524
rect 60936 266484 60942 266496
rect 73114 266484 73120 266496
rect 73172 266484 73178 266536
rect 143034 266484 143040 266536
rect 143092 266524 143098 266536
rect 155730 266524 155736 266536
rect 143092 266496 155736 266524
rect 143092 266484 143098 266496
rect 155730 266484 155736 266496
rect 155788 266484 155794 266536
rect 247178 266484 247184 266536
rect 247236 266524 247242 266536
rect 259690 266524 259696 266536
rect 247236 266496 259696 266524
rect 247236 266484 247242 266496
rect 259690 266484 259696 266496
rect 259748 266484 259754 266536
rect 341754 266484 341760 266536
rect 341812 266524 341818 266536
rect 345802 266524 345808 266536
rect 341812 266496 345808 266524
rect 341812 266484 341818 266496
rect 345802 266484 345808 266496
rect 345860 266484 345866 266536
rect 59498 266416 59504 266468
rect 59556 266456 59562 266468
rect 71090 266456 71096 266468
rect 59556 266428 71096 266456
rect 59556 266416 59562 266428
rect 71090 266416 71096 266428
rect 71148 266416 71154 266468
rect 153246 266416 153252 266468
rect 153304 266456 153310 266468
rect 165942 266456 165948 266468
rect 153304 266428 165948 266456
rect 153304 266416 153310 266428
rect 165942 266416 165948 266428
rect 166000 266416 166006 266468
rect 245706 266416 245712 266468
rect 245764 266456 245770 266468
rect 258402 266456 258408 266468
rect 245764 266428 258408 266456
rect 245764 266416 245770 266428
rect 258402 266416 258408 266428
rect 258460 266416 258466 266468
rect 58118 266348 58124 266400
rect 58176 266388 58182 266400
rect 70078 266388 70084 266400
rect 58176 266360 70084 266388
rect 58176 266348 58182 266360
rect 70078 266348 70084 266360
rect 70136 266348 70142 266400
rect 151774 266348 151780 266400
rect 151832 266388 151838 266400
rect 164562 266388 164568 266400
rect 151832 266360 164568 266388
rect 151832 266348 151838 266360
rect 164562 266348 164568 266360
rect 164620 266348 164626 266400
rect 236874 266348 236880 266400
rect 236932 266388 236938 266400
rect 250030 266388 250036 266400
rect 236932 266360 250036 266388
rect 236932 266348 236938 266360
rect 250030 266348 250036 266360
rect 250088 266348 250094 266400
rect 56738 266280 56744 266332
rect 56796 266320 56802 266332
rect 67962 266320 67968 266332
rect 56796 266292 67968 266320
rect 56796 266280 56802 266292
rect 67962 266280 67968 266292
rect 68020 266280 68026 266332
rect 154626 266280 154632 266332
rect 154684 266320 154690 266332
rect 168702 266320 168708 266332
rect 154684 266292 168708 266320
rect 154684 266280 154690 266292
rect 168702 266280 168708 266292
rect 168760 266280 168766 266332
rect 248466 266280 248472 266332
rect 248524 266320 248530 266332
rect 262450 266320 262456 266332
rect 248524 266292 262456 266320
rect 248524 266280 248530 266292
rect 262450 266280 262456 266292
rect 262508 266280 262514 266332
rect 55358 266212 55364 266264
rect 55416 266252 55422 266264
rect 66950 266252 66956 266264
rect 55416 266224 66956 266252
rect 55416 266212 55422 266224
rect 66950 266212 66956 266224
rect 67008 266212 67014 266264
rect 153338 266212 153344 266264
rect 153396 266252 153402 266264
rect 167322 266252 167328 266264
rect 153396 266224 167328 266252
rect 153396 266212 153402 266224
rect 167322 266212 167328 266224
rect 167380 266212 167386 266264
rect 247086 266212 247092 266264
rect 247144 266252 247150 266264
rect 261070 266252 261076 266264
rect 247144 266224 261076 266252
rect 247144 266212 247150 266224
rect 261070 266212 261076 266224
rect 261128 266212 261134 266264
rect 60786 266144 60792 266196
rect 60844 266184 60850 266196
rect 72102 266184 72108 266196
rect 60844 266156 72108 266184
rect 60844 266144 60850 266156
rect 72102 266144 72108 266156
rect 72160 266144 72166 266196
rect 154534 266144 154540 266196
rect 154592 266184 154598 266196
rect 170082 266184 170088 266196
rect 154592 266156 170088 266184
rect 154592 266144 154598 266156
rect 170082 266144 170088 266156
rect 170140 266144 170146 266196
rect 248558 266144 248564 266196
rect 248616 266184 248622 266196
rect 263830 266184 263836 266196
rect 248616 266156 263836 266184
rect 248616 266144 248622 266156
rect 263830 266144 263836 266156
rect 263888 266144 263894 266196
rect 338534 266144 338540 266196
rect 338592 266184 338598 266196
rect 349482 266184 349488 266196
rect 338592 266156 349488 266184
rect 338592 266144 338598 266156
rect 349482 266144 349488 266156
rect 349540 266144 349546 266196
rect 156837 266119 156895 266125
rect 156837 266085 156849 266119
rect 156883 266116 156895 266119
rect 163090 266116 163096 266128
rect 156883 266088 163096 266116
rect 156883 266085 156895 266088
rect 156837 266079 156895 266085
rect 163090 266076 163096 266088
rect 163148 266076 163154 266128
rect 63822 266008 63828 266060
rect 63880 266048 63886 266060
rect 67870 266048 67876 266060
rect 63880 266020 67876 266048
rect 63880 266008 63886 266020
rect 67870 266008 67876 266020
rect 67928 266008 67934 266060
rect 60694 265804 60700 265856
rect 60752 265844 60758 265856
rect 64374 265844 64380 265856
rect 60752 265816 64380 265844
rect 60752 265804 60758 265816
rect 64374 265804 64380 265816
rect 64432 265804 64438 265856
rect 62810 265736 62816 265788
rect 62868 265776 62874 265788
rect 66490 265776 66496 265788
rect 62868 265748 66496 265776
rect 62868 265736 62874 265748
rect 66490 265736 66496 265748
rect 66548 265736 66554 265788
rect 61798 265668 61804 265720
rect 61856 265708 61862 265720
rect 65754 265708 65760 265720
rect 61856 265680 65760 265708
rect 61856 265668 61862 265680
rect 65754 265668 65760 265680
rect 65812 265668 65818 265720
rect 157846 265668 157852 265720
rect 157904 265708 157910 265720
rect 165114 265708 165120 265720
rect 157904 265680 165120 265708
rect 157904 265668 157910 265680
rect 165114 265668 165120 265680
rect 165172 265668 165178 265720
rect 251870 265668 251876 265720
rect 251928 265708 251934 265720
rect 258954 265708 258960 265720
rect 251928 265680 258960 265708
rect 251928 265668 251934 265680
rect 258954 265668 258960 265680
rect 259012 265668 259018 265720
rect 58670 265600 58676 265652
rect 58728 265640 58734 265652
rect 62994 265640 63000 265652
rect 58728 265612 63000 265640
rect 58728 265600 58734 265612
rect 62994 265600 63000 265612
rect 63052 265600 63058 265652
rect 341846 265600 341852 265652
rect 341904 265640 341910 265652
rect 344790 265640 344796 265652
rect 341904 265612 344796 265640
rect 341904 265600 341910 265612
rect 344790 265600 344796 265612
rect 344848 265600 344854 265652
rect 345894 265600 345900 265652
rect 345952 265640 345958 265652
rect 347918 265640 347924 265652
rect 345952 265612 347924 265640
rect 345952 265600 345958 265612
rect 347918 265600 347924 265612
rect 347976 265600 347982 265652
rect 57658 265532 57664 265584
rect 57716 265572 57722 265584
rect 61614 265572 61620 265584
rect 57716 265544 61620 265572
rect 57716 265532 57722 265544
rect 61614 265532 61620 265544
rect 61672 265532 61678 265584
rect 65938 265532 65944 265584
rect 65996 265572 66002 265584
rect 69250 265572 69256 265584
rect 65996 265544 69256 265572
rect 65996 265532 66002 265544
rect 69250 265532 69256 265544
rect 69308 265532 69314 265584
rect 249018 265532 249024 265584
rect 249076 265572 249082 265584
rect 256194 265572 256200 265584
rect 249076 265544 256200 265572
rect 249076 265532 249082 265544
rect 256194 265532 256200 265544
rect 256252 265532 256258 265584
rect 333382 265532 333388 265584
rect 333440 265572 333446 265584
rect 334118 265572 334124 265584
rect 333440 265544 334124 265572
rect 333440 265532 333446 265544
rect 334118 265532 334124 265544
rect 334176 265532 334182 265584
rect 334394 265532 334400 265584
rect 334452 265572 334458 265584
rect 335406 265572 335412 265584
rect 334452 265544 335412 265572
rect 334452 265532 334458 265544
rect 335406 265532 335412 265544
rect 335464 265532 335470 265584
rect 341938 265532 341944 265584
rect 341996 265572 342002 265584
rect 343778 265572 343784 265584
rect 341996 265544 343784 265572
rect 341996 265532 342002 265544
rect 343778 265532 343784 265544
rect 343836 265532 343842 265584
rect 345986 265532 345992 265584
rect 346044 265572 346050 265584
rect 346814 265572 346820 265584
rect 346044 265544 346820 265572
rect 346044 265532 346050 265544
rect 346814 265532 346820 265544
rect 346872 265532 346878 265584
rect 427590 265464 427596 265516
rect 427648 265504 427654 265516
rect 429430 265504 429436 265516
rect 427648 265476 429436 265504
rect 427648 265464 427654 265476
rect 429430 265464 429436 265476
rect 429488 265464 429494 265516
rect 51310 265056 51316 265108
rect 51368 265096 51374 265108
rect 52046 265096 52052 265108
rect 51368 265068 52052 265096
rect 51368 265056 51374 265068
rect 52046 265056 52052 265068
rect 52104 265056 52110 265108
rect 74034 264416 74040 264428
rect 73995 264388 74040 264416
rect 74034 264376 74040 264388
rect 74092 264376 74098 264428
rect 78910 264036 78916 264088
rect 78968 264076 78974 264088
rect 123254 264076 123260 264088
rect 78968 264048 123260 264076
rect 78968 264036 78974 264048
rect 123254 264036 123260 264048
rect 123312 264076 123318 264088
rect 124358 264076 124364 264088
rect 123312 264048 124364 264076
rect 123312 264036 123318 264048
rect 124358 264036 124364 264048
rect 124416 264036 124422 264088
rect 310750 264036 310756 264088
rect 310808 264076 310814 264088
rect 328414 264076 328420 264088
rect 310808 264048 328420 264076
rect 310808 264036 310814 264048
rect 328414 264036 328420 264048
rect 328472 264036 328478 264088
rect 267234 263492 267240 263544
rect 267292 263532 267298 263544
rect 310750 263532 310756 263544
rect 267292 263504 310756 263532
rect 267292 263492 267298 263504
rect 310750 263492 310756 263504
rect 310808 263492 310814 263544
rect 73942 263464 73948 263476
rect 73903 263436 73948 263464
rect 73942 263424 73948 263436
rect 74000 263424 74006 263476
rect 124358 263424 124364 263476
rect 124416 263464 124422 263476
rect 140274 263464 140280 263476
rect 124416 263436 140280 263464
rect 124416 263424 124422 263436
rect 140274 263424 140280 263436
rect 140332 263424 140338 263476
rect 249938 263424 249944 263476
rect 249996 263464 250002 263476
rect 358406 263464 358412 263476
rect 249996 263436 358412 263464
rect 249996 263424 250002 263436
rect 358406 263424 358412 263436
rect 358464 263424 358470 263476
rect 74037 263399 74095 263405
rect 74037 263365 74049 263399
rect 74083 263396 74095 263399
rect 369538 263396 369544 263408
rect 74083 263368 369544 263396
rect 74083 263365 74095 263368
rect 74037 263359 74095 263365
rect 369538 263356 369544 263368
rect 369596 263356 369602 263408
rect 225834 262880 225840 262932
rect 225892 262920 225898 262932
rect 233470 262920 233476 262932
rect 225892 262892 233476 262920
rect 225892 262880 225898 262892
rect 233470 262880 233476 262892
rect 233528 262880 233534 262932
rect 131994 262744 132000 262796
rect 132052 262784 132058 262796
rect 139814 262784 139820 262796
rect 132052 262756 139820 262784
rect 132052 262744 132058 262756
rect 139814 262744 139820 262756
rect 139872 262744 139878 262796
rect 325194 262744 325200 262796
rect 325252 262784 325258 262796
rect 325838 262784 325844 262796
rect 325252 262756 325844 262784
rect 325252 262744 325258 262756
rect 325838 262744 325844 262756
rect 325896 262784 325902 262796
rect 360706 262784 360712 262796
rect 325896 262756 360712 262784
rect 325896 262744 325902 262756
rect 360706 262744 360712 262756
rect 360764 262744 360770 262796
rect 46986 262676 46992 262728
rect 47044 262716 47050 262728
rect 49194 262716 49200 262728
rect 47044 262688 49200 262716
rect 47044 262676 47050 262688
rect 49194 262676 49200 262688
rect 49252 262716 49258 262728
rect 73945 262719 74003 262725
rect 73945 262716 73957 262719
rect 49252 262688 73957 262716
rect 49252 262676 49258 262688
rect 73945 262685 73957 262688
rect 73991 262685 74003 262719
rect 73945 262679 74003 262685
rect 228686 262608 228692 262660
rect 228744 262648 228750 262660
rect 369722 262648 369728 262660
rect 228744 262620 369728 262648
rect 228744 262608 228750 262620
rect 369722 262608 369728 262620
rect 369780 262608 369786 262660
rect 13406 262540 13412 262592
rect 13464 262580 13470 262592
rect 385270 262580 385276 262592
rect 13464 262552 385276 262580
rect 13464 262540 13470 262552
rect 385270 262540 385276 262552
rect 385328 262540 385334 262592
rect 360430 261996 360436 262048
rect 360488 262036 360494 262048
rect 360798 262036 360804 262048
rect 360488 262008 360804 262036
rect 360488 261996 360494 262008
rect 360798 261996 360804 262008
rect 360856 262036 360862 262048
rect 422530 262036 422536 262048
rect 360856 262008 422536 262036
rect 360856 261996 360862 262008
rect 422530 261996 422536 262008
rect 422588 261996 422594 262048
rect 78910 261384 78916 261436
rect 78968 261424 78974 261436
rect 87190 261424 87196 261436
rect 78968 261396 87196 261424
rect 78968 261384 78974 261396
rect 87190 261384 87196 261396
rect 87248 261384 87254 261436
rect 132086 261384 132092 261436
rect 132144 261424 132150 261436
rect 140366 261424 140372 261436
rect 132144 261396 140372 261424
rect 132144 261384 132150 261396
rect 140366 261384 140372 261396
rect 140424 261384 140430 261436
rect 225742 261384 225748 261436
rect 225800 261424 225806 261436
rect 233470 261424 233476 261436
rect 225800 261396 233476 261424
rect 225800 261384 225806 261396
rect 233470 261384 233476 261396
rect 233528 261384 233534 261436
rect 324642 261384 324648 261436
rect 324700 261424 324706 261436
rect 327678 261424 327684 261436
rect 324700 261396 327684 261424
rect 324700 261384 324706 261396
rect 327678 261384 327684 261396
rect 327736 261384 327742 261436
rect 95562 261316 95568 261368
rect 95620 261356 95626 261368
rect 96206 261356 96212 261368
rect 95620 261328 96212 261356
rect 95620 261316 95626 261328
rect 96206 261316 96212 261328
rect 96264 261316 96270 261368
rect 203846 261248 203852 261300
rect 203904 261288 203910 261300
rect 209918 261288 209924 261300
rect 203904 261260 209924 261288
rect 203904 261248 203910 261260
rect 209918 261248 209924 261260
rect 209976 261248 209982 261300
rect 297870 261248 297876 261300
rect 297928 261288 297934 261300
rect 303758 261288 303764 261300
rect 297928 261260 303764 261288
rect 297928 261248 297934 261260
rect 303758 261248 303764 261260
rect 303816 261248 303822 261300
rect 217186 260636 217192 260688
rect 217244 260676 217250 260688
rect 225190 260676 225196 260688
rect 217244 260648 225196 260676
rect 217244 260636 217250 260648
rect 225190 260636 225196 260648
rect 225248 260636 225254 260688
rect 311210 260636 311216 260688
rect 311268 260676 311274 260688
rect 319214 260676 319220 260688
rect 311268 260648 319220 260676
rect 311268 260636 311274 260648
rect 319214 260636 319220 260648
rect 319272 260636 319278 260688
rect 123530 260568 123536 260620
rect 123588 260608 123594 260620
rect 127762 260608 127768 260620
rect 123588 260580 127768 260608
rect 123588 260568 123594 260580
rect 127762 260568 127768 260580
rect 127820 260568 127826 260620
rect 110190 260432 110196 260484
rect 110248 260472 110254 260484
rect 114790 260472 114796 260484
rect 110248 260444 114796 260472
rect 110248 260432 110254 260444
rect 114790 260432 114796 260444
rect 114848 260432 114854 260484
rect 78910 260024 78916 260076
rect 78968 260064 78974 260076
rect 85074 260064 85080 260076
rect 78968 260036 85080 260064
rect 78968 260024 78974 260036
rect 85074 260024 85080 260036
rect 85132 260024 85138 260076
rect 132454 260024 132460 260076
rect 132512 260064 132518 260076
rect 140366 260064 140372 260076
rect 132512 260036 140372 260064
rect 132512 260024 132518 260036
rect 140366 260024 140372 260036
rect 140424 260024 140430 260076
rect 189310 260024 189316 260076
rect 189368 260064 189374 260076
rect 190506 260064 190512 260076
rect 189368 260036 190512 260064
rect 189368 260024 189374 260036
rect 190506 260024 190512 260036
rect 190564 260024 190570 260076
rect 226202 260024 226208 260076
rect 226260 260064 226266 260076
rect 233470 260064 233476 260076
rect 226260 260036 233476 260064
rect 226260 260024 226266 260036
rect 233470 260024 233476 260036
rect 233528 260024 233534 260076
rect 360614 259276 360620 259328
rect 360672 259316 360678 259328
rect 419770 259316 419776 259328
rect 360672 259288 419776 259316
rect 360672 259276 360678 259288
rect 419770 259276 419776 259288
rect 419828 259276 419834 259328
rect 78910 258664 78916 258716
rect 78968 258704 78974 258716
rect 84430 258704 84436 258716
rect 78968 258676 84436 258704
rect 78968 258664 78974 258676
rect 84430 258664 84436 258676
rect 84488 258664 84494 258716
rect 132178 258596 132184 258648
rect 132236 258636 132242 258648
rect 140550 258636 140556 258648
rect 132236 258608 140556 258636
rect 132236 258596 132242 258608
rect 140550 258596 140556 258608
rect 140608 258596 140614 258648
rect 226294 258596 226300 258648
rect 226352 258636 226358 258648
rect 233470 258636 233476 258648
rect 226352 258608 233476 258636
rect 226352 258596 226358 258608
rect 233470 258596 233476 258608
rect 233528 258596 233534 258648
rect 321054 258528 321060 258580
rect 321112 258568 321118 258580
rect 324642 258568 324648 258580
rect 321112 258540 324648 258568
rect 321112 258528 321118 258540
rect 324642 258528 324648 258540
rect 324700 258528 324706 258580
rect 78910 257304 78916 257356
rect 78968 257344 78974 257356
rect 81670 257344 81676 257356
rect 78968 257316 81676 257344
rect 78968 257304 78974 257316
rect 81670 257304 81676 257316
rect 81728 257304 81734 257356
rect 132270 257304 132276 257356
rect 132328 257344 132334 257356
rect 140550 257344 140556 257356
rect 132328 257316 140556 257344
rect 132328 257304 132334 257316
rect 140550 257304 140556 257316
rect 140608 257304 140614 257356
rect 226478 257304 226484 257356
rect 226536 257344 226542 257356
rect 232826 257344 232832 257356
rect 226536 257316 232832 257344
rect 226536 257304 226542 257316
rect 232826 257304 232832 257316
rect 232884 257304 232890 257356
rect 131350 257236 131356 257288
rect 131408 257276 131414 257288
rect 140642 257276 140648 257288
rect 131408 257248 140648 257276
rect 131408 257236 131414 257248
rect 140642 257236 140648 257248
rect 140700 257236 140706 257288
rect 173118 257236 173124 257288
rect 173176 257276 173182 257288
rect 181030 257276 181036 257288
rect 173176 257248 181036 257276
rect 173176 257236 173182 257248
rect 181030 257236 181036 257248
rect 181088 257236 181094 257288
rect 226110 257236 226116 257288
rect 226168 257276 226174 257288
rect 233470 257276 233476 257288
rect 226168 257248 233476 257276
rect 226168 257236 226174 257248
rect 233470 257236 233476 257248
rect 233528 257236 233534 257288
rect 321054 257168 321060 257220
rect 321112 257208 321118 257220
rect 327954 257208 327960 257220
rect 321112 257180 327960 257208
rect 321112 257168 321118 257180
rect 327954 257168 327960 257180
rect 328012 257168 328018 257220
rect 85074 256828 85080 256880
rect 85132 256868 85138 256880
rect 87190 256868 87196 256880
rect 85132 256840 87196 256868
rect 85132 256828 85138 256840
rect 87190 256828 87196 256840
rect 87248 256828 87254 256880
rect 12854 256556 12860 256608
rect 12912 256596 12918 256608
rect 16258 256596 16264 256608
rect 12912 256568 16264 256596
rect 12912 256556 12918 256568
rect 16258 256556 16264 256568
rect 16316 256556 16322 256608
rect 361166 256488 361172 256540
rect 361224 256528 361230 256540
rect 417010 256528 417016 256540
rect 361224 256500 417016 256528
rect 361224 256488 361230 256500
rect 417010 256488 417016 256500
rect 417068 256488 417074 256540
rect 78910 255876 78916 255928
rect 78968 255916 78974 255928
rect 81762 255916 81768 255928
rect 78968 255888 81768 255916
rect 78968 255876 78974 255888
rect 81762 255876 81768 255888
rect 81820 255876 81826 255928
rect 132362 255876 132368 255928
rect 132420 255916 132426 255928
rect 139722 255916 139728 255928
rect 132420 255888 139728 255916
rect 132420 255876 132426 255888
rect 139722 255876 139728 255888
rect 139780 255876 139786 255928
rect 173302 255876 173308 255928
rect 173360 255916 173366 255928
rect 176154 255916 176160 255928
rect 173360 255888 176160 255916
rect 173360 255876 173366 255888
rect 176154 255876 176160 255888
rect 176212 255876 176218 255928
rect 178270 255876 178276 255928
rect 178328 255916 178334 255928
rect 181030 255916 181036 255928
rect 178328 255888 181036 255916
rect 178328 255876 178334 255888
rect 181030 255876 181036 255888
rect 181088 255876 181094 255928
rect 228686 255876 228692 255928
rect 228744 255916 228750 255928
rect 233470 255916 233476 255928
rect 228744 255888 233476 255916
rect 228744 255876 228750 255888
rect 233470 255876 233476 255888
rect 233528 255876 233534 255928
rect 266590 255876 266596 255928
rect 266648 255916 266654 255928
rect 271374 255916 271380 255928
rect 266648 255888 271380 255916
rect 266648 255876 266654 255888
rect 271374 255876 271380 255888
rect 271432 255876 271438 255928
rect 81670 255808 81676 255860
rect 81728 255848 81734 255860
rect 87190 255848 87196 255860
rect 81728 255820 87196 255848
rect 81728 255808 81734 255820
rect 87190 255808 87196 255820
rect 87248 255808 87254 255860
rect 320594 255808 320600 255860
rect 320652 255848 320658 255860
rect 327126 255848 327132 255860
rect 320652 255820 327132 255848
rect 320652 255808 320658 255820
rect 327126 255808 327132 255820
rect 327184 255808 327190 255860
rect 84430 255740 84436 255792
rect 84488 255780 84494 255792
rect 87282 255780 87288 255792
rect 84488 255752 87288 255780
rect 84488 255740 84494 255752
rect 87282 255740 87288 255752
rect 87340 255740 87346 255792
rect 321606 255740 321612 255792
rect 321664 255780 321670 255792
rect 327218 255780 327224 255792
rect 321664 255752 327224 255780
rect 321664 255740 321670 255752
rect 327218 255740 327224 255752
rect 327276 255740 327282 255792
rect 173578 255536 173584 255588
rect 173636 255576 173642 255588
rect 222706 255576 222712 255588
rect 173636 255548 222712 255576
rect 173636 255536 173642 255548
rect 222706 255536 222712 255548
rect 222764 255536 222770 255588
rect 225834 255128 225840 255180
rect 225892 255128 225898 255180
rect 225926 255128 225932 255180
rect 225984 255168 225990 255180
rect 234574 255168 234580 255180
rect 225984 255140 234580 255168
rect 225984 255128 225990 255140
rect 234574 255128 234580 255140
rect 234632 255128 234638 255180
rect 225852 254976 225880 255128
rect 225834 254924 225840 254976
rect 225892 254924 225898 254976
rect 131350 254584 131356 254636
rect 131408 254624 131414 254636
rect 136134 254624 136140 254636
rect 131408 254596 136140 254624
rect 131408 254584 131414 254596
rect 136134 254584 136140 254596
rect 136192 254584 136198 254636
rect 131994 254516 132000 254568
rect 132052 254556 132058 254568
rect 136226 254556 136232 254568
rect 132052 254528 136232 254556
rect 132052 254516 132058 254528
rect 136226 254516 136232 254528
rect 136284 254516 136290 254568
rect 176338 254516 176344 254568
rect 176396 254556 176402 254568
rect 181030 254556 181036 254568
rect 176396 254528 181036 254556
rect 176396 254516 176402 254528
rect 181030 254516 181036 254528
rect 181088 254516 181094 254568
rect 266590 254516 266596 254568
rect 266648 254556 266654 254568
rect 272754 254556 272760 254568
rect 266648 254528 272760 254556
rect 266648 254516 266654 254528
rect 272754 254516 272760 254528
rect 272812 254516 272818 254568
rect 78910 254448 78916 254500
rect 78968 254488 78974 254500
rect 82682 254488 82688 254500
rect 78968 254460 82688 254488
rect 78968 254448 78974 254460
rect 82682 254448 82688 254460
rect 82740 254448 82746 254500
rect 132546 254448 132552 254500
rect 132604 254488 132610 254500
rect 140550 254488 140556 254500
rect 132604 254460 140556 254488
rect 132604 254448 132610 254460
rect 140550 254448 140556 254460
rect 140608 254448 140614 254500
rect 173302 254448 173308 254500
rect 173360 254488 173366 254500
rect 176246 254488 176252 254500
rect 173360 254460 176252 254488
rect 173360 254448 173366 254460
rect 176246 254448 176252 254460
rect 176304 254448 176310 254500
rect 179190 254448 179196 254500
rect 179248 254488 179254 254500
rect 181582 254488 181588 254500
rect 179248 254460 181588 254488
rect 179248 254448 179254 254460
rect 181582 254448 181588 254460
rect 181640 254448 181646 254500
rect 267878 254448 267884 254500
rect 267936 254488 267942 254500
rect 274870 254488 274876 254500
rect 267936 254460 274876 254488
rect 267936 254448 267942 254460
rect 274870 254448 274876 254460
rect 274928 254448 274934 254500
rect 320502 254448 320508 254500
rect 320560 254488 320566 254500
rect 328414 254488 328420 254500
rect 320560 254460 328420 254488
rect 320560 254448 320566 254460
rect 328414 254448 328420 254460
rect 328472 254448 328478 254500
rect 81762 254380 81768 254432
rect 81820 254420 81826 254432
rect 87190 254420 87196 254432
rect 81820 254392 87196 254420
rect 81820 254380 81826 254392
rect 87190 254380 87196 254392
rect 87248 254380 87254 254432
rect 321606 253904 321612 253956
rect 321664 253944 321670 253956
rect 328506 253944 328512 253956
rect 321664 253916 328512 253944
rect 321664 253904 321670 253916
rect 328506 253904 328512 253916
rect 328564 253904 328570 253956
rect 179006 253428 179012 253480
rect 179064 253468 179070 253480
rect 181030 253468 181036 253480
rect 179064 253440 181036 253468
rect 179064 253428 179070 253440
rect 181030 253428 181036 253440
rect 181088 253428 181094 253480
rect 225742 253360 225748 253412
rect 225800 253400 225806 253412
rect 234206 253400 234212 253412
rect 225800 253372 234212 253400
rect 225800 253360 225806 253372
rect 234206 253360 234212 253372
rect 234264 253360 234270 253412
rect 131350 253156 131356 253208
rect 131408 253196 131414 253208
rect 137698 253196 137704 253208
rect 131408 253168 137704 253196
rect 131408 253156 131414 253168
rect 137698 253156 137704 253168
rect 137756 253156 137762 253208
rect 230066 253156 230072 253208
rect 230124 253196 230130 253208
rect 233470 253196 233476 253208
rect 230124 253168 233476 253196
rect 230124 253156 230130 253168
rect 233470 253156 233476 253168
rect 233528 253156 233534 253208
rect 78910 253088 78916 253140
rect 78968 253128 78974 253140
rect 78968 253100 84476 253128
rect 78968 253088 78974 253100
rect 84448 252992 84476 253100
rect 137514 253088 137520 253140
rect 137572 253128 137578 253140
rect 139814 253128 139820 253140
rect 137572 253100 139820 253128
rect 137572 253088 137578 253100
rect 139814 253088 139820 253100
rect 139872 253088 139878 253140
rect 266590 253088 266596 253140
rect 266648 253128 266654 253140
rect 272846 253128 272852 253140
rect 266648 253100 272852 253128
rect 266648 253088 266654 253100
rect 272846 253088 272852 253100
rect 272904 253088 272910 253140
rect 361166 253020 361172 253072
rect 361224 253060 361230 253072
rect 414250 253060 414256 253072
rect 361224 253032 414256 253060
rect 361224 253020 361230 253032
rect 414250 253020 414256 253032
rect 414308 253020 414314 253072
rect 427498 253020 427504 253072
rect 427556 253060 427562 253072
rect 429430 253060 429436 253072
rect 427556 253032 429436 253060
rect 427556 253020 427562 253032
rect 429430 253020 429436 253032
rect 429488 253020 429494 253072
rect 87282 252992 87288 253004
rect 84448 252964 87288 252992
rect 87282 252952 87288 252964
rect 87340 252952 87346 253004
rect 82682 252884 82688 252936
rect 82740 252924 82746 252936
rect 87190 252924 87196 252936
rect 82740 252896 87196 252924
rect 82740 252884 82746 252896
rect 87190 252884 87196 252896
rect 87248 252884 87254 252936
rect 132270 252408 132276 252460
rect 132328 252408 132334 252460
rect 132288 252256 132316 252408
rect 267326 252340 267332 252392
rect 267384 252380 267390 252392
rect 267786 252380 267792 252392
rect 267384 252352 267792 252380
rect 267384 252340 267390 252352
rect 267786 252340 267792 252352
rect 267844 252340 267850 252392
rect 132270 252204 132276 252256
rect 132328 252204 132334 252256
rect 174038 251864 174044 251916
rect 174096 251904 174102 251916
rect 178914 251904 178920 251916
rect 174096 251876 178920 251904
rect 174096 251864 174102 251876
rect 178914 251864 178920 251876
rect 178972 251864 178978 251916
rect 275974 251904 275980 251916
rect 271392 251876 275980 251904
rect 131350 251796 131356 251848
rect 131408 251836 131414 251848
rect 138986 251836 138992 251848
rect 131408 251808 138992 251836
rect 131408 251796 131414 251808
rect 138986 251796 138992 251808
rect 139044 251796 139050 251848
rect 78910 251728 78916 251780
rect 78968 251768 78974 251780
rect 78968 251740 84476 251768
rect 78968 251728 78974 251740
rect 84448 251632 84476 251740
rect 132638 251728 132644 251780
rect 132696 251768 132702 251780
rect 140550 251768 140556 251780
rect 132696 251740 140556 251768
rect 132696 251728 132702 251740
rect 140550 251728 140556 251740
rect 140608 251728 140614 251780
rect 174038 251728 174044 251780
rect 174096 251768 174102 251780
rect 181582 251768 181588 251780
rect 174096 251740 181588 251768
rect 174096 251728 174102 251740
rect 181582 251728 181588 251740
rect 181640 251728 181646 251780
rect 230158 251728 230164 251780
rect 230216 251768 230222 251780
rect 233562 251768 233568 251780
rect 230216 251740 233568 251768
rect 230216 251728 230222 251740
rect 233562 251728 233568 251740
rect 233620 251728 233626 251780
rect 266590 251728 266596 251780
rect 266648 251768 266654 251780
rect 271392 251768 271420 251876
rect 275974 251864 275980 251876
rect 276032 251864 276038 251916
rect 321606 251864 321612 251916
rect 321664 251904 321670 251916
rect 327126 251904 327132 251916
rect 321664 251876 327132 251904
rect 321664 251864 321670 251876
rect 327126 251864 327132 251876
rect 327184 251864 327190 251916
rect 266648 251740 271420 251768
rect 266648 251728 266654 251740
rect 271466 251728 271472 251780
rect 271524 251768 271530 251780
rect 274870 251768 274876 251780
rect 271524 251740 274876 251768
rect 271524 251728 271530 251740
rect 274870 251728 274876 251740
rect 274928 251728 274934 251780
rect 87190 251632 87196 251644
rect 84448 251604 87196 251632
rect 87190 251592 87196 251604
rect 87248 251592 87254 251644
rect 222798 250980 222804 251032
rect 222856 251020 222862 251032
rect 233470 251020 233476 251032
rect 222856 250992 233476 251020
rect 222856 250980 222862 250992
rect 233470 250980 233476 250992
rect 233528 250980 233534 251032
rect 321606 250980 321612 251032
rect 321664 251020 321670 251032
rect 327218 251020 327224 251032
rect 321664 250992 327224 251020
rect 321664 250980 321670 250992
rect 327218 250980 327224 250992
rect 327276 250980 327282 251032
rect 79738 250300 79744 250352
rect 79796 250340 79802 250352
rect 87190 250340 87196 250352
rect 79796 250312 87196 250340
rect 79796 250300 79802 250312
rect 87190 250300 87196 250312
rect 87248 250300 87254 250352
rect 173578 250300 173584 250352
rect 173636 250340 173642 250352
rect 182318 250340 182324 250352
rect 173636 250312 182324 250340
rect 173636 250300 173642 250312
rect 182318 250300 182324 250312
rect 182376 250300 182382 250352
rect 173486 250232 173492 250284
rect 173544 250272 173550 250284
rect 181490 250272 181496 250284
rect 173544 250244 181496 250272
rect 173544 250232 173550 250244
rect 181490 250232 181496 250244
rect 181548 250232 181554 250284
rect 266590 250232 266596 250284
rect 266648 250272 266654 250284
rect 276158 250272 276164 250284
rect 266648 250244 276164 250272
rect 266648 250232 266654 250244
rect 276158 250232 276164 250244
rect 276216 250232 276222 250284
rect 267418 250164 267424 250216
rect 267476 250204 267482 250216
rect 274870 250204 274876 250216
rect 267476 250176 274876 250204
rect 267476 250164 267482 250176
rect 274870 250164 274876 250176
rect 274928 250164 274934 250216
rect 78910 249552 78916 249604
rect 78968 249592 78974 249604
rect 87190 249592 87196 249604
rect 78968 249564 87196 249592
rect 78968 249552 78974 249564
rect 87190 249552 87196 249564
rect 87248 249552 87254 249604
rect 360706 249552 360712 249604
rect 360764 249592 360770 249604
rect 412870 249592 412876 249604
rect 360764 249564 412876 249592
rect 360764 249552 360770 249564
rect 412870 249552 412876 249564
rect 412928 249552 412934 249604
rect 321054 249484 321060 249536
rect 321112 249524 321118 249536
rect 327218 249524 327224 249536
rect 321112 249496 327224 249524
rect 321112 249484 321118 249496
rect 327218 249484 327224 249496
rect 327276 249484 327282 249536
rect 321606 249076 321612 249128
rect 321664 249116 321670 249128
rect 328414 249116 328420 249128
rect 321664 249088 328420 249116
rect 321664 249076 321670 249088
rect 328414 249076 328420 249088
rect 328472 249076 328478 249128
rect 131994 248940 132000 248992
rect 132052 248980 132058 248992
rect 138894 248980 138900 248992
rect 132052 248952 138900 248980
rect 132052 248940 132058 248952
rect 138894 248940 138900 248952
rect 138952 248940 138958 248992
rect 225834 248940 225840 248992
rect 225892 248980 225898 248992
rect 234114 248980 234120 248992
rect 225892 248952 234120 248980
rect 225892 248940 225898 248952
rect 234114 248940 234120 248952
rect 234172 248940 234178 248992
rect 173394 248872 173400 248924
rect 173452 248912 173458 248924
rect 181950 248912 181956 248924
rect 173452 248884 181956 248912
rect 173452 248872 173458 248884
rect 181950 248872 181956 248884
rect 182008 248872 182014 248924
rect 226570 248872 226576 248924
rect 226628 248912 226634 248924
rect 233470 248912 233476 248924
rect 226628 248884 233476 248912
rect 226628 248872 226634 248884
rect 233470 248872 233476 248884
rect 233528 248872 233534 248924
rect 266590 248872 266596 248924
rect 266648 248912 266654 248924
rect 274962 248912 274968 248924
rect 266648 248884 274968 248912
rect 266648 248872 266654 248884
rect 274962 248872 274968 248884
rect 275020 248872 275026 248924
rect 173762 248804 173768 248856
rect 173820 248844 173826 248856
rect 181858 248844 181864 248856
rect 173820 248816 181864 248844
rect 173820 248804 173826 248816
rect 181858 248804 181864 248816
rect 181916 248804 181922 248856
rect 267510 248804 267516 248856
rect 267568 248844 267574 248856
rect 274870 248844 274876 248856
rect 267568 248816 274876 248844
rect 267568 248804 267574 248816
rect 274870 248804 274876 248816
rect 274928 248804 274934 248856
rect 267602 248736 267608 248788
rect 267660 248776 267666 248788
rect 274962 248776 274968 248788
rect 267660 248748 274968 248776
rect 267660 248736 267666 248748
rect 274962 248736 274968 248748
rect 275020 248736 275026 248788
rect 173486 248668 173492 248720
rect 173544 248708 173550 248720
rect 178270 248708 178276 248720
rect 173544 248680 178276 248708
rect 173544 248668 173550 248680
rect 178270 248668 178276 248680
rect 178328 248668 178334 248720
rect 78910 248192 78916 248244
rect 78968 248232 78974 248244
rect 87190 248232 87196 248244
rect 78968 248204 87196 248232
rect 78968 248192 78974 248204
rect 87190 248192 87196 248204
rect 87248 248192 87254 248244
rect 321606 247648 321612 247700
rect 321664 247688 321670 247700
rect 328414 247688 328420 247700
rect 321664 247660 328420 247688
rect 321664 247648 321670 247660
rect 328414 247648 328420 247660
rect 328472 247648 328478 247700
rect 78910 247512 78916 247564
rect 78968 247552 78974 247564
rect 88478 247552 88484 247564
rect 78968 247524 88484 247552
rect 78968 247512 78974 247524
rect 88478 247512 88484 247524
rect 88536 247512 88542 247564
rect 173854 247512 173860 247564
rect 173912 247552 173918 247564
rect 182318 247552 182324 247564
rect 173912 247524 182324 247552
rect 173912 247512 173918 247524
rect 182318 247512 182324 247524
rect 182376 247512 182382 247564
rect 267786 247512 267792 247564
rect 267844 247552 267850 247564
rect 274870 247552 274876 247564
rect 267844 247524 274876 247552
rect 267844 247512 267850 247524
rect 274870 247512 274876 247524
rect 274928 247512 274934 247564
rect 321790 247512 321796 247564
rect 321848 247552 321854 247564
rect 328414 247552 328420 247564
rect 321848 247524 328420 247552
rect 321848 247512 321854 247524
rect 328414 247512 328420 247524
rect 328472 247512 328478 247564
rect 136226 247240 136232 247292
rect 136284 247280 136290 247292
rect 140642 247280 140648 247292
rect 136284 247252 140648 247280
rect 136284 247240 136290 247252
rect 140642 247240 140648 247252
rect 140700 247240 140706 247292
rect 173302 246492 173308 246544
rect 173360 246532 173366 246544
rect 179190 246532 179196 246544
rect 173360 246504 179196 246532
rect 173360 246492 173366 246504
rect 179190 246492 179196 246504
rect 179248 246492 179254 246544
rect 321422 246220 321428 246272
rect 321480 246260 321486 246272
rect 321480 246232 321836 246260
rect 321480 246220 321486 246232
rect 78910 246152 78916 246204
rect 78968 246192 78974 246204
rect 87190 246192 87196 246204
rect 78968 246164 87196 246192
rect 78968 246152 78974 246164
rect 87190 246152 87196 246164
rect 87248 246152 87254 246204
rect 131350 246152 131356 246204
rect 131408 246192 131414 246204
rect 131408 246164 135996 246192
rect 131408 246152 131414 246164
rect 135968 246124 135996 246164
rect 136134 246152 136140 246204
rect 136192 246192 136198 246204
rect 140366 246192 140372 246204
rect 136192 246164 140372 246192
rect 136192 246152 136198 246164
rect 140366 246152 140372 246164
rect 140424 246152 140430 246204
rect 172750 246152 172756 246204
rect 172808 246192 172814 246204
rect 176338 246192 176344 246204
rect 172808 246164 176344 246192
rect 172808 246152 172814 246164
rect 176338 246152 176344 246164
rect 176396 246152 176402 246204
rect 176433 246195 176491 246201
rect 176433 246161 176445 246195
rect 176479 246192 176491 246195
rect 182318 246192 182324 246204
rect 176479 246164 182324 246192
rect 176479 246161 176491 246164
rect 176433 246155 176491 246161
rect 182318 246152 182324 246164
rect 182376 246152 182382 246204
rect 226386 246152 226392 246204
rect 226444 246192 226450 246204
rect 233470 246192 233476 246204
rect 226444 246164 233476 246192
rect 226444 246152 226450 246164
rect 233470 246152 233476 246164
rect 233528 246152 233534 246204
rect 267694 246152 267700 246204
rect 267752 246192 267758 246204
rect 274870 246192 274876 246204
rect 267752 246164 274876 246192
rect 267752 246152 267758 246164
rect 274870 246152 274876 246164
rect 274928 246152 274934 246204
rect 321808 246192 321836 246232
rect 327862 246192 327868 246204
rect 321808 246164 327868 246192
rect 327862 246152 327868 246164
rect 327920 246152 327926 246204
rect 140550 246124 140556 246136
rect 135968 246096 140556 246124
rect 140550 246084 140556 246096
rect 140608 246084 140614 246136
rect 176154 246084 176160 246136
rect 176212 246124 176218 246136
rect 181582 246124 181588 246136
rect 176212 246096 181588 246124
rect 176212 246084 176218 246096
rect 181582 246084 181588 246096
rect 181640 246084 181646 246136
rect 266590 246084 266596 246136
rect 266648 246124 266654 246136
rect 275790 246124 275796 246136
rect 266648 246096 275796 246124
rect 266648 246084 266654 246096
rect 275790 246084 275796 246096
rect 275848 246084 275854 246136
rect 173670 246016 173676 246068
rect 173728 246056 173734 246068
rect 176433 246059 176491 246065
rect 176433 246056 176445 246059
rect 173728 246028 176445 246056
rect 173728 246016 173734 246028
rect 176433 246025 176445 246028
rect 176479 246025 176491 246059
rect 176433 246019 176491 246025
rect 271374 246016 271380 246068
rect 271432 246056 271438 246068
rect 274962 246056 274968 246068
rect 271432 246028 274968 246056
rect 271432 246016 271438 246028
rect 274962 246016 274968 246028
rect 275020 246016 275026 246068
rect 225558 245200 225564 245252
rect 225616 245240 225622 245252
rect 228686 245240 228692 245252
rect 225616 245212 228692 245240
rect 225616 245200 225622 245212
rect 228686 245200 228692 245212
rect 228744 245200 228750 245252
rect 321698 244860 321704 244912
rect 321756 244900 321762 244912
rect 323170 244900 323176 244912
rect 321756 244872 323176 244900
rect 321756 244860 321762 244872
rect 323170 244860 323176 244872
rect 323228 244860 323234 244912
rect 321606 244792 321612 244844
rect 321664 244832 321670 244844
rect 321664 244804 321836 244832
rect 321664 244792 321670 244804
rect 78910 244724 78916 244776
rect 78968 244764 78974 244776
rect 87190 244764 87196 244776
rect 78968 244736 87196 244764
rect 78968 244724 78974 244736
rect 87190 244724 87196 244736
rect 87248 244724 87254 244776
rect 137698 244724 137704 244776
rect 137756 244764 137762 244776
rect 140090 244764 140096 244776
rect 137756 244736 140096 244764
rect 137756 244724 137762 244736
rect 140090 244724 140096 244736
rect 140148 244724 140154 244776
rect 176246 244724 176252 244776
rect 176304 244764 176310 244776
rect 182318 244764 182324 244776
rect 176304 244736 182324 244764
rect 176304 244724 176310 244736
rect 182318 244724 182324 244736
rect 182376 244724 182382 244776
rect 225558 244724 225564 244776
rect 225616 244764 225622 244776
rect 232734 244764 232740 244776
rect 225616 244736 232740 244764
rect 225616 244724 225622 244736
rect 232734 244724 232740 244736
rect 232792 244724 232798 244776
rect 266590 244724 266596 244776
rect 266648 244764 266654 244776
rect 266648 244736 271972 244764
rect 266648 244724 266654 244736
rect 271944 244628 271972 244736
rect 272754 244724 272760 244776
rect 272812 244764 272818 244776
rect 274870 244764 274876 244776
rect 272812 244736 274876 244764
rect 272812 244724 272818 244736
rect 274870 244724 274876 244736
rect 274928 244724 274934 244776
rect 321808 244764 321836 244804
rect 327862 244764 327868 244776
rect 321808 244736 327868 244764
rect 327862 244724 327868 244736
rect 327920 244724 327926 244776
rect 275882 244628 275888 244640
rect 271944 244600 275888 244628
rect 275882 244588 275888 244600
rect 275940 244588 275946 244640
rect 173118 243976 173124 244028
rect 173176 244016 173182 244028
rect 179006 244016 179012 244028
rect 173176 243988 179012 244016
rect 173176 243976 173182 243988
rect 179006 243976 179012 243988
rect 179064 243976 179070 244028
rect 321606 243432 321612 243484
rect 321664 243472 321670 243484
rect 327218 243472 327224 243484
rect 321664 243444 327224 243472
rect 321664 243432 321670 243444
rect 327218 243432 327224 243444
rect 327276 243432 327282 243484
rect 13130 243364 13136 243416
rect 13188 243404 13194 243416
rect 16166 243404 16172 243416
rect 13188 243376 16172 243404
rect 13188 243364 13194 243376
rect 16166 243364 16172 243376
rect 16224 243364 16230 243416
rect 173946 243364 173952 243416
rect 174004 243404 174010 243416
rect 181030 243404 181036 243416
rect 174004 243376 181036 243404
rect 174004 243364 174010 243376
rect 181030 243364 181036 243376
rect 181088 243364 181094 243416
rect 272846 243364 272852 243416
rect 272904 243404 272910 243416
rect 275422 243404 275428 243416
rect 272904 243376 275428 243404
rect 272904 243364 272910 243376
rect 275422 243364 275428 243376
rect 275480 243364 275486 243416
rect 323170 243364 323176 243416
rect 323228 243404 323234 243416
rect 327862 243404 327868 243416
rect 323228 243376 327868 243404
rect 323228 243364 323234 243376
rect 327862 243364 327868 243376
rect 327920 243364 327926 243416
rect 226478 243228 226484 243280
rect 226536 243268 226542 243280
rect 233470 243268 233476 243280
rect 226536 243240 233476 243268
rect 226536 243228 226542 243240
rect 233470 243228 233476 243240
rect 233528 243228 233534 243280
rect 132546 243160 132552 243212
rect 132604 243200 132610 243212
rect 137514 243200 137520 243212
rect 132604 243172 137520 243200
rect 132604 243160 132610 243172
rect 137514 243160 137520 243172
rect 137572 243160 137578 243212
rect 226478 243092 226484 243144
rect 226536 243132 226542 243144
rect 230066 243132 230072 243144
rect 226536 243104 230072 243132
rect 226536 243092 226542 243104
rect 230066 243092 230072 243104
rect 230124 243092 230130 243144
rect 78910 243024 78916 243076
rect 78968 243064 78974 243076
rect 87098 243064 87104 243076
rect 78968 243036 87104 243064
rect 78968 243024 78974 243036
rect 87098 243024 87104 243036
rect 87156 243024 87162 243076
rect 178914 242956 178920 243008
rect 178972 242996 178978 243008
rect 181214 242996 181220 243008
rect 178972 242968 181220 242996
rect 178972 242956 178978 242968
rect 181214 242956 181220 242968
rect 181272 242956 181278 243008
rect 225742 242888 225748 242940
rect 225800 242928 225806 242940
rect 230158 242928 230164 242940
rect 225800 242900 230164 242928
rect 225800 242888 225806 242900
rect 230158 242888 230164 242900
rect 230216 242888 230222 242940
rect 321606 242208 321612 242260
rect 321664 242248 321670 242260
rect 328046 242248 328052 242260
rect 321664 242220 328052 242248
rect 321664 242208 321670 242220
rect 328046 242208 328052 242220
rect 328104 242208 328110 242260
rect 79094 242140 79100 242192
rect 79152 242180 79158 242192
rect 87190 242180 87196 242192
rect 79152 242152 87196 242180
rect 79152 242140 79158 242152
rect 87190 242140 87196 242152
rect 87248 242140 87254 242192
rect 267878 242140 267884 242192
rect 267936 242180 267942 242192
rect 271466 242180 271472 242192
rect 267936 242152 271472 242180
rect 267936 242140 267942 242152
rect 271466 242140 271472 242152
rect 271524 242140 271530 242192
rect 79002 242072 79008 242124
rect 79060 242112 79066 242124
rect 87282 242112 87288 242124
rect 79060 242084 87288 242112
rect 79060 242072 79066 242084
rect 87282 242072 87288 242084
rect 87340 242072 87346 242124
rect 320502 242072 320508 242124
rect 320560 242112 320566 242124
rect 327862 242112 327868 242124
rect 320560 242084 327868 242112
rect 320560 242072 320566 242084
rect 327862 242072 327868 242084
rect 327920 242072 327926 242124
rect 123070 241596 123076 241648
rect 123128 241636 123134 241648
rect 124312 241636 124318 241648
rect 123128 241608 124318 241636
rect 123128 241596 123134 241608
rect 124312 241596 124318 241608
rect 124370 241596 124376 241648
rect 133374 240576 133380 240628
rect 133432 240616 133438 240628
rect 140550 240616 140556 240628
rect 133432 240588 140556 240616
rect 133432 240576 133438 240588
rect 140550 240576 140556 240588
rect 140608 240576 140614 240628
rect 173578 240576 173584 240628
rect 173636 240616 173642 240628
rect 181582 240616 181588 240628
rect 173636 240588 181588 240616
rect 173636 240576 173642 240588
rect 181582 240576 181588 240588
rect 181640 240576 181646 240628
rect 227214 240576 227220 240628
rect 227272 240616 227278 240628
rect 233470 240616 233476 240628
rect 227272 240588 233476 240616
rect 227272 240576 227278 240588
rect 233470 240576 233476 240588
rect 233528 240576 233534 240628
rect 267878 240576 267884 240628
rect 267936 240616 267942 240628
rect 275606 240616 275612 240628
rect 267936 240588 275612 240616
rect 267936 240576 267942 240588
rect 275606 240576 275612 240588
rect 275664 240576 275670 240628
rect 427406 240576 427412 240628
rect 427464 240616 427470 240628
rect 429522 240616 429528 240628
rect 427464 240588 429528 240616
rect 427464 240576 427470 240588
rect 429522 240576 429528 240588
rect 429580 240576 429586 240628
rect 358590 239964 358596 240016
rect 358648 240004 358654 240016
rect 389870 240004 389876 240016
rect 358648 239976 389876 240004
rect 358648 239964 358654 239976
rect 389870 239964 389876 239976
rect 389928 239964 389934 240016
rect 358498 239896 358504 239948
rect 358556 239936 358562 239948
rect 393826 239936 393832 239948
rect 358556 239908 393832 239936
rect 358556 239896 358562 239908
rect 393826 239896 393832 239908
rect 393884 239896 393890 239948
rect 314890 239828 314896 239880
rect 314948 239868 314954 239880
rect 316086 239868 316092 239880
rect 314948 239840 316092 239868
rect 314948 239828 314954 239840
rect 316086 239828 316092 239840
rect 316144 239828 316150 239880
rect 78910 239624 78916 239676
rect 78968 239664 78974 239676
rect 87006 239664 87012 239676
rect 78968 239636 87012 239664
rect 78968 239624 78974 239636
rect 87006 239624 87012 239636
rect 87064 239624 87070 239676
rect 364478 239352 364484 239404
rect 364536 239392 364542 239404
rect 377818 239392 377824 239404
rect 364536 239364 377824 239392
rect 364536 239352 364542 239364
rect 377818 239352 377824 239364
rect 377876 239352 377882 239404
rect 185630 239284 185636 239336
rect 185688 239324 185694 239336
rect 186458 239324 186464 239336
rect 185688 239296 186464 239324
rect 185688 239284 185694 239296
rect 186458 239284 186464 239296
rect 186516 239284 186522 239336
rect 279654 239284 279660 239336
rect 279712 239324 279718 239336
rect 280298 239324 280304 239336
rect 279712 239296 280304 239324
rect 279712 239284 279718 239296
rect 280298 239284 280304 239296
rect 280356 239284 280362 239336
rect 358317 239327 358375 239333
rect 358317 239293 358329 239327
rect 358363 239324 358375 239327
rect 381866 239324 381872 239336
rect 358363 239296 381872 239324
rect 358363 239293 358375 239296
rect 358317 239287 358375 239293
rect 381866 239284 381872 239296
rect 381924 239284 381930 239336
rect 132178 239216 132184 239268
rect 132236 239256 132242 239268
rect 140550 239256 140556 239268
rect 132236 239228 140556 239256
rect 132236 239216 132242 239228
rect 140550 239216 140556 239228
rect 140608 239216 140614 239268
rect 173394 239216 173400 239268
rect 173452 239256 173458 239268
rect 181950 239256 181956 239268
rect 173452 239228 181956 239256
rect 173452 239216 173458 239228
rect 181950 239216 181956 239228
rect 182008 239216 182014 239268
rect 226018 239216 226024 239268
rect 226076 239256 226082 239268
rect 233470 239256 233476 239268
rect 226076 239228 233476 239256
rect 226076 239216 226082 239228
rect 233470 239216 233476 239228
rect 233528 239216 233534 239268
rect 267602 239216 267608 239268
rect 267660 239256 267666 239268
rect 275698 239256 275704 239268
rect 267660 239228 275704 239256
rect 267660 239216 267666 239228
rect 275698 239216 275704 239228
rect 275756 239216 275762 239268
rect 266774 239148 266780 239200
rect 266832 239188 266838 239200
rect 275514 239188 275520 239200
rect 266832 239160 275520 239188
rect 266832 239148 266838 239160
rect 275514 239148 275520 239160
rect 275572 239148 275578 239200
rect 200166 238536 200172 238588
rect 200224 238576 200230 238588
rect 230894 238576 230900 238588
rect 200224 238548 230900 238576
rect 200224 238536 200230 238548
rect 230894 238536 230900 238548
rect 230952 238536 230958 238588
rect 290050 238536 290056 238588
rect 290108 238576 290114 238588
rect 290510 238576 290516 238588
rect 290108 238548 290516 238576
rect 290108 238536 290114 238548
rect 290510 238536 290516 238548
rect 290568 238576 290574 238588
rect 325194 238576 325200 238588
rect 290568 238548 325200 238576
rect 290568 238536 290574 238548
rect 325194 238536 325200 238548
rect 325252 238536 325258 238588
rect 221050 237788 221056 237840
rect 221108 237828 221114 237840
rect 222154 237828 222160 237840
rect 221108 237800 222160 237828
rect 221108 237788 221114 237800
rect 222154 237788 222160 237800
rect 222212 237788 222218 237840
rect 128130 237176 128136 237228
rect 128188 237216 128194 237228
rect 140366 237216 140372 237228
rect 128188 237188 140372 237216
rect 128188 237176 128194 237188
rect 140366 237176 140372 237188
rect 140424 237176 140430 237228
rect 172934 237176 172940 237228
rect 172992 237216 172998 237228
rect 219762 237216 219768 237228
rect 172992 237188 219768 237216
rect 172992 237176 172998 237188
rect 219762 237176 219768 237188
rect 219820 237216 219826 237228
rect 233470 237216 233476 237228
rect 219820 237188 233476 237216
rect 219820 237176 219826 237188
rect 233470 237176 233476 237188
rect 233528 237176 233534 237228
rect 267326 237176 267332 237228
rect 267384 237216 267390 237228
rect 316270 237216 316276 237228
rect 267384 237188 316276 237216
rect 267384 237176 267390 237188
rect 316270 237176 316276 237188
rect 316328 237176 316334 237228
rect 78910 236564 78916 236616
rect 78968 236604 78974 236616
rect 128130 236604 128136 236616
rect 78968 236576 128136 236604
rect 78968 236564 78974 236576
rect 128130 236564 128136 236576
rect 128188 236564 128194 236616
rect 316270 236564 316276 236616
rect 316328 236604 316334 236616
rect 328414 236604 328420 236616
rect 316328 236576 328420 236604
rect 316328 236564 316334 236576
rect 328414 236564 328420 236576
rect 328472 236564 328478 236616
rect 296950 236332 296956 236344
rect 262652 236304 296956 236332
rect 262652 236208 262680 236304
rect 296950 236292 296956 236304
rect 297008 236332 297014 236344
rect 298238 236332 298244 236344
rect 297008 236304 298244 236332
rect 297008 236292 297014 236304
rect 298238 236292 298244 236304
rect 298296 236292 298302 236344
rect 262634 236156 262640 236208
rect 262692 236156 262698 236208
rect 298238 235884 298244 235936
rect 298296 235924 298302 235936
rect 324826 235924 324832 235936
rect 298296 235896 324832 235924
rect 298296 235884 298302 235896
rect 324826 235884 324832 235896
rect 324884 235884 324890 235936
rect 203110 235816 203116 235868
rect 203168 235856 203174 235868
rect 230986 235856 230992 235868
rect 203168 235828 230992 235856
rect 203168 235816 203174 235828
rect 230986 235816 230992 235828
rect 231044 235816 231050 235868
rect 286922 235816 286928 235868
rect 286980 235856 286986 235868
rect 325378 235856 325384 235868
rect 286980 235828 325384 235856
rect 286980 235816 286986 235828
rect 325378 235816 325384 235828
rect 325436 235816 325442 235868
rect 145334 235612 145340 235664
rect 145392 235652 145398 235664
rect 146208 235652 146214 235664
rect 145392 235624 146214 235652
rect 145392 235612 145398 235624
rect 146208 235612 146214 235624
rect 146266 235612 146272 235664
rect 136870 235272 136876 235324
rect 136928 235312 136934 235324
rect 137238 235312 137244 235324
rect 136928 235284 137244 235312
rect 136928 235272 136934 235284
rect 137238 235272 137244 235284
rect 137296 235312 137302 235324
rect 145150 235312 145156 235324
rect 137296 235284 145156 235312
rect 137296 235272 137302 235284
rect 145150 235272 145156 235284
rect 145208 235312 145214 235324
rect 152602 235312 152608 235324
rect 145208 235284 152608 235312
rect 145208 235272 145214 235284
rect 152602 235272 152608 235284
rect 152660 235272 152666 235324
rect 137054 235204 137060 235256
rect 137112 235244 137118 235256
rect 150394 235244 150400 235256
rect 137112 235216 150400 235244
rect 137112 235204 137118 235216
rect 150394 235204 150400 235216
rect 150452 235244 150458 235256
rect 167690 235244 167696 235256
rect 150452 235216 167696 235244
rect 150452 235204 150458 235216
rect 167690 235204 167696 235216
rect 167748 235204 167754 235256
rect 149106 235136 149112 235188
rect 149164 235176 149170 235188
rect 167966 235176 167972 235188
rect 149164 235148 167972 235176
rect 149164 235136 149170 235148
rect 167966 235136 167972 235148
rect 168024 235136 168030 235188
rect 230986 235136 230992 235188
rect 231044 235176 231050 235188
rect 244970 235176 244976 235188
rect 231044 235148 244976 235176
rect 231044 235136 231050 235148
rect 244970 235136 244976 235148
rect 245028 235176 245034 235188
rect 262542 235176 262548 235188
rect 245028 235148 262548 235176
rect 245028 235136 245034 235148
rect 262542 235136 262548 235148
rect 262600 235136 262606 235188
rect 76058 235068 76064 235120
rect 76116 235108 76122 235120
rect 113502 235108 113508 235120
rect 76116 235080 113508 235108
rect 76116 235068 76122 235080
rect 113502 235068 113508 235080
rect 113560 235108 113566 235120
rect 113870 235108 113876 235120
rect 113560 235080 113876 235108
rect 113560 235068 113566 235080
rect 113870 235068 113876 235080
rect 113928 235068 113934 235120
rect 359694 235068 359700 235120
rect 359752 235108 359758 235120
rect 368710 235108 368716 235120
rect 359752 235080 368716 235108
rect 359752 235068 359758 235080
rect 368710 235068 368716 235080
rect 368768 235068 368774 235120
rect 113870 234388 113876 234440
rect 113928 234428 113934 234440
rect 137330 234428 137336 234440
rect 113928 234400 137336 234428
rect 113928 234388 113934 234400
rect 137330 234388 137336 234400
rect 137388 234388 137394 234440
rect 301090 234388 301096 234440
rect 301148 234428 301154 234440
rect 324918 234428 324924 234440
rect 301148 234400 324924 234428
rect 301148 234388 301154 234400
rect 324918 234388 324924 234400
rect 324976 234388 324982 234440
rect 346538 234388 346544 234440
rect 346596 234428 346602 234440
rect 360614 234428 360620 234440
rect 346596 234400 360620 234428
rect 346596 234388 346602 234400
rect 360614 234388 360620 234400
rect 360672 234388 360678 234440
rect 324918 233776 324924 233828
rect 324976 233816 324982 233828
rect 345250 233816 345256 233828
rect 324976 233788 345256 233816
rect 324976 233776 324982 233788
rect 345250 233776 345256 233788
rect 345308 233816 345314 233828
rect 346538 233816 346544 233828
rect 345308 233788 346544 233816
rect 345308 233776 345314 233788
rect 346538 233776 346544 233788
rect 346596 233776 346602 233828
rect 63638 233708 63644 233760
rect 63696 233748 63702 233760
rect 63696 233720 69940 233748
rect 63696 233708 63702 233720
rect 61798 233572 61804 233624
rect 61856 233612 61862 233624
rect 65754 233612 65760 233624
rect 61856 233584 65760 233612
rect 61856 233572 61862 233584
rect 65754 233572 65760 233584
rect 65812 233572 65818 233624
rect 62810 233504 62816 233556
rect 62868 233544 62874 233556
rect 65846 233544 65852 233556
rect 62868 233516 65852 233544
rect 62868 233504 62874 233516
rect 65846 233504 65852 233516
rect 65904 233504 65910 233556
rect 69912 233544 69940 233720
rect 138158 233708 138164 233760
rect 138216 233748 138222 233760
rect 146806 233748 146812 233760
rect 138216 233720 146812 233748
rect 138216 233708 138222 233720
rect 146806 233708 146812 233720
rect 146864 233708 146870 233760
rect 149290 233708 149296 233760
rect 149348 233748 149354 233760
rect 162262 233748 162268 233760
rect 149348 233720 162268 233748
rect 149348 233708 149354 233720
rect 162262 233708 162268 233720
rect 162320 233708 162326 233760
rect 234758 233708 234764 233760
rect 234816 233748 234822 233760
rect 241474 233748 241480 233760
rect 234816 233720 241480 233748
rect 234816 233708 234822 233720
rect 241474 233708 241480 233720
rect 241532 233708 241538 233760
rect 246258 233708 246264 233760
rect 246316 233748 246322 233760
rect 259230 233748 259236 233760
rect 246316 233720 259236 233748
rect 246316 233708 246322 233720
rect 259230 233708 259236 233720
rect 259288 233708 259294 233760
rect 323814 233708 323820 233760
rect 323872 233748 323878 233760
rect 368710 233748 368716 233760
rect 323872 233720 368716 233748
rect 323872 233708 323878 233720
rect 368710 233708 368716 233720
rect 368768 233708 368774 233760
rect 154718 233640 154724 233692
rect 154776 233680 154782 233692
rect 168058 233680 168064 233692
rect 154776 233652 168064 233680
rect 154776 233640 154782 233652
rect 168058 233640 168064 233652
rect 168116 233640 168122 233692
rect 248926 233640 248932 233692
rect 248984 233680 248990 233692
rect 262082 233680 262088 233692
rect 248984 233652 262088 233680
rect 248984 233640 248990 233652
rect 262082 233640 262088 233652
rect 262140 233640 262146 233692
rect 243590 233572 243596 233624
rect 243648 233612 243654 233624
rect 256286 233612 256292 233624
rect 243648 233584 256292 233612
rect 243648 233572 243654 233584
rect 256286 233572 256292 233584
rect 256344 233572 256350 233624
rect 362454 233572 362460 233624
rect 362512 233612 362518 233624
rect 368802 233612 368808 233624
rect 362512 233584 368808 233612
rect 362512 233572 362518 233584
rect 368802 233572 368808 233584
rect 368860 233572 368866 233624
rect 75230 233544 75236 233556
rect 69912 233516 75236 233544
rect 75230 233504 75236 233516
rect 75288 233504 75294 233556
rect 153338 233504 153344 233556
rect 153396 233544 153402 233556
rect 166126 233544 166132 233556
rect 153396 233516 166132 233544
rect 153396 233504 153402 233516
rect 166126 233504 166132 233516
rect 166184 233504 166190 233556
rect 248006 233504 248012 233556
rect 248064 233544 248070 233556
rect 261162 233544 261168 233556
rect 248064 233516 261168 233544
rect 248064 233504 248070 233516
rect 261162 233504 261168 233516
rect 261220 233504 261226 233556
rect 340926 233504 340932 233556
rect 340984 233544 340990 233556
rect 347918 233544 347924 233556
rect 340984 233516 347924 233544
rect 340984 233504 340990 233516
rect 347918 233504 347924 233516
rect 347976 233504 347982 233556
rect 64834 233436 64840 233488
rect 64892 233476 64898 233488
rect 67134 233476 67140 233488
rect 64892 233448 67140 233476
rect 64892 233436 64898 233448
rect 67134 233436 67140 233448
rect 67192 233436 67198 233488
rect 249938 233436 249944 233488
rect 249996 233476 250002 233488
rect 263094 233476 263100 233488
rect 249996 233448 263100 233476
rect 249996 233436 250002 233448
rect 263094 233436 263100 233448
rect 263152 233436 263158 233488
rect 63822 233368 63828 233420
rect 63880 233408 63886 233420
rect 67226 233408 67232 233420
rect 63880 233380 67232 233408
rect 63880 233368 63886 233380
rect 67226 233368 67232 233380
rect 67284 233368 67290 233420
rect 151958 233368 151964 233420
rect 152016 233408 152022 233420
rect 165206 233408 165212 233420
rect 152016 233380 165212 233408
rect 152016 233368 152022 233380
rect 165206 233368 165212 233380
rect 165264 233368 165270 233420
rect 340834 233368 340840 233420
rect 340892 233408 340898 233420
rect 346814 233408 346820 233420
rect 340892 233380 346820 233408
rect 340892 233368 340898 233380
rect 346814 233368 346820 233380
rect 346872 233368 346878 233420
rect 365214 233368 365220 233420
rect 365272 233408 365278 233420
rect 368710 233408 368716 233420
rect 365272 233380 368716 233408
rect 365272 233368 365278 233380
rect 368710 233368 368716 233380
rect 368768 233368 368774 233420
rect 58118 233300 58124 233352
rect 58176 233340 58182 233352
rect 70078 233340 70084 233352
rect 58176 233312 70084 233340
rect 58176 233300 58182 233312
rect 70078 233300 70084 233312
rect 70136 233300 70142 233352
rect 231446 233300 231452 233352
rect 231504 233340 231510 233352
rect 234758 233340 234764 233352
rect 231504 233312 234764 233340
rect 231504 233300 231510 233312
rect 234758 233300 234764 233312
rect 234816 233300 234822 233352
rect 250674 233300 250680 233352
rect 250732 233340 250738 233352
rect 264014 233340 264020 233352
rect 250732 233312 264020 233340
rect 250732 233300 250738 233312
rect 264014 233300 264020 233312
rect 264072 233300 264078 233352
rect 56738 233232 56744 233284
rect 56796 233272 56802 233284
rect 67962 233272 67968 233284
rect 56796 233244 67968 233272
rect 56796 233232 56802 233244
rect 67962 233232 67968 233244
rect 68020 233232 68026 233284
rect 153706 233232 153712 233284
rect 153764 233272 153770 233284
rect 167322 233272 167328 233284
rect 153764 233244 167328 233272
rect 153764 233232 153770 233244
rect 167322 233232 167328 233244
rect 167380 233232 167386 233284
rect 231722 233232 231728 233284
rect 231780 233272 231786 233284
rect 243038 233272 243044 233284
rect 231780 233244 243044 233272
rect 231780 233232 231786 233244
rect 243038 233232 243044 233244
rect 243096 233232 243102 233284
rect 245338 233232 245344 233284
rect 245396 233272 245402 233284
rect 258402 233272 258408 233284
rect 245396 233244 258408 233272
rect 245396 233232 245402 233244
rect 258402 233232 258408 233244
rect 258460 233232 258466 233284
rect 62258 233164 62264 233216
rect 62316 233204 62322 233216
rect 74218 233204 74224 233216
rect 62316 233176 74224 233204
rect 62316 233164 62322 233176
rect 74218 233164 74224 233176
rect 74276 233164 74282 233216
rect 96761 233207 96819 233213
rect 96761 233173 96773 233207
rect 96807 233204 96819 233207
rect 150670 233204 150676 233216
rect 96807 233176 96896 233204
rect 96807 233173 96819 233176
rect 96761 233167 96819 233173
rect 55358 233096 55364 233148
rect 55416 233136 55422 233148
rect 66950 233136 66956 233148
rect 55416 233108 66956 233136
rect 55416 233096 55422 233108
rect 66950 233096 66956 233108
rect 67008 233096 67014 233148
rect 74126 233096 74132 233148
rect 74184 233136 74190 233148
rect 96868 233145 96896 233176
rect 138176 233176 150676 233204
rect 77533 233139 77591 233145
rect 77533 233136 77545 233139
rect 74184 233108 77545 233136
rect 74184 233096 74190 233108
rect 77533 233105 77545 233108
rect 77579 233105 77591 233139
rect 95381 233139 95439 233145
rect 95381 233136 95393 233139
rect 77533 233099 77591 233105
rect 87024 233108 95393 233136
rect 60786 233028 60792 233080
rect 60844 233068 60850 233080
rect 73114 233068 73120 233080
rect 60844 233040 73120 233068
rect 60844 233028 60850 233040
rect 73114 233028 73120 233040
rect 73172 233028 73178 233080
rect 77533 233003 77591 233009
rect 77533 232969 77545 233003
rect 77579 233000 77591 233003
rect 87024 233000 87052 233108
rect 95381 233105 95393 233108
rect 95427 233105 95439 233139
rect 95381 233099 95439 233105
rect 96853 233139 96911 233145
rect 96853 233105 96865 233139
rect 96899 233105 96911 233139
rect 96853 233099 96911 233105
rect 101637 233139 101695 233145
rect 101637 233105 101649 233139
rect 101683 233136 101695 233139
rect 105133 233139 105191 233145
rect 105133 233136 105145 233139
rect 101683 233108 105145 233136
rect 101683 233105 101695 233108
rect 101637 233099 101695 233105
rect 105133 233105 105145 233108
rect 105179 233105 105191 233139
rect 137146 233136 137152 233148
rect 105133 233099 105191 233105
rect 128608 233108 137152 233136
rect 77579 232972 87052 233000
rect 95381 233003 95439 233009
rect 77579 232969 77591 232972
rect 77533 232963 77591 232969
rect 95381 232969 95393 233003
rect 95427 233000 95439 233003
rect 96761 233003 96819 233009
rect 96761 233000 96773 233003
rect 95427 232972 96773 233000
rect 95427 232969 95439 232972
rect 95381 232963 95439 232969
rect 96761 232969 96773 232972
rect 96807 232969 96819 233003
rect 96761 232963 96819 232969
rect 96853 233003 96911 233009
rect 96853 232969 96865 233003
rect 96899 233000 96911 233003
rect 101637 233003 101695 233009
rect 101637 233000 101649 233003
rect 96899 232972 101649 233000
rect 96899 232969 96911 232972
rect 96853 232963 96911 232969
rect 101637 232969 101649 232972
rect 101683 232969 101695 233003
rect 101637 232963 101695 232969
rect 120957 233003 121015 233009
rect 120957 232969 120969 233003
rect 121003 233000 121015 233003
rect 128608 233000 128636 233108
rect 137146 233096 137152 233108
rect 137204 233136 137210 233148
rect 138176 233136 138204 233176
rect 150670 233164 150676 233176
rect 150728 233164 150734 233216
rect 151038 233164 151044 233216
rect 151096 233204 151102 233216
rect 164562 233204 164568 233216
rect 151096 233176 164568 233204
rect 151096 233164 151102 233176
rect 164562 233164 164568 233176
rect 164620 233164 164626 233216
rect 231630 233164 231636 233216
rect 231688 233204 231694 233216
rect 242118 233204 242124 233216
rect 231688 233176 242124 233204
rect 231688 233164 231694 233176
rect 242118 233164 242124 233176
rect 242176 233164 242182 233216
rect 244326 233164 244332 233216
rect 244384 233204 244390 233216
rect 257298 233204 257304 233216
rect 244384 233176 257304 233204
rect 244384 233164 244390 233176
rect 257298 233164 257304 233176
rect 257356 233164 257362 233216
rect 137204 233108 138204 233136
rect 137204 233096 137210 233108
rect 144598 233096 144604 233148
rect 144656 233136 144662 233148
rect 165114 233136 165120 233148
rect 144656 233108 165120 233136
rect 144656 233096 144662 233108
rect 165114 233096 165120 233108
rect 165172 233096 165178 233148
rect 238622 233096 238628 233148
rect 238680 233136 238686 233148
rect 250125 233139 250183 233145
rect 238680 233108 240278 233136
rect 238680 233096 238686 233108
rect 145242 233028 145248 233080
rect 145300 233068 145306 233080
rect 222433 233071 222491 233077
rect 222433 233068 222445 233071
rect 145300 233040 222445 233068
rect 145300 233028 145306 233040
rect 222433 233037 222445 233040
rect 222479 233037 222491 233071
rect 222433 233031 222491 233037
rect 121003 232972 128636 233000
rect 121003 232969 121015 232972
rect 120957 232963 121015 232969
rect 156374 232960 156380 233012
rect 156432 233000 156438 233012
rect 169990 233000 169996 233012
rect 156432 232972 169996 233000
rect 156432 232960 156438 232972
rect 169990 232960 169996 232972
rect 170048 232960 170054 233012
rect 222525 233003 222583 233009
rect 222525 232969 222537 233003
rect 222571 233000 222583 233003
rect 222571 232972 240140 233000
rect 222571 232969 222583 232972
rect 222525 232963 222583 232969
rect 59498 232892 59504 232944
rect 59556 232932 59562 232944
rect 71090 232932 71096 232944
rect 59556 232904 71096 232932
rect 59556 232892 59562 232904
rect 71090 232892 71096 232904
rect 71148 232892 71154 232944
rect 114701 232935 114759 232941
rect 114701 232901 114713 232935
rect 114747 232932 114759 232935
rect 116173 232935 116231 232941
rect 116173 232932 116185 232935
rect 114747 232904 116185 232932
rect 114747 232901 114759 232904
rect 114701 232895 114759 232901
rect 116173 232901 116185 232904
rect 116219 232901 116231 232935
rect 116173 232895 116231 232901
rect 155454 232892 155460 232944
rect 155512 232932 155518 232944
rect 169070 232932 169076 232944
rect 155512 232904 169076 232932
rect 155512 232892 155518 232904
rect 169070 232892 169076 232904
rect 169128 232892 169134 232944
rect 60878 232824 60884 232876
rect 60936 232864 60942 232876
rect 72102 232864 72108 232876
rect 60936 232836 72108 232864
rect 60936 232824 60942 232836
rect 72102 232824 72108 232836
rect 72160 232824 72166 232876
rect 150578 232824 150584 232876
rect 150636 232864 150642 232876
rect 163274 232864 163280 232876
rect 150636 232836 163280 232864
rect 150636 232824 150642 232836
rect 163274 232824 163280 232836
rect 163332 232824 163338 232876
rect 105133 232799 105191 232805
rect 105133 232765 105145 232799
rect 105179 232796 105191 232799
rect 109270 232796 109276 232808
rect 105179 232768 109276 232796
rect 105179 232765 105191 232768
rect 105133 232759 105191 232765
rect 109270 232756 109276 232768
rect 109328 232796 109334 232808
rect 114701 232799 114759 232805
rect 114701 232796 114713 232799
rect 109328 232768 114713 232796
rect 109328 232756 109334 232768
rect 114701 232765 114713 232768
rect 114747 232765 114759 232799
rect 114701 232759 114759 232765
rect 116173 232799 116231 232805
rect 116173 232765 116185 232799
rect 116219 232796 116231 232799
rect 120957 232799 121015 232805
rect 120957 232796 120969 232799
rect 116219 232768 120969 232796
rect 116219 232765 116231 232768
rect 116173 232759 116231 232765
rect 120957 232765 120969 232768
rect 121003 232765 121015 232799
rect 240112 232796 240140 232972
rect 240250 232864 240278 233108
rect 250125 233105 250137 233139
rect 250171 233136 250183 233139
rect 250171 233108 254308 233136
rect 250171 233105 250183 233108
rect 250125 233099 250183 233105
rect 250033 233071 250091 233077
rect 250033 233037 250045 233071
rect 250079 233037 250091 233071
rect 254280 233068 254308 233108
rect 352886 233068 352892 233080
rect 254280 233040 352892 233068
rect 250033 233031 250091 233037
rect 244513 233003 244571 233009
rect 244513 232969 244525 233003
rect 244559 233000 244571 233003
rect 250048 233000 250076 233031
rect 352886 233028 352892 233040
rect 352944 233028 352950 233080
rect 244559 232972 250076 233000
rect 244559 232969 244571 232972
rect 244513 232963 244571 232969
rect 247086 232892 247092 232944
rect 247144 232932 247150 232944
rect 260150 232932 260156 232944
rect 247144 232904 260156 232932
rect 247144 232892 247150 232904
rect 260150 232892 260156 232904
rect 260208 232892 260214 232944
rect 258954 232864 258960 232876
rect 240250 232836 258960 232864
rect 258954 232824 258960 232836
rect 259012 232824 259018 232876
rect 244513 232799 244571 232805
rect 244513 232796 244525 232799
rect 240112 232768 244525 232796
rect 120957 232759 121015 232765
rect 244513 232765 244525 232768
rect 244559 232765 244571 232799
rect 244513 232759 244571 232765
rect 158858 232688 158864 232740
rect 158916 232728 158922 232740
rect 161802 232728 161808 232740
rect 158916 232700 161808 232728
rect 158916 232688 158922 232700
rect 161802 232688 161808 232700
rect 161860 232688 161866 232740
rect 58670 232620 58676 232672
rect 58728 232660 58734 232672
rect 63086 232660 63092 232672
rect 58728 232632 63092 232660
rect 58728 232620 58734 232632
rect 63086 232620 63092 232632
rect 63144 232620 63150 232672
rect 156098 232620 156104 232672
rect 156156 232660 156162 232672
rect 158030 232660 158036 232672
rect 156156 232632 158036 232660
rect 156156 232620 156162 232632
rect 158030 232620 158036 232632
rect 158088 232620 158094 232672
rect 158122 232620 158128 232672
rect 158180 232660 158186 232672
rect 160330 232660 160336 232672
rect 158180 232632 160336 232660
rect 158180 232620 158186 232632
rect 160330 232620 160336 232632
rect 160388 232620 160394 232672
rect 256010 232620 256016 232672
rect 256068 232660 256074 232672
rect 258310 232660 258316 232672
rect 256068 232632 258316 232660
rect 256068 232620 256074 232632
rect 258310 232620 258316 232632
rect 258368 232620 258374 232672
rect 59682 232552 59688 232604
rect 59740 232592 59746 232604
rect 63178 232592 63184 232604
rect 59740 232564 63184 232592
rect 59740 232552 59746 232564
rect 63178 232552 63184 232564
rect 63236 232552 63242 232604
rect 155178 232552 155184 232604
rect 155236 232592 155242 232604
rect 157570 232592 157576 232604
rect 155236 232564 157576 232592
rect 155236 232552 155242 232564
rect 157570 232552 157576 232564
rect 157628 232552 157634 232604
rect 252698 232552 252704 232604
rect 252756 232592 252762 232604
rect 255550 232592 255556 232604
rect 252756 232564 255556 232592
rect 252756 232552 252762 232564
rect 255550 232552 255556 232564
rect 255608 232552 255614 232604
rect 57658 232484 57664 232536
rect 57716 232524 57722 232536
rect 61614 232524 61620 232536
rect 57716 232496 61620 232524
rect 57716 232484 57722 232496
rect 61614 232484 61620 232496
rect 61672 232484 61678 232536
rect 65938 232484 65944 232536
rect 65996 232524 66002 232536
rect 68514 232524 68520 232536
rect 65996 232496 68520 232524
rect 65996 232484 66002 232496
rect 68514 232484 68520 232496
rect 68572 232484 68578 232536
rect 157110 232484 157116 232536
rect 157168 232524 157174 232536
rect 159134 232524 159140 232536
rect 157168 232496 159140 232524
rect 157168 232484 157174 232496
rect 159134 232484 159140 232496
rect 159192 232484 159198 232536
rect 160054 232484 160060 232536
rect 160112 232524 160118 232536
rect 162262 232524 162268 232536
rect 160112 232496 162268 232524
rect 160112 232484 160118 232496
rect 162262 232484 162268 232496
rect 162320 232484 162326 232536
rect 254078 232484 254084 232536
rect 254136 232524 254142 232536
rect 255642 232524 255648 232536
rect 254136 232496 255648 232524
rect 254136 232484 254142 232496
rect 255642 232484 255648 232496
rect 255700 232484 255706 232536
rect 60694 232416 60700 232468
rect 60752 232456 60758 232468
rect 62994 232456 63000 232468
rect 60752 232428 63000 232456
rect 60752 232416 60758 232428
rect 62994 232416 63000 232428
rect 63052 232416 63058 232468
rect 67318 232416 67324 232468
rect 67376 232456 67382 232468
rect 68974 232456 68980 232468
rect 67376 232428 68980 232456
rect 67376 232416 67382 232428
rect 68974 232416 68980 232428
rect 69032 232416 69038 232468
rect 154258 232416 154264 232468
rect 154316 232456 154322 232468
rect 156742 232456 156748 232468
rect 154316 232428 156748 232456
rect 154316 232416 154322 232428
rect 156742 232416 156748 232428
rect 156800 232416 156806 232468
rect 160974 232416 160980 232468
rect 161032 232456 161038 232468
rect 163182 232456 163188 232468
rect 161032 232428 163188 232456
rect 161032 232416 161038 232428
rect 163182 232416 163188 232428
rect 163240 232416 163246 232468
rect 248282 232416 248288 232468
rect 248340 232456 248346 232468
rect 250766 232456 250772 232468
rect 248340 232428 250772 232456
rect 248340 232416 248346 232428
rect 250766 232416 250772 232428
rect 250824 232416 250830 232468
rect 252146 232416 252152 232468
rect 252204 232456 252210 232468
rect 254170 232456 254176 232468
rect 252204 232428 254176 232456
rect 252204 232416 252210 232428
rect 254170 232416 254176 232428
rect 254228 232416 254234 232468
rect 254998 232416 255004 232468
rect 255056 232456 255062 232468
rect 256930 232456 256936 232468
rect 255056 232428 256936 232456
rect 255056 232416 255062 232428
rect 256930 232416 256936 232428
rect 256988 232416 256994 232468
rect 333382 232416 333388 232468
rect 333440 232456 333446 232468
rect 334118 232456 334124 232468
rect 333440 232428 334124 232456
rect 333440 232416 333446 232428
rect 334118 232416 334124 232428
rect 334176 232416 334182 232468
rect 334394 232416 334400 232468
rect 334452 232456 334458 232468
rect 335406 232456 335412 232468
rect 334452 232428 335412 232456
rect 334452 232416 334458 232428
rect 335406 232416 335412 232428
rect 335464 232416 335470 232468
rect 338534 232416 338540 232468
rect 338592 232456 338598 232468
rect 339638 232456 339644 232468
rect 338592 232428 339644 232456
rect 338592 232416 338598 232428
rect 339638 232416 339644 232428
rect 339696 232416 339702 232468
rect 342674 232416 342680 232468
rect 342732 232456 342738 232468
rect 344790 232456 344796 232468
rect 342732 232428 344796 232456
rect 342732 232416 342738 232428
rect 344790 232416 344796 232428
rect 344848 232416 344854 232468
rect 348102 232416 348108 232468
rect 348160 232456 348166 232468
rect 349942 232456 349948 232468
rect 348160 232428 349948 232456
rect 348160 232416 348166 232428
rect 349942 232416 349948 232428
rect 350000 232416 350006 232468
rect 134846 232348 134852 232400
rect 134904 232388 134910 232400
rect 368894 232388 368900 232400
rect 134904 232360 368900 232388
rect 134904 232348 134910 232360
rect 368894 232348 368900 232360
rect 368952 232348 368958 232400
rect 229974 232280 229980 232332
rect 230032 232320 230038 232332
rect 368710 232320 368716 232332
rect 230032 232292 368716 232320
rect 230032 232280 230038 232292
rect 368710 232280 368716 232292
rect 368768 232280 368774 232332
rect 326574 232212 326580 232264
rect 326632 232252 326638 232264
rect 368802 232252 368808 232264
rect 326632 232224 368808 232252
rect 326632 232212 326638 232224
rect 368802 232212 368808 232224
rect 368860 232212 368866 232264
rect 345710 231668 345716 231720
rect 345768 231708 345774 231720
rect 360522 231708 360528 231720
rect 345768 231680 360528 231708
rect 345768 231668 345774 231680
rect 360522 231668 360528 231680
rect 360580 231668 360586 231720
rect 222614 230988 222620 231040
rect 222672 231028 222678 231040
rect 222798 231028 222804 231040
rect 222672 231000 222804 231028
rect 222672 230988 222678 231000
rect 222798 230988 222804 231000
rect 222856 230988 222862 231040
rect 324826 230988 324832 231040
rect 324884 231028 324890 231040
rect 325746 231028 325752 231040
rect 324884 231000 325752 231028
rect 324884 230988 324890 231000
rect 325746 230988 325752 231000
rect 325804 231028 325810 231040
rect 345434 231028 345440 231040
rect 325804 231000 345440 231028
rect 325804 230988 325810 231000
rect 345434 230988 345440 231000
rect 345492 231028 345498 231040
rect 345710 231028 345716 231040
rect 345492 231000 345716 231028
rect 345492 230988 345498 231000
rect 345710 230988 345716 231000
rect 345768 230988 345774 231040
rect 358314 231028 358320 231040
rect 358275 231000 358320 231028
rect 358314 230988 358320 231000
rect 358372 230988 358378 231040
rect 47078 230920 47084 230972
rect 47136 230960 47142 230972
rect 368894 230960 368900 230972
rect 47136 230932 368900 230960
rect 47136 230920 47142 230932
rect 368894 230920 368900 230932
rect 368952 230920 368958 230972
rect 76794 230852 76800 230904
rect 76852 230892 76858 230904
rect 368710 230892 368716 230904
rect 76852 230864 368716 230892
rect 76852 230852 76858 230864
rect 368710 230852 368716 230864
rect 368768 230852 368774 230904
rect 134754 230784 134760 230836
rect 134812 230824 134818 230836
rect 368802 230824 368808 230836
rect 134812 230796 368808 230824
rect 134812 230784 134818 230796
rect 368802 230784 368808 230796
rect 368860 230784 368866 230836
rect 115986 230376 115992 230428
rect 116044 230416 116050 230428
rect 127210 230416 127216 230428
rect 116044 230388 127216 230416
rect 116044 230376 116050 230388
rect 127210 230376 127216 230388
rect 127268 230376 127274 230428
rect 210010 230376 210016 230428
rect 210068 230416 210074 230428
rect 221050 230416 221056 230428
rect 210068 230388 221056 230416
rect 210068 230376 210074 230388
rect 221050 230376 221056 230388
rect 221108 230376 221114 230428
rect 304034 230376 304040 230428
rect 304092 230416 304098 230428
rect 314890 230416 314896 230428
rect 304092 230388 314896 230416
rect 304092 230376 304098 230388
rect 314890 230376 314896 230388
rect 314948 230376 314954 230428
rect 103474 230308 103480 230360
rect 103532 230348 103538 230360
rect 123070 230348 123076 230360
rect 103532 230320 123076 230348
rect 103532 230308 103538 230320
rect 123070 230308 123076 230320
rect 123128 230308 123134 230360
rect 197498 230308 197504 230360
rect 197556 230348 197562 230360
rect 218290 230348 218296 230360
rect 197556 230320 218296 230348
rect 197556 230308 197562 230320
rect 218290 230308 218296 230320
rect 218348 230308 218354 230360
rect 291522 230308 291528 230360
rect 291580 230348 291586 230360
rect 312130 230348 312136 230360
rect 291580 230320 312136 230348
rect 291580 230308 291586 230320
rect 312130 230308 312136 230320
rect 312188 230308 312194 230360
rect 91054 230240 91060 230292
rect 91112 230280 91118 230292
rect 120310 230280 120316 230292
rect 91112 230252 120316 230280
rect 91112 230240 91118 230252
rect 120310 230240 120316 230252
rect 120368 230240 120374 230292
rect 185078 230240 185084 230292
rect 185136 230280 185142 230292
rect 214150 230280 214156 230292
rect 185136 230252 214156 230280
rect 185136 230240 185142 230252
rect 214150 230240 214156 230252
rect 214208 230240 214214 230292
rect 279102 230240 279108 230292
rect 279160 230280 279166 230292
rect 307990 230280 307996 230292
rect 279160 230252 307996 230280
rect 279160 230240 279166 230252
rect 307990 230240 307996 230252
rect 308048 230240 308054 230292
rect 343778 230240 343784 230292
rect 343836 230280 343842 230292
rect 360890 230280 360896 230292
rect 343836 230252 360896 230280
rect 343836 230240 343842 230252
rect 360890 230240 360896 230252
rect 360948 230240 360954 230292
rect 324642 229628 324648 229680
rect 324700 229668 324706 229680
rect 325470 229668 325476 229680
rect 324700 229640 325476 229668
rect 324700 229628 324706 229640
rect 325470 229628 325476 229640
rect 325528 229668 325534 229680
rect 343226 229668 343232 229680
rect 325528 229640 343232 229668
rect 325528 229628 325534 229640
rect 343226 229628 343232 229640
rect 343284 229668 343290 229680
rect 343778 229668 343784 229680
rect 343284 229640 343784 229668
rect 343284 229628 343290 229640
rect 343778 229628 343784 229640
rect 343836 229628 343842 229680
rect 13038 229560 13044 229612
rect 13096 229600 13102 229612
rect 16074 229600 16080 229612
rect 13096 229572 16080 229600
rect 13096 229560 13102 229572
rect 16074 229560 16080 229572
rect 16132 229560 16138 229612
rect 22238 229560 22244 229612
rect 22296 229600 22302 229612
rect 368710 229600 368716 229612
rect 22296 229572 368716 229600
rect 22296 229560 22302 229572
rect 368710 229560 368716 229572
rect 368768 229560 368774 229612
rect 369909 229059 369967 229065
rect 369909 229025 369921 229059
rect 369955 229056 369967 229059
rect 369998 229056 370004 229068
rect 369955 229028 370004 229056
rect 369955 229025 369967 229028
rect 369909 229019 369967 229025
rect 369998 229016 370004 229028
rect 370056 229016 370062 229068
rect 345250 228880 345256 228932
rect 345308 228920 345314 228932
rect 346078 228920 346084 228932
rect 345308 228892 346084 228920
rect 345308 228880 345314 228892
rect 346078 228880 346084 228892
rect 346136 228880 346142 228932
rect 354910 228880 354916 228932
rect 354968 228920 354974 228932
rect 355830 228920 355836 228932
rect 354968 228892 355836 228920
rect 354968 228880 354974 228892
rect 355830 228880 355836 228892
rect 355888 228880 355894 228932
rect 369814 228880 369820 228932
rect 369872 228920 369878 228932
rect 369998 228920 370004 228932
rect 369872 228892 370004 228920
rect 369872 228880 369878 228892
rect 369998 228880 370004 228892
rect 370056 228880 370062 228932
rect 74034 228404 74040 228456
rect 74092 228444 74098 228456
rect 368710 228444 368716 228456
rect 74092 228416 368716 228444
rect 74092 228404 74098 228416
rect 368710 228404 368716 228416
rect 368768 228404 368774 228456
rect 47078 228336 47084 228388
rect 47136 228376 47142 228388
rect 368802 228376 368808 228388
rect 47136 228348 368808 228376
rect 47136 228336 47142 228348
rect 368802 228336 368808 228348
rect 368860 228336 368866 228388
rect 34014 228268 34020 228320
rect 34072 228308 34078 228320
rect 368710 228308 368716 228320
rect 34072 228280 368716 228308
rect 34072 228268 34078 228280
rect 368710 228268 368716 228280
rect 368768 228268 368774 228320
rect 305138 227656 305144 227708
rect 305196 227696 305202 227708
rect 322986 227696 322992 227708
rect 305196 227668 322992 227696
rect 305196 227656 305202 227668
rect 322986 227656 322992 227668
rect 323044 227656 323050 227708
rect 345158 227656 345164 227708
rect 345216 227696 345222 227708
rect 360798 227696 360804 227708
rect 345216 227668 360804 227696
rect 345216 227656 345222 227668
rect 360798 227656 360804 227668
rect 360856 227656 360862 227708
rect 222430 227588 222436 227640
rect 222488 227628 222494 227640
rect 222614 227628 222620 227640
rect 222488 227600 222620 227628
rect 222488 227588 222494 227600
rect 222614 227588 222620 227600
rect 222672 227588 222678 227640
rect 280298 227588 280304 227640
rect 280356 227628 280362 227640
rect 353070 227628 353076 227640
rect 280356 227600 353076 227628
rect 280356 227588 280362 227600
rect 353070 227588 353076 227600
rect 353128 227588 353134 227640
rect 186458 227520 186464 227572
rect 186516 227560 186522 227572
rect 369262 227560 369268 227572
rect 186516 227532 369268 227560
rect 186516 227520 186522 227532
rect 369262 227520 369268 227532
rect 369320 227520 369326 227572
rect 325378 226976 325384 227028
rect 325436 227016 325442 227028
rect 325654 227016 325660 227028
rect 325436 226988 325660 227016
rect 325436 226976 325442 226988
rect 325654 226976 325660 226988
rect 325712 227016 325718 227028
rect 343870 227016 343876 227028
rect 325712 226988 343876 227016
rect 325712 226976 325718 226988
rect 343870 226976 343876 226988
rect 343928 227016 343934 227028
rect 345158 227016 345164 227028
rect 343928 226988 345164 227016
rect 343928 226976 343934 226988
rect 345158 226976 345164 226988
rect 345216 226976 345222 227028
rect 76794 226908 76800 226960
rect 76852 226948 76858 226960
rect 368802 226948 368808 226960
rect 76852 226920 368808 226948
rect 76852 226908 76858 226920
rect 368802 226908 368808 226920
rect 368860 226908 368866 226960
rect 34566 226840 34572 226892
rect 34624 226880 34630 226892
rect 368710 226880 368716 226892
rect 34624 226852 368716 226880
rect 34624 226840 34630 226852
rect 368710 226840 368716 226852
rect 368768 226840 368774 226892
rect 324734 226296 324740 226348
rect 324792 226336 324798 226348
rect 347182 226336 347188 226348
rect 324792 226308 347188 226336
rect 324792 226296 324798 226308
rect 347182 226296 347188 226308
rect 347240 226296 347246 226348
rect 239542 226228 239548 226280
rect 239600 226268 239606 226280
rect 353162 226268 353168 226280
rect 239600 226240 353168 226268
rect 239600 226228 239606 226240
rect 353162 226228 353168 226240
rect 353220 226228 353226 226280
rect 231354 226160 231360 226212
rect 231412 226200 231418 226212
rect 353254 226200 353260 226212
rect 231412 226172 353260 226200
rect 231412 226160 231418 226172
rect 353254 226160 353260 226172
rect 353312 226160 353318 226212
rect 137606 226092 137612 226144
rect 137664 226132 137670 226144
rect 353346 226132 353352 226144
rect 137664 226104 353352 226132
rect 137664 226092 137670 226104
rect 353346 226092 353352 226104
rect 353404 226092 353410 226144
rect 360430 225996 360436 226008
rect 360356 225968 360436 225996
rect 359694 225860 359700 225872
rect 350788 225832 359700 225860
rect 347182 225684 347188 225736
rect 347240 225724 347246 225736
rect 350788 225724 350816 225832
rect 359694 225820 359700 225832
rect 359752 225860 359758 225872
rect 360356 225860 360384 225968
rect 360430 225956 360436 225968
rect 360488 225956 360494 226008
rect 359752 225832 360384 225860
rect 359752 225820 359758 225832
rect 347240 225696 350816 225724
rect 347240 225684 347246 225696
rect 172014 225616 172020 225668
rect 172072 225656 172078 225668
rect 368802 225656 368808 225668
rect 172072 225628 368808 225656
rect 172072 225616 172078 225628
rect 368802 225616 368808 225628
rect 368860 225616 368866 225668
rect 137514 225548 137520 225600
rect 137572 225588 137578 225600
rect 368710 225588 368716 225600
rect 137572 225560 368716 225588
rect 137572 225548 137578 225560
rect 368710 225548 368716 225560
rect 368768 225548 368774 225600
rect 134754 225480 134760 225532
rect 134812 225520 134818 225532
rect 368894 225520 368900 225532
rect 134812 225492 368900 225520
rect 134812 225480 134818 225492
rect 368894 225480 368900 225492
rect 368952 225480 368958 225532
rect 158030 225412 158036 225464
rect 158088 225452 158094 225464
rect 159042 225452 159048 225464
rect 158088 225424 159048 225452
rect 158088 225412 158094 225424
rect 159042 225412 159048 225424
rect 159100 225412 159106 225464
rect 161986 225412 161992 225464
rect 162044 225452 162050 225464
rect 164378 225452 164384 225464
rect 162044 225424 164384 225452
rect 162044 225412 162050 225424
rect 164378 225412 164384 225424
rect 164436 225412 164442 225464
rect 251318 225412 251324 225464
rect 251376 225452 251382 225464
rect 253986 225452 253992 225464
rect 251376 225424 253992 225452
rect 251376 225412 251382 225424
rect 253986 225412 253992 225424
rect 254044 225412 254050 225464
rect 338350 225412 338356 225464
rect 338408 225452 338414 225464
rect 343502 225452 343508 225464
rect 338408 225424 343508 225452
rect 338408 225412 338414 225424
rect 343502 225412 343508 225424
rect 343560 225412 343566 225464
rect 345897 225455 345955 225461
rect 345897 225421 345909 225455
rect 345943 225452 345955 225455
rect 350954 225452 350960 225464
rect 345943 225424 350960 225452
rect 345943 225421 345955 225424
rect 345897 225415 345955 225421
rect 350954 225412 350960 225424
rect 351012 225412 351018 225464
rect 62994 225344 63000 225396
rect 63052 225384 63058 225396
rect 65938 225384 65944 225396
rect 63052 225356 65944 225384
rect 63052 225344 63058 225356
rect 65938 225344 65944 225356
rect 65996 225344 66002 225396
rect 67134 225344 67140 225396
rect 67192 225384 67198 225396
rect 69434 225384 69440 225396
rect 67192 225356 69440 225384
rect 67192 225344 67198 225356
rect 69434 225344 69440 225356
rect 69492 225344 69498 225396
rect 228686 225344 228692 225396
rect 228744 225384 228750 225396
rect 368710 225384 368716 225396
rect 228744 225356 368716 225384
rect 228744 225344 228750 225356
rect 368710 225344 368716 225356
rect 368768 225344 368774 225396
rect 56094 225276 56100 225328
rect 56152 225316 56158 225328
rect 56738 225316 56744 225328
rect 56152 225288 56744 225316
rect 56152 225276 56158 225288
rect 56738 225276 56744 225288
rect 56796 225276 56802 225328
rect 59682 225276 59688 225328
rect 59740 225316 59746 225328
rect 60878 225316 60884 225328
rect 59740 225288 60884 225316
rect 59740 225276 59746 225288
rect 60878 225276 60884 225288
rect 60936 225276 60942 225328
rect 61430 225276 61436 225328
rect 61488 225316 61494 225328
rect 62258 225316 62264 225328
rect 61488 225288 62264 225316
rect 61488 225276 61494 225288
rect 62258 225276 62264 225288
rect 62316 225276 62322 225328
rect 62350 225276 62356 225328
rect 62408 225316 62414 225328
rect 63638 225316 63644 225328
rect 62408 225288 63644 225316
rect 62408 225276 62414 225288
rect 63638 225276 63644 225288
rect 63696 225276 63702 225328
rect 65754 225276 65760 225328
rect 65812 225316 65818 225328
rect 66766 225316 66772 225328
rect 65812 225288 66772 225316
rect 65812 225276 65818 225288
rect 66766 225276 66772 225288
rect 66824 225276 66830 225328
rect 68514 225276 68520 225328
rect 68572 225316 68578 225328
rect 70354 225316 70360 225328
rect 68572 225288 70360 225316
rect 68572 225276 68578 225288
rect 70354 225276 70360 225288
rect 70412 225276 70418 225328
rect 137606 225276 137612 225328
rect 137664 225316 137670 225328
rect 368986 225316 368992 225328
rect 137664 225288 368992 225316
rect 137664 225276 137670 225288
rect 368986 225276 368992 225288
rect 369044 225276 369050 225328
rect 249202 225208 249208 225260
rect 249260 225248 249266 225260
rect 252146 225248 252152 225260
rect 249260 225220 252152 225248
rect 249260 225208 249266 225220
rect 252146 225208 252152 225220
rect 252204 225208 252210 225260
rect 337154 225208 337160 225260
rect 337212 225248 337218 225260
rect 341110 225248 341116 225260
rect 337212 225220 341116 225248
rect 337212 225208 337218 225220
rect 341110 225208 341116 225220
rect 341168 225208 341174 225260
rect 341202 225208 341208 225260
rect 341260 225248 341266 225260
rect 352242 225248 352248 225260
rect 341260 225220 352248 225248
rect 341260 225208 341266 225220
rect 352242 225208 352248 225220
rect 352300 225208 352306 225260
rect 65846 225140 65852 225192
rect 65904 225180 65910 225192
rect 67686 225180 67692 225192
rect 65904 225152 67692 225180
rect 65904 225140 65910 225152
rect 67686 225140 67692 225152
rect 67744 225140 67750 225192
rect 249754 225140 249760 225192
rect 249812 225180 249818 225192
rect 253066 225180 253072 225192
rect 249812 225152 253072 225180
rect 249812 225140 249818 225152
rect 253066 225140 253072 225152
rect 253124 225140 253130 225192
rect 338994 225140 339000 225192
rect 339052 225180 339058 225192
rect 341941 225183 341999 225189
rect 341941 225180 341953 225183
rect 339052 225152 341953 225180
rect 339052 225140 339058 225152
rect 341941 225149 341953 225152
rect 341987 225149 341999 225183
rect 341941 225143 341999 225149
rect 342030 225140 342036 225192
rect 342088 225180 342094 225192
rect 348102 225180 348108 225192
rect 342088 225152 348108 225180
rect 342088 225140 342094 225152
rect 348102 225140 348108 225152
rect 348160 225140 348166 225192
rect 63086 225072 63092 225124
rect 63144 225112 63150 225124
rect 64098 225112 64104 225124
rect 63144 225084 64104 225112
rect 63144 225072 63150 225084
rect 64098 225072 64104 225084
rect 64156 225072 64162 225124
rect 337706 225072 337712 225124
rect 337764 225112 337770 225124
rect 342490 225112 342496 225124
rect 337764 225084 342496 225112
rect 337764 225072 337770 225084
rect 342490 225072 342496 225084
rect 342548 225072 342554 225124
rect 347921 225115 347979 225121
rect 347921 225081 347933 225115
rect 347967 225112 347979 225115
rect 348013 225115 348071 225121
rect 348013 225112 348025 225115
rect 347967 225084 348025 225112
rect 347967 225081 347979 225084
rect 347921 225075 347979 225081
rect 348013 225081 348025 225084
rect 348059 225081 348071 225115
rect 348013 225075 348071 225081
rect 58762 225004 58768 225056
rect 58820 225044 58826 225056
rect 59498 225044 59504 225056
rect 58820 225016 59504 225044
rect 58820 225004 58826 225016
rect 59498 225004 59504 225016
rect 59556 225004 59562 225056
rect 335406 225004 335412 225056
rect 335464 225044 335470 225056
rect 348562 225044 348568 225056
rect 335464 225016 348568 225044
rect 335464 225004 335470 225016
rect 348562 225004 348568 225016
rect 348620 225004 348626 225056
rect 332738 224936 332744 224988
rect 332796 224976 332802 224988
rect 347274 224976 347280 224988
rect 332796 224948 347280 224976
rect 332796 224936 332802 224948
rect 347274 224936 347280 224948
rect 347332 224936 347338 224988
rect 360706 224936 360712 224988
rect 360764 224976 360770 224988
rect 361166 224976 361172 224988
rect 360764 224948 361172 224976
rect 360764 224936 360770 224948
rect 361166 224936 361172 224948
rect 361224 224936 361230 224988
rect 334118 224868 334124 224920
rect 334176 224908 334182 224920
rect 347918 224908 347924 224920
rect 334176 224880 347924 224908
rect 334176 224868 334182 224880
rect 347918 224868 347924 224880
rect 347976 224868 347982 224920
rect 335498 224800 335504 224852
rect 335556 224840 335562 224852
rect 349390 224840 349396 224852
rect 335556 224812 349396 224840
rect 335556 224800 335562 224812
rect 349390 224800 349396 224812
rect 349448 224800 349454 224852
rect 349500 224812 350816 224840
rect 57014 224732 57020 224784
rect 57072 224772 57078 224784
rect 67318 224772 67324 224784
rect 57072 224744 67324 224772
rect 57072 224732 57078 224744
rect 67318 224732 67324 224744
rect 67376 224732 67382 224784
rect 339638 224732 339644 224784
rect 339696 224772 339702 224784
rect 345897 224775 345955 224781
rect 345897 224772 345909 224775
rect 339696 224744 345909 224772
rect 339696 224732 339702 224744
rect 345897 224741 345909 224744
rect 345943 224741 345955 224775
rect 345897 224735 345955 224741
rect 348013 224775 348071 224781
rect 348013 224741 348025 224775
rect 348059 224772 348071 224775
rect 349500 224772 349528 224812
rect 348059 224744 349528 224772
rect 350788 224772 350816 224812
rect 358038 224800 358044 224852
rect 358096 224840 358102 224852
rect 358222 224840 358228 224852
rect 358096 224812 358228 224840
rect 358096 224800 358102 224812
rect 358222 224800 358228 224812
rect 358280 224800 358286 224852
rect 360982 224772 360988 224784
rect 350788 224744 360988 224772
rect 348059 224741 348071 224744
rect 348013 224735 348071 224741
rect 360982 224732 360988 224744
rect 361040 224732 361046 224784
rect 339546 224664 339552 224716
rect 339604 224704 339610 224716
rect 341941 224707 341999 224713
rect 339604 224676 341892 224704
rect 339604 224664 339610 224676
rect 341864 224636 341892 224676
rect 341941 224673 341953 224707
rect 341987 224704 341999 224707
rect 342674 224704 342680 224716
rect 341987 224676 342680 224704
rect 341987 224673 341999 224676
rect 341941 224667 341999 224673
rect 342674 224664 342680 224676
rect 342732 224664 342738 224716
rect 345342 224636 345348 224648
rect 341864 224608 345348 224636
rect 345342 224596 345348 224608
rect 345400 224596 345406 224648
rect 336878 224528 336884 224580
rect 336936 224568 336942 224580
rect 349758 224568 349764 224580
rect 336936 224540 349764 224568
rect 336936 224528 336942 224540
rect 349758 224528 349764 224540
rect 349816 224528 349822 224580
rect 341386 224460 341392 224512
rect 341444 224500 341450 224512
rect 348010 224500 348016 224512
rect 341444 224472 348016 224500
rect 341444 224460 341450 224472
rect 348010 224460 348016 224472
rect 348068 224460 348074 224512
rect 338258 224392 338264 224444
rect 338316 224432 338322 224444
rect 350678 224432 350684 224444
rect 338316 224404 350684 224432
rect 338316 224392 338322 224404
rect 350678 224392 350684 224404
rect 350736 224392 350742 224444
rect 339454 224324 339460 224376
rect 339512 224364 339518 224376
rect 351598 224364 351604 224376
rect 339512 224336 351604 224364
rect 339512 224324 339518 224336
rect 351598 224324 351604 224336
rect 351656 224324 351662 224376
rect 63178 224256 63184 224308
rect 63236 224296 63242 224308
rect 65018 224296 65024 224308
rect 63236 224268 65024 224296
rect 63236 224256 63242 224268
rect 65018 224256 65024 224268
rect 65076 224256 65082 224308
rect 67226 224256 67232 224308
rect 67284 224296 67290 224308
rect 68606 224296 68612 224308
rect 67284 224268 68612 224296
rect 67284 224256 67290 224268
rect 68606 224256 68612 224268
rect 68664 224256 68670 224308
rect 325838 224256 325844 224308
rect 325896 224296 325902 224308
rect 345158 224296 345164 224308
rect 325896 224268 345164 224296
rect 325896 224256 325902 224268
rect 345158 224256 345164 224268
rect 345216 224256 345222 224308
rect 61614 224188 61620 224240
rect 61672 224228 61678 224240
rect 63270 224228 63276 224240
rect 61672 224200 63276 224228
rect 61672 224188 61678 224200
rect 63270 224188 63276 224200
rect 63328 224188 63334 224240
rect 324918 224188 324924 224240
rect 324976 224228 324982 224240
rect 325194 224228 325200 224240
rect 324976 224200 325200 224228
rect 324976 224188 324982 224200
rect 325194 224188 325200 224200
rect 325252 224228 325258 224240
rect 344514 224228 344520 224240
rect 325252 224200 344520 224228
rect 325252 224188 325258 224200
rect 344514 224188 344520 224200
rect 344572 224228 344578 224240
rect 361166 224228 361172 224240
rect 344572 224200 361172 224228
rect 344572 224188 344578 224200
rect 361166 224188 361172 224200
rect 361224 224188 361230 224240
rect 322526 224120 322532 224172
rect 322584 224160 322590 224172
rect 368802 224160 368808 224172
rect 322584 224132 368808 224160
rect 322584 224120 322590 224132
rect 368802 224120 368808 224132
rect 368860 224120 368866 224172
rect 369170 224160 369176 224172
rect 369131 224132 369176 224160
rect 369170 224120 369176 224132
rect 369228 224120 369234 224172
rect 369078 223984 369084 224036
rect 369136 224024 369142 224036
rect 369354 224024 369360 224036
rect 369136 223996 369360 224024
rect 369136 223984 369142 223996
rect 369354 223984 369360 223996
rect 369412 223984 369418 224036
rect 342720 223032 342726 223084
rect 342778 223072 342784 223084
rect 347921 223075 347979 223081
rect 347921 223072 347933 223075
rect 342778 223044 347933 223072
rect 342778 223032 342784 223044
rect 347921 223041 347933 223044
rect 347967 223041 347979 223075
rect 347921 223035 347979 223041
rect 325562 222896 325568 222948
rect 325620 222936 325626 222948
rect 342720 222936 342726 222948
rect 325620 222908 342726 222936
rect 325620 222896 325626 222908
rect 342720 222896 342726 222908
rect 342778 222896 342784 222948
rect 362454 222896 362460 222948
rect 362512 222936 362518 222948
rect 369078 222936 369084 222948
rect 362512 222908 369084 222936
rect 362512 222896 362518 222908
rect 369078 222896 369084 222908
rect 369136 222896 369142 222948
rect 323814 222828 323820 222880
rect 323872 222868 323878 222880
rect 368710 222868 368716 222880
rect 323872 222840 368716 222868
rect 323872 222828 323878 222840
rect 368710 222828 368716 222840
rect 368768 222828 368774 222880
rect 322618 222760 322624 222812
rect 322676 222800 322682 222812
rect 368802 222800 368808 222812
rect 322676 222772 368808 222800
rect 322676 222760 322682 222772
rect 368802 222760 368808 222772
rect 368860 222760 368866 222812
rect 38522 222012 38528 222064
rect 38580 222052 38586 222064
rect 50574 222052 50580 222064
rect 38580 222024 50580 222052
rect 38580 222012 38586 222024
rect 50574 222012 50580 222024
rect 50632 222012 50638 222064
rect 34566 221740 34572 221792
rect 34624 221780 34630 221792
rect 34934 221780 34940 221792
rect 34624 221752 34940 221780
rect 34624 221740 34630 221752
rect 34934 221740 34940 221752
rect 34992 221740 34998 221792
rect 34014 221672 34020 221724
rect 34072 221712 34078 221724
rect 34750 221712 34756 221724
rect 34072 221684 34756 221712
rect 34072 221672 34078 221684
rect 34750 221672 34756 221684
rect 34808 221672 34814 221724
rect 361074 221468 361080 221520
rect 361132 221508 361138 221520
rect 369078 221508 369084 221520
rect 361132 221480 369084 221508
rect 361132 221468 361138 221480
rect 369078 221468 369084 221480
rect 369136 221468 369142 221520
rect 325194 221400 325200 221452
rect 325252 221440 325258 221452
rect 368802 221440 368808 221452
rect 325252 221412 368808 221440
rect 325252 221400 325258 221412
rect 368802 221400 368808 221412
rect 368860 221400 368866 221452
rect 322802 221332 322808 221384
rect 322860 221372 322866 221384
rect 368710 221372 368716 221384
rect 322860 221344 368716 221372
rect 322860 221332 322866 221344
rect 368710 221332 368716 221344
rect 368768 221332 368774 221384
rect 369906 221372 369912 221384
rect 369867 221344 369912 221372
rect 369906 221332 369912 221344
rect 369964 221332 369970 221384
rect 325286 220584 325292 220636
rect 325344 220624 325350 220636
rect 353438 220624 353444 220636
rect 325344 220596 353444 220624
rect 325344 220584 325350 220596
rect 353438 220584 353444 220596
rect 353496 220584 353502 220636
rect 34658 220516 34664 220568
rect 34716 220556 34722 220568
rect 34934 220556 34940 220568
rect 34716 220528 34940 220556
rect 34716 220516 34722 220528
rect 34934 220516 34940 220528
rect 34992 220516 34998 220568
rect 325378 220516 325384 220568
rect 325436 220556 325442 220568
rect 368802 220556 368808 220568
rect 325436 220528 368808 220556
rect 325436 220516 325442 220528
rect 368802 220516 368808 220528
rect 368860 220516 368866 220568
rect 34750 220448 34756 220500
rect 34808 220488 34814 220500
rect 34845 220491 34903 220497
rect 34845 220488 34857 220491
rect 34808 220460 34857 220488
rect 34808 220448 34814 220460
rect 34845 220457 34857 220460
rect 34891 220457 34903 220491
rect 34845 220451 34903 220457
rect 322710 220448 322716 220500
rect 322768 220488 322774 220500
rect 368710 220488 368716 220500
rect 322768 220460 368716 220488
rect 322768 220448 322774 220460
rect 368710 220448 368716 220460
rect 368768 220448 368774 220500
rect 359786 220040 359792 220092
rect 359844 220080 359850 220092
rect 368986 220080 368992 220092
rect 359844 220052 368992 220080
rect 359844 220040 359850 220052
rect 368986 220040 368992 220052
rect 369044 220040 369050 220092
rect 38062 219904 38068 219956
rect 38120 219944 38126 219956
rect 52046 219944 52052 219956
rect 38120 219916 52052 219944
rect 38120 219904 38126 219916
rect 52046 219904 52052 219916
rect 52104 219904 52110 219956
rect 76150 219496 76156 219548
rect 76208 219536 76214 219548
rect 81670 219536 81676 219548
rect 76208 219508 81676 219536
rect 76208 219496 76214 219508
rect 81670 219496 81676 219508
rect 81728 219496 81734 219548
rect 165114 219224 165120 219276
rect 165172 219264 165178 219276
rect 178914 219264 178920 219276
rect 165172 219236 178920 219264
rect 165172 219224 165178 219236
rect 178914 219224 178920 219236
rect 178972 219224 178978 219276
rect 258954 219224 258960 219276
rect 259012 219264 259018 219276
rect 272938 219264 272944 219276
rect 259012 219236 272944 219264
rect 259012 219224 259018 219236
rect 272938 219224 272944 219236
rect 272996 219224 273002 219276
rect 365214 218680 365220 218732
rect 365272 218720 365278 218732
rect 368802 218720 368808 218732
rect 365272 218692 368808 218720
rect 365272 218680 365278 218692
rect 368802 218680 368808 218692
rect 368860 218680 368866 218732
rect 352794 218612 352800 218664
rect 352852 218652 352858 218664
rect 368710 218652 368716 218664
rect 352852 218624 368716 218652
rect 352852 218612 352858 218624
rect 368710 218612 368716 218624
rect 368768 218612 368774 218664
rect 394838 218612 394844 218664
rect 394896 218652 394902 218664
rect 405970 218652 405976 218664
rect 394896 218624 405976 218652
rect 394896 218612 394902 218624
rect 405970 218612 405976 218624
rect 406028 218612 406034 218664
rect 352886 218544 352892 218596
rect 352944 218584 352950 218596
rect 368802 218584 368808 218596
rect 352944 218556 368808 218584
rect 352944 218544 352950 218556
rect 368802 218544 368808 218556
rect 368860 218544 368866 218596
rect 352978 217184 352984 217236
rect 353036 217224 353042 217236
rect 368710 217224 368716 217236
rect 353036 217196 368716 217224
rect 353036 217184 353042 217196
rect 368710 217184 368716 217196
rect 368768 217184 368774 217236
rect 38522 217116 38528 217168
rect 38580 217156 38586 217168
rect 53242 217156 53248 217168
rect 38580 217128 53248 217156
rect 38580 217116 38586 217128
rect 53242 217116 53248 217128
rect 53300 217116 53306 217168
rect 353346 217048 353352 217100
rect 353404 217088 353410 217100
rect 368710 217088 368716 217100
rect 353404 217060 368716 217088
rect 353404 217048 353410 217060
rect 368710 217048 368716 217060
rect 368768 217048 368774 217100
rect 368986 216436 368992 216488
rect 369044 216476 369050 216488
rect 369173 216479 369231 216485
rect 369173 216476 369185 216479
rect 369044 216448 369185 216476
rect 369044 216436 369050 216448
rect 369173 216445 369185 216448
rect 369219 216445 369231 216479
rect 369173 216439 369231 216445
rect 137698 215824 137704 215876
rect 137756 215864 137762 215876
rect 145150 215864 145156 215876
rect 137756 215836 145156 215864
rect 137756 215824 137762 215836
rect 145150 215824 145156 215836
rect 145208 215824 145214 215876
rect 231354 215824 231360 215876
rect 231412 215864 231418 215876
rect 240922 215864 240928 215876
rect 231412 215836 240928 215864
rect 231412 215824 231418 215836
rect 240922 215824 240928 215836
rect 240980 215824 240986 215876
rect 325286 215824 325292 215876
rect 325344 215864 325350 215876
rect 334210 215864 334216 215876
rect 325344 215836 334216 215864
rect 325344 215824 325350 215836
rect 334210 215824 334216 215836
rect 334268 215824 334274 215876
rect 353162 215756 353168 215808
rect 353220 215796 353226 215808
rect 368710 215796 368716 215808
rect 353220 215768 368716 215796
rect 353220 215756 353226 215768
rect 368710 215756 368716 215768
rect 368768 215756 368774 215808
rect 427314 215756 427320 215808
rect 427372 215796 427378 215808
rect 429706 215796 429712 215808
rect 427372 215768 429712 215796
rect 427372 215756 427378 215768
rect 429706 215756 429712 215768
rect 429764 215756 429770 215808
rect 353254 215688 353260 215740
rect 353312 215728 353318 215740
rect 368802 215728 368808 215740
rect 353312 215700 368808 215728
rect 353312 215688 353318 215700
rect 368802 215688 368808 215700
rect 368860 215688 368866 215740
rect 358406 215620 358412 215672
rect 358464 215660 358470 215672
rect 368710 215660 368716 215672
rect 358464 215632 368716 215660
rect 358464 215620 358470 215632
rect 368710 215620 368716 215632
rect 368768 215620 368774 215672
rect 358222 215484 358228 215536
rect 358280 215524 358286 215536
rect 358406 215524 358412 215536
rect 358280 215496 358412 215524
rect 358280 215484 358286 215496
rect 358406 215484 358412 215496
rect 358464 215484 358470 215536
rect 368986 214464 368992 214516
rect 369044 214504 369050 214516
rect 369170 214504 369176 214516
rect 369044 214476 369176 214504
rect 369044 214464 369050 214476
rect 369170 214464 369176 214476
rect 369228 214464 369234 214516
rect 38522 214396 38528 214448
rect 38580 214436 38586 214448
rect 51402 214436 51408 214448
rect 38580 214408 51408 214436
rect 38580 214396 38586 214408
rect 51402 214396 51408 214408
rect 51460 214396 51466 214448
rect 353070 214260 353076 214312
rect 353128 214300 353134 214312
rect 368710 214300 368716 214312
rect 353128 214272 368716 214300
rect 353128 214260 353134 214272
rect 368710 214260 368716 214272
rect 368768 214260 368774 214312
rect 361258 214192 361264 214244
rect 361316 214232 361322 214244
rect 368894 214232 368900 214244
rect 361316 214204 368900 214232
rect 361316 214192 361322 214204
rect 368894 214192 368900 214204
rect 368952 214192 368958 214244
rect 356198 214056 356204 214108
rect 356256 214096 356262 214108
rect 405970 214096 405976 214108
rect 356256 214068 405976 214096
rect 356256 214056 356262 214068
rect 405970 214056 405976 214068
rect 406028 214056 406034 214108
rect 357670 213988 357676 214040
rect 357728 214028 357734 214040
rect 406614 214028 406620 214040
rect 357728 214000 406620 214028
rect 357728 213988 357734 214000
rect 406614 213988 406620 214000
rect 406672 213988 406678 214040
rect 355094 213920 355100 213972
rect 355152 213960 355158 213972
rect 394838 213960 394844 213972
rect 355152 213932 394844 213960
rect 355152 213920 355158 213932
rect 394838 213920 394844 213932
rect 394896 213920 394902 213972
rect 34842 213892 34848 213904
rect 34803 213864 34848 213892
rect 34842 213852 34848 213864
rect 34900 213852 34906 213904
rect 353438 213036 353444 213088
rect 353496 213076 353502 213088
rect 368710 213076 368716 213088
rect 353496 213048 368716 213076
rect 353496 213036 353502 213048
rect 368710 213036 368716 213048
rect 368768 213036 368774 213088
rect 369906 211608 369912 211660
rect 369964 211648 369970 211660
rect 370734 211648 370740 211660
rect 369964 211620 370740 211648
rect 369964 211608 369970 211620
rect 370734 211608 370740 211620
rect 370792 211608 370798 211660
rect 38706 210928 38712 210980
rect 38764 210968 38770 210980
rect 54070 210968 54076 210980
rect 38764 210940 54076 210968
rect 38764 210928 38770 210940
rect 54070 210928 54076 210940
rect 54128 210928 54134 210980
rect 354910 210928 354916 210980
rect 354968 210968 354974 210980
rect 405970 210968 405976 210980
rect 354968 210940 405976 210968
rect 354968 210928 354974 210940
rect 405970 210928 405976 210940
rect 406028 210928 406034 210980
rect 383890 210860 383896 210912
rect 383948 210900 383954 210912
rect 385178 210900 385184 210912
rect 383948 210872 385184 210900
rect 383948 210860 383954 210872
rect 385178 210860 385184 210872
rect 385236 210860 385242 210912
rect 369538 209636 369544 209688
rect 369596 209676 369602 209688
rect 369906 209676 369912 209688
rect 369596 209648 369912 209676
rect 369596 209636 369602 209648
rect 369906 209636 369912 209648
rect 369964 209636 369970 209688
rect 38522 209568 38528 209620
rect 38580 209608 38586 209620
rect 51402 209608 51408 209620
rect 38580 209580 51408 209608
rect 38580 209568 38586 209580
rect 51402 209568 51408 209580
rect 51460 209568 51466 209620
rect 356198 209568 356204 209620
rect 356256 209608 356262 209620
rect 405970 209608 405976 209620
rect 356256 209580 405976 209608
rect 356256 209568 356262 209580
rect 405970 209568 405976 209580
rect 406028 209568 406034 209620
rect 34842 206888 34848 206900
rect 34803 206860 34848 206888
rect 34842 206848 34848 206860
rect 34900 206848 34906 206900
rect 38522 206780 38528 206832
rect 38580 206820 38586 206832
rect 51402 206820 51408 206832
rect 38580 206792 51408 206820
rect 38580 206780 38586 206792
rect 51402 206780 51408 206792
rect 51460 206780 51466 206832
rect 355002 206780 355008 206832
rect 355060 206820 355066 206832
rect 405970 206820 405976 206832
rect 355060 206792 405976 206820
rect 355060 206780 355066 206792
rect 405970 206780 405976 206792
rect 406028 206780 406034 206832
rect 38522 204740 38528 204792
rect 38580 204780 38586 204792
rect 51402 204780 51408 204792
rect 38580 204752 51408 204780
rect 38580 204740 38586 204752
rect 51402 204740 51408 204752
rect 51460 204740 51466 204792
rect 136870 204740 136876 204792
rect 136928 204780 136934 204792
rect 145334 204780 145340 204792
rect 136928 204752 145340 204780
rect 136928 204740 136934 204752
rect 145334 204740 145340 204752
rect 145392 204740 145398 204792
rect 356198 204740 356204 204792
rect 356256 204780 356262 204792
rect 406062 204780 406068 204792
rect 356256 204752 406068 204780
rect 356256 204740 356262 204752
rect 406062 204740 406068 204752
rect 406120 204740 406126 204792
rect 34842 204712 34848 204724
rect 34803 204684 34848 204712
rect 34842 204672 34848 204684
rect 34900 204672 34906 204724
rect 368986 204672 368992 204724
rect 369044 204712 369050 204724
rect 369170 204712 369176 204724
rect 369044 204684 369176 204712
rect 369044 204672 369050 204684
rect 369170 204672 369176 204684
rect 369228 204672 369234 204724
rect 231630 204060 231636 204112
rect 231688 204100 231694 204112
rect 237518 204100 237524 204112
rect 231688 204072 237524 204100
rect 231688 204060 231694 204072
rect 237518 204060 237524 204072
rect 237576 204060 237582 204112
rect 74218 203312 74224 203364
rect 74276 203352 74282 203364
rect 81670 203352 81676 203364
rect 74276 203324 81676 203352
rect 74276 203312 74282 203324
rect 81670 203312 81676 203324
rect 81728 203312 81734 203364
rect 167874 203312 167880 203364
rect 167932 203352 167938 203364
rect 178914 203352 178920 203364
rect 167932 203324 178920 203352
rect 167932 203312 167938 203324
rect 178914 203312 178920 203324
rect 178972 203312 178978 203364
rect 261714 203312 261720 203364
rect 261772 203352 261778 203364
rect 272938 203352 272944 203364
rect 261772 203324 272944 203352
rect 261772 203312 261778 203324
rect 272938 203312 272944 203324
rect 272996 203312 273002 203364
rect 13958 202020 13964 202072
rect 14016 202060 14022 202072
rect 16442 202060 16448 202072
rect 14016 202032 16448 202060
rect 14016 202020 14022 202032
rect 16442 202020 16448 202032
rect 16500 202020 16506 202072
rect 137790 202020 137796 202072
rect 137848 202060 137854 202072
rect 145150 202060 145156 202072
rect 137848 202032 145156 202060
rect 137848 202020 137854 202032
rect 145150 202020 145156 202032
rect 145208 202020 145214 202072
rect 231446 202020 231452 202072
rect 231504 202060 231510 202072
rect 240370 202060 240376 202072
rect 231504 202032 240376 202060
rect 231504 202020 231510 202032
rect 240370 202020 240376 202032
rect 240428 202020 240434 202072
rect 325470 202020 325476 202072
rect 325528 202060 325534 202072
rect 334210 202060 334216 202072
rect 325528 202032 334216 202060
rect 325528 202020 325534 202032
rect 334210 202020 334216 202032
rect 334268 202020 334274 202072
rect 358406 202020 358412 202072
rect 358464 202060 358470 202072
rect 358590 202060 358596 202072
rect 358464 202032 358596 202060
rect 358464 202020 358470 202032
rect 358590 202020 358596 202032
rect 358648 202020 358654 202072
rect 38522 201272 38528 201324
rect 38580 201312 38586 201324
rect 51494 201312 51500 201324
rect 38580 201284 51500 201312
rect 38580 201272 38586 201284
rect 51494 201272 51500 201284
rect 51552 201272 51558 201324
rect 353530 201272 353536 201324
rect 353588 201312 353594 201324
rect 405970 201312 405976 201324
rect 353588 201284 405976 201312
rect 353588 201272 353594 201284
rect 405970 201272 405976 201284
rect 406028 201272 406034 201324
rect 369538 199912 369544 199964
rect 369596 199952 369602 199964
rect 369906 199952 369912 199964
rect 369596 199924 369912 199952
rect 369596 199912 369602 199924
rect 369906 199912 369912 199924
rect 369964 199912 369970 199964
rect 427130 199708 427136 199760
rect 427188 199748 427194 199760
rect 428786 199748 428792 199760
rect 427188 199720 428792 199748
rect 427188 199708 427194 199720
rect 428786 199708 428792 199720
rect 428844 199708 428850 199760
rect 13406 199300 13412 199352
rect 13464 199340 13470 199352
rect 17638 199340 17644 199352
rect 13464 199312 17644 199340
rect 13464 199300 13470 199312
rect 17638 199300 17644 199312
rect 17696 199300 17702 199352
rect 38522 199232 38528 199284
rect 38580 199272 38586 199284
rect 51218 199272 51224 199284
rect 38580 199244 51224 199272
rect 38580 199232 38586 199244
rect 51218 199232 51224 199244
rect 51276 199232 51282 199284
rect 356198 199232 356204 199284
rect 356256 199272 356262 199284
rect 405970 199272 405976 199284
rect 356256 199244 405976 199272
rect 356256 199232 356262 199244
rect 405970 199232 405976 199244
rect 406028 199232 406034 199284
rect 38522 195764 38528 195816
rect 38580 195804 38586 195816
rect 51310 195804 51316 195816
rect 38580 195776 51316 195804
rect 38580 195764 38586 195776
rect 51310 195764 51316 195776
rect 51368 195764 51374 195816
rect 352702 195764 352708 195816
rect 352760 195804 352766 195816
rect 405970 195804 405976 195816
rect 352760 195776 405976 195804
rect 352760 195764 352766 195776
rect 405970 195764 405976 195776
rect 406028 195764 406034 195816
rect 368713 195263 368771 195269
rect 368713 195229 368725 195263
rect 368759 195260 368771 195263
rect 368802 195260 368808 195272
rect 368759 195232 368808 195260
rect 368759 195229 368771 195232
rect 368713 195223 368771 195229
rect 368802 195220 368808 195232
rect 368860 195220 368866 195272
rect 51310 195192 51316 195204
rect 48476 195164 51316 195192
rect 38798 195084 38804 195136
rect 38856 195124 38862 195136
rect 48476 195124 48504 195164
rect 51310 195152 51316 195164
rect 51368 195152 51374 195204
rect 369078 195152 369084 195204
rect 369136 195192 369142 195204
rect 369354 195192 369360 195204
rect 369136 195164 369360 195192
rect 369136 195152 369142 195164
rect 369354 195152 369360 195164
rect 369412 195152 369418 195204
rect 38856 195096 48504 195124
rect 38856 195084 38862 195096
rect 356198 195084 356204 195136
rect 356256 195124 356262 195136
rect 406062 195124 406068 195136
rect 356256 195096 406068 195124
rect 356256 195084 356262 195096
rect 406062 195084 406068 195096
rect 406120 195084 406126 195136
rect 167966 192568 167972 192620
rect 168024 192608 168030 192620
rect 173394 192608 173400 192620
rect 168024 192580 173400 192608
rect 168024 192568 168030 192580
rect 173394 192568 173400 192580
rect 173452 192568 173458 192620
rect 262358 192364 262364 192416
rect 262416 192404 262422 192416
rect 273122 192404 273128 192416
rect 262416 192376 273128 192404
rect 262416 192364 262422 192376
rect 273122 192364 273128 192376
rect 273180 192364 273186 192416
rect 368710 192404 368716 192416
rect 368671 192376 368716 192404
rect 368710 192364 368716 192376
rect 368768 192364 368774 192416
rect 38798 191616 38804 191668
rect 38856 191656 38862 191668
rect 49930 191656 49936 191668
rect 38856 191628 49936 191656
rect 38856 191616 38862 191628
rect 49930 191616 49936 191628
rect 49988 191616 49994 191668
rect 173394 191616 173400 191668
rect 173452 191656 173458 191668
rect 178914 191656 178920 191668
rect 173452 191628 178920 191656
rect 173452 191616 173458 191628
rect 178914 191616 178920 191628
rect 178972 191616 178978 191668
rect 352794 191616 352800 191668
rect 352852 191656 352858 191668
rect 405970 191656 405976 191668
rect 352852 191628 405976 191656
rect 352852 191616 352858 191628
rect 405970 191616 405976 191628
rect 406028 191616 406034 191668
rect 368986 190256 368992 190308
rect 369044 190296 369050 190308
rect 369354 190296 369360 190308
rect 369044 190268 369360 190296
rect 369044 190256 369050 190268
rect 369354 190256 369360 190268
rect 369412 190256 369418 190308
rect 369538 190256 369544 190308
rect 369596 190296 369602 190308
rect 369906 190296 369912 190308
rect 369596 190268 369912 190296
rect 369596 190256 369602 190268
rect 369906 190256 369912 190268
rect 369964 190256 369970 190308
rect 13314 189576 13320 189628
rect 13372 189616 13378 189628
rect 13498 189616 13504 189628
rect 13372 189588 13504 189616
rect 13372 189576 13378 189588
rect 13498 189576 13504 189588
rect 13556 189576 13562 189628
rect 38062 189576 38068 189628
rect 38120 189616 38126 189628
rect 51218 189616 51224 189628
rect 38120 189588 51224 189616
rect 38120 189576 38126 189588
rect 51218 189576 51224 189588
rect 51276 189576 51282 189628
rect 137330 189576 137336 189628
rect 137388 189616 137394 189628
rect 137698 189616 137704 189628
rect 137388 189588 137704 189616
rect 137388 189576 137394 189588
rect 137698 189576 137704 189588
rect 137756 189576 137762 189628
rect 356198 189576 356204 189628
rect 356256 189616 356262 189628
rect 405970 189616 405976 189628
rect 356256 189588 405976 189616
rect 356256 189576 356262 189588
rect 405970 189576 405976 189588
rect 406028 189576 406034 189628
rect 13314 189372 13320 189424
rect 13372 189412 13378 189424
rect 17454 189412 17460 189424
rect 13372 189384 17460 189412
rect 13372 189372 13378 189384
rect 17454 189372 17460 189384
rect 17512 189372 17518 189424
rect 324550 188896 324556 188948
rect 324608 188936 324614 188948
rect 330070 188936 330076 188948
rect 324608 188908 330076 188936
rect 324608 188896 324614 188908
rect 330070 188896 330076 188908
rect 330128 188896 330134 188948
rect 231998 188760 232004 188812
rect 232056 188800 232062 188812
rect 236230 188800 236236 188812
rect 232056 188772 236236 188800
rect 232056 188760 232062 188772
rect 236230 188760 236236 188772
rect 236288 188800 236294 188812
rect 236874 188800 236880 188812
rect 236288 188772 236880 188800
rect 236288 188760 236294 188772
rect 236874 188760 236880 188772
rect 236932 188760 236938 188812
rect 137790 188284 137796 188336
rect 137848 188324 137854 188336
rect 142390 188324 142396 188336
rect 137848 188296 142396 188324
rect 137848 188284 137854 188296
rect 142390 188284 142396 188296
rect 142448 188324 142454 188336
rect 143034 188324 143040 188336
rect 142448 188296 143040 188324
rect 142448 188284 142454 188296
rect 143034 188284 143040 188296
rect 143092 188284 143098 188336
rect 232734 188284 232740 188336
rect 232792 188324 232798 188336
rect 240370 188324 240376 188336
rect 232792 188296 240376 188324
rect 232792 188284 232798 188296
rect 240370 188284 240376 188296
rect 240428 188284 240434 188336
rect 138894 188216 138900 188268
rect 138952 188256 138958 188268
rect 145610 188256 145616 188268
rect 138952 188228 145616 188256
rect 138952 188216 138958 188228
rect 145610 188216 145616 188228
rect 145668 188216 145674 188268
rect 326574 188216 326580 188268
rect 326632 188256 326638 188268
rect 334210 188256 334216 188268
rect 326632 188228 334216 188256
rect 326632 188216 326638 188228
rect 334210 188216 334216 188228
rect 334268 188216 334274 188268
rect 75414 186788 75420 186840
rect 75472 186828 75478 186840
rect 81670 186828 81676 186840
rect 75472 186800 81676 186828
rect 75472 186788 75478 186800
rect 81670 186788 81676 186800
rect 81728 186788 81734 186840
rect 38062 186108 38068 186160
rect 38120 186148 38126 186160
rect 48550 186148 48556 186160
rect 38120 186120 48556 186148
rect 38120 186108 38126 186120
rect 48550 186108 48556 186120
rect 48608 186108 48614 186160
rect 352794 186108 352800 186160
rect 352852 186148 352858 186160
rect 405970 186148 405976 186160
rect 352852 186120 405976 186148
rect 352852 186108 352858 186120
rect 405970 186108 405976 186120
rect 406028 186108 406034 186160
rect 368710 185496 368716 185548
rect 368768 185496 368774 185548
rect 13498 185428 13504 185480
rect 13556 185468 13562 185480
rect 17454 185468 17460 185480
rect 13556 185440 17460 185468
rect 13556 185428 13562 185440
rect 17454 185428 17460 185440
rect 17512 185428 17518 185480
rect 368728 185400 368756 185496
rect 427222 185428 427228 185480
rect 427280 185468 427286 185480
rect 430074 185468 430080 185480
rect 427280 185440 430080 185468
rect 427280 185428 427286 185440
rect 430074 185428 430080 185440
rect 430132 185428 430138 185480
rect 368802 185400 368808 185412
rect 368728 185372 368808 185400
rect 368802 185360 368808 185372
rect 368860 185360 368866 185412
rect 38798 184000 38804 184052
rect 38856 184040 38862 184052
rect 51402 184040 51408 184052
rect 38856 184012 51408 184040
rect 38856 184000 38862 184012
rect 51402 184000 51408 184012
rect 51460 184000 51466 184052
rect 356198 184000 356204 184052
rect 356256 184040 356262 184052
rect 405970 184040 405976 184052
rect 356256 184012 405976 184040
rect 356256 184000 356262 184012
rect 405970 184000 405976 184012
rect 406028 184000 406034 184052
rect 34382 183184 34388 183236
rect 34440 183224 34446 183236
rect 34934 183224 34940 183236
rect 34440 183196 34940 183224
rect 34440 183184 34446 183196
rect 34934 183184 34940 183196
rect 34992 183184 34998 183236
rect 34566 182640 34572 182692
rect 34624 182680 34630 182692
rect 34750 182680 34756 182692
rect 34624 182652 34756 182680
rect 34624 182640 34630 182652
rect 34750 182640 34756 182652
rect 34808 182640 34814 182692
rect 348013 181731 348071 181737
rect 348013 181697 348025 181731
rect 348059 181728 348071 181731
rect 352150 181728 352156 181740
rect 348059 181700 352156 181728
rect 348059 181697 348071 181700
rect 348013 181691 348071 181697
rect 352150 181688 352156 181700
rect 352208 181688 352214 181740
rect 21594 181280 21600 181332
rect 21652 181320 21658 181332
rect 34382 181320 34388 181332
rect 21652 181292 34388 181320
rect 21652 181280 21658 181292
rect 34382 181280 34388 181292
rect 34440 181280 34446 181332
rect 59682 181280 59688 181332
rect 59740 181320 59746 181332
rect 60878 181320 60884 181332
rect 59740 181292 60884 181320
rect 59740 181280 59746 181292
rect 60878 181280 60884 181292
rect 60936 181280 60942 181332
rect 61430 181280 61436 181332
rect 61488 181320 61494 181332
rect 62258 181320 62264 181332
rect 61488 181292 62264 181320
rect 61488 181280 61494 181292
rect 62258 181280 62264 181292
rect 62316 181280 62322 181332
rect 62994 181280 63000 181332
rect 63052 181320 63058 181332
rect 64098 181320 64104 181332
rect 63052 181292 64104 181320
rect 63052 181280 63058 181292
rect 64098 181280 64104 181292
rect 64156 181280 64162 181332
rect 65754 181280 65760 181332
rect 65812 181320 65818 181332
rect 66766 181320 66772 181332
rect 65812 181292 66772 181320
rect 65812 181280 65818 181292
rect 66766 181280 66772 181292
rect 66824 181280 66830 181332
rect 151038 181280 151044 181332
rect 151096 181320 151102 181332
rect 151866 181320 151872 181332
rect 151096 181292 151872 181320
rect 151096 181280 151102 181292
rect 151866 181280 151872 181292
rect 151924 181280 151930 181332
rect 152234 181280 152240 181332
rect 152292 181320 152298 181332
rect 153246 181320 153252 181332
rect 152292 181292 153252 181320
rect 152292 181280 152298 181292
rect 153246 181280 153252 181292
rect 153304 181280 153310 181332
rect 153430 181280 153436 181332
rect 153488 181320 153494 181332
rect 154718 181320 154724 181332
rect 153488 181292 154724 181320
rect 153488 181280 153494 181292
rect 154718 181280 154724 181292
rect 154776 181280 154782 181332
rect 245338 181280 245344 181332
rect 245396 181320 245402 181332
rect 245798 181320 245804 181332
rect 245396 181292 245804 181320
rect 245396 181280 245402 181292
rect 245798 181280 245804 181292
rect 245856 181280 245862 181332
rect 252054 181280 252060 181332
rect 252112 181320 252118 181332
rect 257574 181320 257580 181332
rect 252112 181292 257580 181320
rect 252112 181280 252118 181292
rect 257574 181280 257580 181292
rect 257632 181280 257638 181332
rect 337614 181280 337620 181332
rect 337672 181320 337678 181332
rect 341110 181320 341116 181332
rect 337672 181292 341116 181320
rect 337672 181280 337678 181292
rect 341110 181280 341116 181292
rect 341168 181280 341174 181332
rect 345158 181280 345164 181332
rect 345216 181320 345222 181332
rect 359786 181320 359792 181332
rect 345216 181292 359792 181320
rect 345216 181280 345222 181292
rect 359786 181280 359792 181292
rect 359844 181280 359850 181332
rect 361166 181280 361172 181332
rect 361224 181320 361230 181332
rect 412870 181320 412876 181332
rect 361224 181292 412876 181320
rect 361224 181280 361230 181292
rect 412870 181280 412876 181292
rect 412928 181280 412934 181332
rect 346170 181252 346176 181264
rect 336804 181224 346176 181252
rect 149198 181144 149204 181196
rect 149256 181184 149262 181196
rect 158214 181184 158220 181196
rect 149256 181156 158220 181184
rect 149256 181144 149262 181156
rect 158214 181144 158220 181156
rect 158272 181144 158278 181196
rect 149750 181076 149756 181128
rect 149808 181116 149814 181128
rect 160330 181116 160336 181128
rect 149808 181088 160336 181116
rect 149808 181076 149814 181088
rect 160330 181076 160336 181088
rect 160388 181076 160394 181128
rect 150578 181008 150584 181060
rect 150636 181048 150642 181060
rect 162722 181048 162728 181060
rect 150636 181020 162728 181048
rect 150636 181008 150642 181020
rect 162722 181008 162728 181020
rect 162780 181008 162786 181060
rect 243498 181008 243504 181060
rect 243556 181048 243562 181060
rect 252790 181048 252796 181060
rect 243556 181020 252796 181048
rect 243556 181008 243562 181020
rect 252790 181008 252796 181020
rect 252848 181008 252854 181060
rect 151958 180940 151964 180992
rect 152016 180980 152022 180992
rect 163274 180980 163280 180992
rect 152016 180952 163280 180980
rect 152016 180940 152022 180952
rect 163274 180940 163280 180952
rect 163332 180940 163338 180992
rect 244050 180940 244056 180992
rect 244108 180980 244114 180992
rect 254170 180980 254176 180992
rect 244108 180952 254176 180980
rect 244108 180940 244114 180952
rect 254170 180940 254176 180952
rect 254228 180940 254234 180992
rect 334118 180940 334124 180992
rect 334176 180980 334182 180992
rect 336804 180980 336832 181224
rect 346170 181212 346176 181224
rect 346228 181212 346234 181264
rect 370734 181212 370740 181264
rect 370792 181252 370798 181264
rect 410202 181252 410208 181264
rect 370792 181224 410208 181252
rect 370792 181212 370798 181224
rect 410202 181212 410208 181224
rect 410260 181212 410266 181264
rect 338258 181144 338264 181196
rect 338316 181184 338322 181196
rect 341846 181184 341852 181196
rect 338316 181156 341852 181184
rect 338316 181144 338322 181156
rect 341846 181144 341852 181156
rect 341904 181144 341910 181196
rect 340098 181076 340104 181128
rect 340156 181116 340162 181128
rect 343870 181116 343876 181128
rect 340156 181088 343876 181116
rect 340156 181076 340162 181088
rect 343870 181076 343876 181088
rect 343928 181076 343934 181128
rect 336878 181008 336884 181060
rect 336936 181048 336942 181060
rect 348746 181048 348752 181060
rect 336936 181020 348752 181048
rect 336936 181008 336942 181020
rect 348746 181008 348752 181020
rect 348804 181008 348810 181060
rect 334176 180952 336832 180980
rect 334176 180940 334182 180952
rect 339638 180940 339644 180992
rect 339696 180980 339702 180992
rect 351230 180980 351236 180992
rect 339696 180952 351236 180980
rect 339696 180940 339702 180952
rect 351230 180940 351236 180952
rect 351288 180940 351294 180992
rect 34658 180872 34664 180924
rect 34716 180912 34722 180924
rect 46986 180912 46992 180924
rect 34716 180884 46992 180912
rect 34716 180872 34722 180884
rect 46986 180872 46992 180884
rect 47044 180872 47050 180924
rect 149198 180872 149204 180924
rect 149256 180912 149262 180924
rect 162078 180912 162084 180924
rect 149256 180884 162084 180912
rect 149256 180872 149262 180884
rect 162078 180872 162084 180884
rect 162136 180872 162142 180924
rect 243038 180872 243044 180924
rect 243096 180912 243102 180924
rect 255734 180912 255740 180924
rect 243096 180884 255740 180912
rect 243096 180872 243102 180884
rect 255734 180872 255740 180884
rect 255792 180872 255798 180924
rect 31806 180804 31812 180856
rect 31864 180844 31870 180856
rect 45790 180844 45796 180856
rect 31864 180816 45796 180844
rect 31864 180804 31870 180816
rect 45790 180804 45796 180816
rect 45848 180804 45854 180856
rect 147818 180804 147824 180856
rect 147876 180844 147882 180856
rect 161434 180844 161440 180856
rect 147876 180816 161440 180844
rect 147876 180804 147882 180816
rect 161434 180804 161440 180816
rect 161492 180804 161498 180856
rect 240278 180804 240284 180856
rect 240336 180844 240342 180856
rect 254538 180844 254544 180856
rect 240336 180816 254544 180844
rect 240336 180804 240342 180816
rect 254538 180804 254544 180816
rect 254596 180804 254602 180856
rect 341018 180804 341024 180856
rect 341076 180844 341082 180856
rect 348013 180847 348071 180853
rect 348013 180844 348025 180847
rect 341076 180816 348025 180844
rect 341076 180804 341082 180816
rect 348013 180813 348025 180816
rect 348059 180813 348071 180847
rect 348013 180807 348071 180813
rect 29506 180736 29512 180788
rect 29564 180776 29570 180788
rect 46618 180776 46624 180788
rect 29564 180748 46624 180776
rect 29564 180736 29570 180748
rect 46618 180736 46624 180748
rect 46676 180736 46682 180788
rect 145058 180736 145064 180788
rect 145116 180776 145122 180788
rect 160238 180776 160244 180788
rect 145116 180748 160244 180776
rect 145116 180736 145122 180748
rect 160238 180736 160244 180748
rect 160296 180736 160302 180788
rect 241658 180736 241664 180788
rect 241716 180776 241722 180788
rect 255090 180776 255096 180788
rect 241716 180748 255096 180776
rect 241716 180736 241722 180748
rect 255090 180736 255096 180748
rect 255148 180736 255154 180788
rect 335406 180736 335412 180788
rect 335464 180776 335470 180788
rect 346998 180776 347004 180788
rect 335464 180748 347004 180776
rect 335464 180736 335470 180748
rect 346998 180736 347004 180748
rect 347056 180736 347062 180788
rect 26930 180668 26936 180720
rect 26988 180708 26994 180720
rect 46526 180708 46532 180720
rect 26988 180680 46532 180708
rect 26988 180668 26994 180680
rect 46526 180668 46532 180680
rect 46584 180668 46590 180720
rect 238898 180668 238904 180720
rect 238956 180708 238962 180720
rect 254262 180708 254268 180720
rect 238956 180680 254268 180708
rect 238956 180668 238962 180680
rect 254262 180668 254268 180680
rect 254320 180668 254326 180720
rect 332738 180668 332744 180720
rect 332796 180708 332802 180720
rect 345342 180708 345348 180720
rect 332796 180680 345348 180708
rect 332796 180668 332802 180680
rect 345342 180668 345348 180680
rect 345400 180668 345406 180720
rect 24170 180600 24176 180652
rect 24228 180640 24234 180652
rect 46434 180640 46440 180652
rect 24228 180612 46440 180640
rect 24228 180600 24234 180612
rect 46434 180600 46440 180612
rect 46492 180600 46498 180652
rect 57014 180600 57020 180652
rect 57072 180640 57078 180652
rect 68054 180640 68060 180652
rect 57072 180612 68060 180640
rect 57072 180600 57078 180612
rect 68054 180600 68060 180612
rect 68112 180600 68118 180652
rect 146438 180600 146444 180652
rect 146496 180640 146502 180652
rect 160882 180640 160888 180652
rect 146496 180612 160888 180640
rect 146496 180600 146502 180612
rect 160882 180600 160888 180612
rect 160940 180600 160946 180652
rect 237518 180600 237524 180652
rect 237576 180640 237582 180652
rect 253434 180640 253440 180652
rect 237576 180612 253440 180640
rect 237576 180600 237582 180612
rect 253434 180600 253440 180612
rect 253492 180600 253498 180652
rect 335498 180600 335504 180652
rect 335556 180640 335562 180652
rect 348010 180640 348016 180652
rect 335556 180612 348016 180640
rect 335556 180600 335562 180612
rect 348010 180600 348016 180612
rect 348068 180600 348074 180652
rect 143678 180532 143684 180584
rect 143736 180572 143742 180584
rect 159594 180572 159600 180584
rect 143736 180544 159600 180572
rect 143736 180532 143742 180544
rect 159594 180532 159600 180544
rect 159652 180532 159658 180584
rect 338258 180532 338264 180584
rect 338316 180572 338322 180584
rect 349574 180572 349580 180584
rect 338316 180544 349580 180572
rect 338316 180532 338322 180544
rect 349574 180532 349580 180544
rect 349632 180532 349638 180584
rect 62350 180464 62356 180516
rect 62408 180504 62414 180516
rect 63638 180504 63644 180516
rect 62408 180476 63644 180504
rect 62408 180464 62414 180476
rect 63638 180464 63644 180476
rect 63696 180464 63702 180516
rect 68514 180464 68520 180516
rect 68572 180504 68578 180516
rect 69434 180504 69440 180516
rect 68572 180476 69440 180504
rect 68572 180464 68578 180476
rect 69434 180464 69440 180476
rect 69492 180464 69498 180516
rect 247730 180464 247736 180516
rect 247788 180504 247794 180516
rect 248558 180504 248564 180516
rect 247788 180476 248564 180504
rect 247788 180464 247794 180476
rect 248558 180464 248564 180476
rect 248616 180464 248622 180516
rect 339270 180464 339276 180516
rect 339328 180504 339334 180516
rect 341754 180504 341760 180516
rect 339328 180476 341760 180504
rect 339328 180464 339334 180476
rect 341754 180464 341760 180476
rect 341812 180464 341818 180516
rect 340926 180396 340932 180448
rect 340984 180436 340990 180448
rect 344606 180436 344612 180448
rect 340984 180408 344612 180436
rect 340984 180396 340990 180408
rect 344606 180396 344612 180408
rect 344664 180396 344670 180448
rect 246534 180328 246540 180380
rect 246592 180368 246598 180380
rect 247178 180368 247184 180380
rect 246592 180340 247184 180368
rect 246592 180328 246598 180340
rect 247178 180328 247184 180340
rect 247236 180328 247242 180380
rect 343502 180124 343508 180176
rect 343560 180164 343566 180176
rect 348010 180164 348016 180176
rect 343560 180136 348016 180164
rect 343560 180124 343566 180136
rect 348010 180124 348016 180136
rect 348068 180124 348074 180176
rect 341662 180056 341668 180108
rect 341720 180096 341726 180108
rect 344698 180096 344704 180108
rect 341720 180068 344704 180096
rect 341720 180056 341726 180068
rect 344698 180056 344704 180068
rect 344756 180056 344762 180108
rect 344330 179988 344336 180040
rect 344388 180028 344394 180040
rect 347274 180028 347280 180040
rect 344388 180000 347280 180028
rect 344388 179988 344394 180000
rect 347274 179988 347280 180000
rect 347332 179988 347338 180040
rect 254814 179920 254820 179972
rect 254872 179960 254878 179972
rect 258402 179960 258408 179972
rect 254872 179932 258408 179960
rect 254872 179920 254878 179932
rect 258402 179920 258408 179932
rect 258460 179920 258466 179972
rect 342398 179920 342404 179972
rect 342456 179960 342462 179972
rect 344514 179960 344520 179972
rect 342456 179932 344520 179960
rect 342456 179920 342462 179932
rect 344514 179920 344520 179932
rect 344572 179920 344578 179972
rect 368986 179920 368992 179972
rect 369044 179960 369050 179972
rect 369354 179960 369360 179972
rect 369044 179932 369360 179960
rect 369044 179920 369050 179932
rect 369354 179920 369360 179932
rect 369412 179920 369418 179972
rect 369538 179920 369544 179972
rect 369596 179960 369602 179972
rect 369906 179960 369912 179972
rect 369596 179932 369912 179960
rect 369596 179920 369602 179932
rect 369906 179920 369912 179932
rect 369964 179920 369970 179972
rect 324550 179852 324556 179904
rect 324608 179892 324614 179904
rect 326574 179892 326580 179904
rect 324608 179864 326580 179892
rect 324608 179852 324614 179864
rect 326574 179852 326580 179864
rect 326632 179852 326638 179904
rect 230986 179716 230992 179768
rect 231044 179756 231050 179768
rect 232734 179756 232740 179768
rect 231044 179728 232740 179756
rect 231044 179716 231050 179728
rect 232734 179716 232740 179728
rect 232792 179716 232798 179768
rect 427590 178492 427596 178544
rect 427648 178532 427654 178544
rect 429890 178532 429896 178544
rect 427648 178504 429896 178532
rect 427648 178492 427654 178504
rect 429890 178492 429896 178504
rect 429948 178492 429954 178544
rect 368526 177880 368532 177932
rect 368584 177920 368590 177932
rect 368710 177920 368716 177932
rect 368584 177892 368716 177920
rect 368584 177880 368590 177892
rect 368710 177880 368716 177892
rect 368768 177880 368774 177932
rect 358314 175908 358320 175960
rect 358372 175908 358378 175960
rect 358332 175824 358360 175908
rect 88386 175772 88392 175824
rect 88444 175812 88450 175824
rect 178270 175812 178276 175824
rect 88444 175784 178276 175812
rect 88444 175772 88450 175784
rect 178270 175772 178276 175784
rect 178328 175772 178334 175824
rect 182410 175772 182416 175824
rect 182468 175812 182474 175824
rect 182870 175812 182876 175824
rect 182468 175784 182876 175812
rect 182468 175772 182474 175784
rect 182870 175772 182876 175784
rect 182928 175812 182934 175824
rect 276434 175812 276440 175824
rect 182928 175784 276440 175812
rect 182928 175772 182934 175784
rect 276434 175772 276440 175784
rect 276492 175772 276498 175824
rect 358314 175772 358320 175824
rect 358372 175772 358378 175824
rect 95470 175704 95476 175756
rect 95528 175744 95534 175756
rect 170634 175744 170640 175756
rect 95528 175716 170640 175744
rect 95528 175704 95534 175716
rect 170634 175704 170640 175716
rect 170692 175744 170698 175756
rect 189494 175744 189500 175756
rect 170692 175716 189500 175744
rect 170692 175704 170698 175716
rect 189494 175704 189500 175716
rect 189552 175744 189558 175756
rect 283518 175744 283524 175756
rect 189552 175716 283524 175744
rect 189552 175704 189558 175716
rect 283518 175704 283524 175716
rect 283576 175704 283582 175756
rect 196670 175636 196676 175688
rect 196728 175676 196734 175688
rect 268614 175676 268620 175688
rect 196728 175648 268620 175676
rect 196728 175636 196734 175648
rect 268614 175636 268620 175648
rect 268672 175676 268678 175688
rect 290694 175676 290700 175688
rect 268672 175648 290700 175676
rect 268672 175636 268678 175648
rect 290694 175636 290700 175648
rect 290752 175636 290758 175688
rect 96758 175160 96764 175212
rect 96816 175200 96822 175212
rect 109730 175200 109736 175212
rect 96816 175172 109736 175200
rect 96816 175160 96822 175172
rect 109730 175160 109736 175172
rect 109788 175160 109794 175212
rect 190598 175160 190604 175212
rect 190656 175200 190662 175212
rect 203754 175200 203760 175212
rect 190656 175172 203760 175200
rect 190656 175160 190662 175172
rect 203754 175160 203760 175172
rect 203812 175160 203818 175212
rect 102646 175092 102652 175144
rect 102704 175132 102710 175144
rect 176154 175132 176160 175144
rect 102704 175104 176160 175132
rect 102704 175092 102710 175104
rect 176154 175092 176160 175104
rect 176212 175132 176218 175144
rect 196670 175132 196676 175144
rect 176212 175104 196676 175132
rect 176212 175092 176218 175104
rect 196670 175092 196676 175104
rect 196728 175092 196734 175144
rect 285818 175092 285824 175144
rect 285876 175132 285882 175144
rect 297778 175132 297784 175144
rect 285876 175104 297784 175132
rect 285876 175092 285882 175104
rect 297778 175092 297784 175104
rect 297836 175092 297842 175144
rect 124358 174412 124364 174464
rect 124416 174452 124422 174464
rect 131166 174452 131172 174464
rect 124416 174424 131172 174452
rect 124416 174412 124422 174424
rect 131166 174412 131172 174424
rect 131224 174412 131230 174464
rect 60694 172984 60700 173036
rect 60752 173024 60758 173036
rect 65938 173024 65944 173036
rect 60752 172996 65944 173024
rect 60752 172984 60758 172996
rect 65938 172984 65944 172996
rect 65996 172984 66002 173036
rect 153154 172984 153160 173036
rect 153212 173024 153218 173036
rect 153338 173024 153344 173036
rect 153212 172996 153344 173024
rect 153212 172984 153218 172996
rect 153338 172984 153344 172996
rect 153396 172984 153402 173036
rect 158214 172984 158220 173036
rect 158272 173024 158278 173036
rect 158950 173024 158956 173036
rect 158272 172996 158956 173024
rect 158272 172984 158278 172996
rect 158950 172984 158956 172996
rect 159008 172984 159014 173036
rect 249018 172984 249024 173036
rect 249076 173024 249082 173036
rect 254814 173024 254820 173036
rect 249076 172996 254820 173024
rect 249076 172984 249082 172996
rect 254814 172984 254820 172996
rect 254872 172984 254878 173036
rect 333382 172984 333388 173036
rect 333440 173024 333446 173036
rect 334118 173024 334124 173036
rect 333440 172996 334124 173024
rect 333440 172984 333446 172996
rect 334118 172984 334124 172996
rect 334176 172984 334182 173036
rect 341846 172984 341852 173036
rect 341904 173024 341910 173036
rect 342674 173024 342680 173036
rect 341904 172996 342680 173024
rect 341904 172984 341910 172996
rect 342674 172984 342680 172996
rect 342732 172984 342738 173036
rect 347274 172984 347280 173036
rect 347332 173024 347338 173036
rect 349942 173024 349948 173036
rect 347332 172996 349948 173024
rect 347332 172984 347338 172996
rect 349942 172984 349948 172996
rect 350000 172984 350006 173036
rect 64834 172916 64840 172968
rect 64892 172956 64898 172968
rect 68514 172956 68520 172968
rect 64892 172928 68520 172956
rect 64892 172916 64898 172928
rect 68514 172916 68520 172928
rect 68572 172916 68578 172968
rect 154534 172916 154540 172968
rect 154592 172956 154598 172968
rect 164654 172956 164660 172968
rect 154592 172928 164660 172956
rect 154592 172916 154598 172928
rect 164654 172916 164660 172928
rect 164712 172916 164718 172968
rect 246258 172916 246264 172968
rect 246316 172956 246322 172968
rect 257298 172956 257304 172968
rect 246316 172928 257304 172956
rect 246316 172916 246322 172928
rect 257298 172916 257304 172928
rect 257356 172916 257362 172968
rect 341754 172916 341760 172968
rect 341812 172956 341818 172968
rect 343778 172956 343784 172968
rect 341812 172928 343784 172956
rect 341812 172916 341818 172928
rect 343778 172916 343784 172928
rect 343836 172916 343842 172968
rect 59682 172848 59688 172900
rect 59740 172888 59746 172900
rect 65018 172888 65024 172900
rect 59740 172860 65024 172888
rect 59740 172848 59746 172860
rect 65018 172848 65024 172860
rect 65076 172848 65082 172900
rect 153338 172848 153344 172900
rect 153396 172888 153402 172900
rect 163918 172888 163924 172900
rect 153396 172860 163924 172888
rect 153396 172848 153402 172860
rect 163918 172848 163924 172860
rect 163976 172848 163982 172900
rect 244878 172848 244884 172900
rect 244936 172888 244942 172900
rect 256746 172888 256752 172900
rect 244936 172860 256752 172888
rect 244936 172848 244942 172860
rect 256746 172848 256752 172860
rect 256804 172848 256810 172900
rect 63638 172780 63644 172832
rect 63696 172820 63702 172832
rect 75230 172820 75236 172832
rect 63696 172792 75236 172820
rect 63696 172780 63702 172792
rect 75230 172780 75236 172792
rect 75288 172780 75294 172832
rect 150302 172780 150308 172832
rect 150360 172820 150366 172832
rect 161710 172820 161716 172832
rect 150360 172792 161716 172820
rect 150360 172780 150366 172792
rect 161710 172780 161716 172792
rect 161768 172780 161774 172832
rect 245798 172780 245804 172832
rect 245856 172820 245862 172832
rect 256930 172820 256936 172832
rect 245856 172792 256936 172820
rect 245856 172780 245862 172792
rect 256930 172780 256936 172792
rect 256988 172780 256994 172832
rect 60878 172712 60884 172764
rect 60936 172752 60942 172764
rect 72102 172752 72108 172764
rect 60936 172724 72108 172752
rect 60936 172712 60942 172724
rect 72102 172712 72108 172724
rect 72160 172712 72166 172764
rect 151866 172712 151872 172764
rect 151924 172752 151930 172764
rect 163090 172752 163096 172764
rect 151924 172724 163096 172752
rect 151924 172712 151930 172724
rect 163090 172712 163096 172724
rect 163148 172712 163154 172764
rect 244418 172712 244424 172764
rect 244476 172752 244482 172764
rect 255550 172752 255556 172764
rect 244476 172724 255556 172752
rect 244476 172712 244482 172724
rect 255550 172712 255556 172724
rect 255608 172712 255614 172764
rect 62258 172644 62264 172696
rect 62316 172684 62322 172696
rect 74218 172684 74224 172696
rect 62316 172656 74224 172684
rect 62316 172644 62322 172656
rect 74218 172644 74224 172656
rect 74276 172644 74282 172696
rect 143034 172644 143040 172696
rect 143092 172684 143098 172696
rect 155730 172684 155736 172696
rect 143092 172656 155736 172684
rect 143092 172644 143098 172656
rect 155730 172644 155736 172656
rect 155788 172644 155794 172696
rect 157846 172644 157852 172696
rect 157904 172684 157910 172696
rect 165114 172684 165120 172696
rect 157904 172656 165120 172684
rect 157904 172644 157910 172656
rect 165114 172644 165120 172656
rect 165172 172644 165178 172696
rect 247178 172644 247184 172696
rect 247236 172684 247242 172696
rect 259690 172684 259696 172696
rect 247236 172656 259696 172684
rect 247236 172644 247242 172656
rect 259690 172644 259696 172656
rect 259748 172644 259754 172696
rect 59498 172576 59504 172628
rect 59556 172616 59562 172628
rect 71090 172616 71096 172628
rect 59556 172588 71096 172616
rect 59556 172576 59562 172588
rect 71090 172576 71096 172588
rect 71148 172576 71154 172628
rect 153246 172576 153252 172628
rect 153304 172616 153310 172628
rect 165850 172616 165856 172628
rect 153304 172588 165856 172616
rect 153304 172576 153310 172588
rect 165850 172576 165856 172588
rect 165908 172576 165914 172628
rect 246810 172576 246816 172628
rect 246868 172616 246874 172628
rect 252241 172619 252299 172625
rect 252241 172616 252253 172619
rect 246868 172588 252253 172616
rect 246868 172576 246874 172588
rect 252241 172585 252253 172588
rect 252287 172585 252299 172619
rect 252241 172579 252299 172585
rect 252333 172619 252391 172625
rect 252333 172585 252345 172619
rect 252379 172616 252391 172619
rect 258310 172616 258316 172628
rect 252379 172588 258316 172616
rect 252379 172585 252391 172588
rect 252333 172579 252391 172585
rect 258310 172576 258316 172588
rect 258368 172576 258374 172628
rect 354910 172576 354916 172628
rect 354968 172616 354974 172628
rect 355830 172616 355836 172628
rect 354968 172588 355836 172616
rect 354968 172576 354974 172588
rect 355830 172576 355836 172588
rect 355888 172576 355894 172628
rect 58026 172508 58032 172560
rect 58084 172548 58090 172560
rect 70078 172548 70084 172560
rect 58084 172520 70084 172548
rect 58084 172508 58090 172520
rect 70078 172508 70084 172520
rect 70136 172508 70142 172560
rect 151682 172508 151688 172560
rect 151740 172548 151746 172560
rect 164470 172548 164476 172560
rect 151740 172520 164476 172548
rect 151740 172508 151746 172520
rect 164470 172508 164476 172520
rect 164528 172508 164534 172560
rect 236874 172508 236880 172560
rect 236932 172548 236938 172560
rect 250030 172548 250036 172560
rect 236932 172520 250036 172548
rect 236932 172508 236938 172520
rect 250030 172508 250036 172520
rect 250088 172508 250094 172560
rect 55358 172440 55364 172492
rect 55416 172480 55422 172492
rect 66950 172480 66956 172492
rect 55416 172452 66956 172480
rect 55416 172440 55422 172452
rect 66950 172440 66956 172452
rect 67008 172440 67014 172492
rect 154718 172440 154724 172492
rect 154776 172480 154782 172492
rect 168610 172480 168616 172492
rect 154776 172452 168616 172480
rect 154776 172440 154782 172452
rect 168610 172440 168616 172452
rect 168668 172440 168674 172492
rect 247638 172440 247644 172492
rect 247696 172480 247702 172492
rect 252054 172480 252060 172492
rect 247696 172452 252060 172480
rect 247696 172440 247702 172452
rect 252054 172440 252060 172452
rect 252112 172440 252118 172492
rect 262450 172480 262456 172492
rect 252164 172452 262456 172480
rect 56738 172372 56744 172424
rect 56796 172412 56802 172424
rect 67962 172412 67968 172424
rect 56796 172384 67968 172412
rect 56796 172372 56802 172384
rect 67962 172372 67968 172384
rect 68020 172372 68026 172424
rect 153154 172372 153160 172424
rect 153212 172412 153218 172424
rect 167230 172412 167236 172424
rect 153212 172384 167236 172412
rect 153212 172372 153218 172384
rect 167230 172372 167236 172384
rect 167288 172372 167294 172424
rect 248558 172372 248564 172424
rect 248616 172412 248622 172424
rect 252164 172412 252192 172452
rect 262450 172440 262456 172452
rect 262508 172440 262514 172492
rect 248616 172384 252192 172412
rect 252241 172415 252299 172421
rect 248616 172372 248622 172384
rect 252241 172381 252253 172415
rect 252287 172412 252299 172415
rect 261162 172412 261168 172424
rect 252287 172384 261168 172412
rect 252287 172381 252299 172384
rect 252241 172375 252299 172381
rect 261162 172372 261168 172384
rect 261220 172372 261226 172424
rect 60602 172304 60608 172356
rect 60660 172344 60666 172356
rect 73114 172344 73120 172356
rect 60660 172316 73120 172344
rect 60660 172304 60666 172316
rect 73114 172304 73120 172316
rect 73172 172304 73178 172356
rect 154626 172304 154632 172356
rect 154684 172344 154690 172356
rect 169990 172344 169996 172356
rect 154684 172316 169996 172344
rect 154684 172304 154690 172316
rect 169990 172304 169996 172316
rect 170048 172304 170054 172356
rect 248006 172304 248012 172356
rect 248064 172344 248070 172356
rect 263830 172344 263836 172356
rect 248064 172316 263836 172344
rect 248064 172304 248070 172316
rect 263830 172304 263836 172316
rect 263888 172304 263894 172356
rect 338534 172304 338540 172356
rect 338592 172344 338598 172356
rect 350678 172344 350684 172356
rect 338592 172316 350684 172344
rect 338592 172304 338598 172316
rect 350678 172304 350684 172316
rect 350736 172304 350742 172356
rect 63822 172236 63828 172288
rect 63880 172276 63886 172288
rect 68606 172276 68612 172288
rect 63880 172248 68612 172276
rect 63880 172236 63886 172248
rect 68606 172236 68612 172248
rect 68664 172236 68670 172288
rect 245522 172236 245528 172288
rect 245580 172276 245586 172288
rect 252333 172279 252391 172285
rect 252333 172276 252345 172279
rect 245580 172248 252345 172276
rect 245580 172236 245586 172248
rect 252333 172245 252345 172248
rect 252379 172245 252391 172279
rect 252333 172239 252391 172245
rect 58670 172032 58676 172084
rect 58728 172072 58734 172084
rect 62994 172072 63000 172084
rect 58728 172044 63000 172072
rect 58728 172032 58734 172044
rect 62994 172032 63000 172044
rect 63052 172032 63058 172084
rect 65938 172032 65944 172084
rect 65996 172072 66002 172084
rect 70446 172072 70452 172084
rect 65996 172044 70452 172072
rect 65996 172032 66002 172044
rect 70446 172032 70452 172044
rect 70504 172032 70510 172084
rect 334394 172032 334400 172084
rect 334452 172072 334458 172084
rect 335406 172072 335412 172084
rect 334452 172044 335412 172072
rect 334452 172032 334458 172044
rect 335406 172032 335412 172044
rect 335464 172032 335470 172084
rect 57658 171896 57664 171948
rect 57716 171936 57722 171948
rect 63270 171936 63276 171948
rect 57716 171908 63276 171936
rect 57716 171896 57722 171908
rect 63270 171896 63276 171908
rect 63328 171896 63334 171948
rect 62810 171828 62816 171880
rect 62868 171868 62874 171880
rect 67686 171868 67692 171880
rect 62868 171840 67692 171868
rect 62868 171828 62874 171840
rect 67686 171828 67692 171840
rect 67744 171828 67750 171880
rect 344514 171828 344520 171880
rect 344572 171868 344578 171880
rect 347918 171868 347924 171880
rect 344572 171840 347924 171868
rect 344572 171828 344578 171840
rect 347918 171828 347924 171840
rect 347976 171828 347982 171880
rect 344698 171760 344704 171812
rect 344756 171800 344762 171812
rect 346814 171800 346820 171812
rect 344756 171772 346820 171800
rect 344756 171760 344762 171772
rect 346814 171760 346820 171772
rect 346872 171760 346878 171812
rect 61798 171692 61804 171744
rect 61856 171732 61862 171744
rect 65754 171732 65760 171744
rect 61856 171704 65760 171732
rect 61856 171692 61862 171704
rect 65754 171692 65760 171704
rect 65812 171692 65818 171744
rect 251870 171692 251876 171744
rect 251928 171732 251934 171744
rect 258954 171732 258960 171744
rect 251928 171704 258960 171732
rect 251928 171692 251934 171704
rect 258954 171692 258960 171704
rect 259012 171692 259018 171744
rect 344606 171692 344612 171744
rect 344664 171732 344670 171744
rect 345802 171732 345808 171744
rect 344664 171704 345808 171732
rect 344664 171692 344670 171704
rect 345802 171692 345808 171704
rect 345860 171692 345866 171744
rect 358406 171556 358412 171608
rect 358464 171596 358470 171608
rect 358590 171596 358596 171608
rect 358464 171568 358596 171596
rect 358464 171556 358470 171568
rect 358590 171556 358596 171568
rect 358648 171556 358654 171608
rect 79738 170196 79744 170248
rect 79796 170236 79802 170248
rect 123990 170236 123996 170248
rect 79796 170208 123996 170236
rect 79796 170196 79802 170208
rect 123990 170196 123996 170208
rect 124048 170196 124054 170248
rect 312038 170196 312044 170248
rect 312096 170236 312102 170248
rect 328414 170236 328420 170248
rect 312096 170208 328420 170236
rect 312096 170196 312102 170208
rect 328414 170196 328420 170208
rect 328472 170196 328478 170248
rect 123990 169516 123996 169568
rect 124048 169556 124054 169568
rect 140274 169556 140280 169568
rect 124048 169528 140280 169556
rect 124048 169516 124054 169528
rect 140274 169516 140280 169528
rect 140332 169516 140338 169568
rect 267234 169516 267240 169568
rect 267292 169556 267298 169568
rect 312038 169556 312044 169568
rect 267292 169528 312044 169556
rect 267292 169516 267298 169528
rect 312038 169516 312044 169528
rect 312096 169516 312102 169568
rect 71642 169420 71648 169432
rect 71603 169392 71648 169420
rect 71642 169380 71648 169392
rect 71700 169380 71706 169432
rect 132178 168904 132184 168956
rect 132236 168944 132242 168956
rect 140550 168944 140556 168956
rect 132236 168916 140556 168944
rect 132236 168904 132242 168916
rect 140550 168904 140556 168916
rect 140608 168904 140614 168956
rect 225834 168904 225840 168956
rect 225892 168944 225898 168956
rect 233470 168944 233476 168956
rect 225892 168916 233476 168944
rect 225892 168904 225898 168916
rect 233470 168904 233476 168916
rect 233528 168904 233534 168956
rect 46986 168836 46992 168888
rect 47044 168876 47050 168888
rect 49194 168876 49200 168888
rect 47044 168848 49200 168876
rect 47044 168836 47050 168848
rect 49194 168836 49200 168848
rect 49252 168876 49258 168888
rect 71645 168879 71703 168885
rect 71645 168876 71657 168879
rect 49252 168848 71657 168876
rect 49252 168836 49258 168848
rect 71645 168845 71657 168848
rect 71691 168845 71703 168879
rect 71645 168839 71703 168845
rect 359694 168836 359700 168888
rect 359752 168876 359758 168888
rect 423634 168876 423640 168888
rect 359752 168848 423640 168876
rect 359752 168836 359758 168848
rect 423634 168836 423640 168848
rect 423692 168836 423698 168888
rect 222154 168564 222160 168616
rect 222212 168604 222218 168616
rect 369262 168604 369268 168616
rect 222212 168576 369268 168604
rect 222212 168564 222218 168576
rect 369262 168564 369268 168576
rect 369320 168564 369326 168616
rect 128130 168496 128136 168548
rect 128188 168536 128194 168548
rect 368986 168536 368992 168548
rect 128188 168508 368992 168536
rect 128188 168496 128194 168508
rect 368986 168496 368992 168508
rect 369044 168496 369050 168548
rect 368710 168156 368716 168208
rect 368768 168196 368774 168208
rect 368986 168196 368992 168208
rect 368768 168168 368992 168196
rect 368768 168156 368774 168168
rect 368986 168156 368992 168168
rect 369044 168156 369050 168208
rect 77254 167544 77260 167596
rect 77312 167584 77318 167596
rect 87190 167584 87196 167596
rect 77312 167556 87196 167584
rect 77312 167544 77318 167556
rect 87190 167544 87196 167556
rect 87248 167544 87254 167596
rect 132270 167544 132276 167596
rect 132328 167584 132334 167596
rect 140550 167584 140556 167596
rect 132328 167556 140556 167584
rect 132328 167544 132334 167556
rect 140550 167544 140556 167556
rect 140608 167544 140614 167596
rect 226018 167544 226024 167596
rect 226076 167584 226082 167596
rect 233470 167584 233476 167596
rect 226076 167556 233476 167584
rect 226076 167544 226082 167556
rect 233470 167544 233476 167556
rect 233528 167544 233534 167596
rect 203846 166932 203852 166984
rect 203904 166972 203910 166984
rect 210930 166972 210936 166984
rect 203904 166944 210936 166972
rect 203904 166932 203910 166944
rect 210930 166932 210936 166944
rect 210988 166932 210994 166984
rect 110190 166796 110196 166848
rect 110248 166836 110254 166848
rect 116906 166836 116912 166848
rect 110248 166808 116912 166836
rect 110248 166796 110254 166808
rect 116906 166796 116912 166808
rect 116964 166796 116970 166848
rect 217186 166796 217192 166848
rect 217244 166836 217250 166848
rect 225190 166836 225196 166848
rect 217244 166808 225196 166836
rect 217244 166796 217250 166808
rect 225190 166796 225196 166808
rect 225248 166796 225254 166848
rect 297870 166796 297876 166848
rect 297928 166836 297934 166848
rect 304954 166836 304960 166848
rect 297928 166808 304960 166836
rect 297928 166796 297934 166808
rect 304954 166796 304960 166808
rect 305012 166796 305018 166848
rect 311210 166796 311216 166848
rect 311268 166836 311274 166848
rect 319214 166836 319220 166848
rect 311268 166808 319220 166836
rect 311268 166796 311274 166808
rect 319214 166796 319220 166808
rect 319272 166796 319278 166848
rect 123530 166320 123536 166372
rect 123588 166360 123594 166372
rect 124358 166360 124364 166372
rect 123588 166332 124364 166360
rect 123588 166320 123594 166332
rect 124358 166320 124364 166332
rect 124416 166320 124422 166372
rect 284530 166252 284536 166304
rect 284588 166292 284594 166304
rect 285818 166292 285824 166304
rect 284588 166264 285824 166292
rect 284588 166252 284594 166264
rect 285818 166252 285824 166264
rect 285876 166252 285882 166304
rect 77254 166184 77260 166236
rect 77312 166224 77318 166236
rect 85718 166224 85724 166236
rect 77312 166196 85724 166224
rect 77312 166184 77318 166196
rect 85718 166184 85724 166196
rect 85776 166184 85782 166236
rect 132086 166184 132092 166236
rect 132144 166224 132150 166236
rect 140550 166224 140556 166236
rect 132144 166196 140556 166224
rect 132144 166184 132150 166196
rect 140550 166184 140556 166196
rect 140608 166184 140614 166236
rect 225926 166184 225932 166236
rect 225984 166224 225990 166236
rect 233470 166224 233476 166236
rect 225984 166196 233476 166224
rect 225984 166184 225990 166196
rect 233470 166184 233476 166196
rect 233528 166184 233534 166236
rect 324550 166184 324556 166236
rect 324608 166224 324614 166236
rect 328414 166224 328420 166236
rect 324608 166196 328420 166224
rect 324608 166184 324614 166196
rect 328414 166184 328420 166196
rect 328472 166184 328478 166236
rect 361258 165436 361264 165488
rect 361316 165476 361322 165488
rect 420874 165476 420880 165488
rect 361316 165448 420880 165476
rect 361316 165436 361322 165448
rect 420874 165436 420880 165448
rect 420932 165436 420938 165488
rect 79738 164824 79744 164876
rect 79796 164864 79802 164876
rect 85626 164864 85632 164876
rect 79796 164836 85632 164864
rect 79796 164824 79802 164836
rect 85626 164824 85632 164836
rect 85684 164824 85690 164876
rect 132546 164756 132552 164808
rect 132604 164796 132610 164808
rect 139630 164796 139636 164808
rect 132604 164768 139636 164796
rect 132604 164756 132610 164768
rect 139630 164756 139636 164768
rect 139688 164756 139694 164808
rect 225742 164756 225748 164808
rect 225800 164796 225806 164808
rect 233470 164796 233476 164808
rect 225800 164768 233476 164796
rect 225800 164756 225806 164768
rect 233470 164756 233476 164768
rect 233528 164756 233534 164808
rect 321790 164756 321796 164808
rect 321848 164796 321854 164808
rect 328506 164796 328512 164808
rect 321848 164768 328512 164796
rect 321848 164756 321854 164768
rect 328506 164756 328512 164768
rect 328564 164756 328570 164808
rect 132638 163464 132644 163516
rect 132696 163504 132702 163516
rect 139630 163504 139636 163516
rect 132696 163476 139636 163504
rect 132696 163464 132702 163476
rect 139630 163464 139636 163476
rect 139688 163464 139694 163516
rect 226294 163464 226300 163516
rect 226352 163504 226358 163516
rect 232826 163504 232832 163516
rect 226352 163476 232832 163504
rect 226352 163464 226358 163476
rect 232826 163464 232832 163476
rect 232884 163464 232890 163516
rect 321606 163464 321612 163516
rect 321664 163504 321670 163516
rect 327218 163504 327224 163516
rect 321664 163476 327224 163504
rect 321664 163464 321670 163476
rect 327218 163464 327224 163476
rect 327276 163464 327282 163516
rect 131350 163396 131356 163448
rect 131408 163436 131414 163448
rect 140550 163436 140556 163448
rect 131408 163408 140556 163436
rect 131408 163396 131414 163408
rect 140550 163396 140556 163408
rect 140608 163396 140614 163448
rect 179006 163396 179012 163448
rect 179064 163436 179070 163448
rect 182318 163436 182324 163448
rect 179064 163408 182324 163436
rect 179064 163396 179070 163408
rect 182318 163396 182324 163408
rect 182376 163396 182382 163448
rect 226110 163396 226116 163448
rect 226168 163436 226174 163448
rect 233470 163436 233476 163448
rect 226168 163408 233476 163436
rect 226168 163396 226174 163408
rect 233470 163396 233476 163408
rect 233528 163396 233534 163448
rect 85718 163328 85724 163380
rect 85776 163368 85782 163380
rect 87190 163368 87196 163380
rect 85776 163340 87196 163368
rect 85776 163328 85782 163340
rect 87190 163328 87196 163340
rect 87248 163328 87254 163380
rect 320962 163328 320968 163380
rect 321020 163368 321026 163380
rect 324550 163368 324556 163380
rect 321020 163340 324556 163368
rect 321020 163328 321026 163340
rect 324550 163328 324556 163340
rect 324608 163328 324614 163380
rect 358590 163368 358596 163380
rect 358551 163340 358596 163368
rect 358590 163328 358596 163340
rect 358648 163328 358654 163380
rect 12854 163192 12860 163244
rect 12912 163232 12918 163244
rect 16350 163232 16356 163244
rect 12912 163204 16356 163232
rect 12912 163192 12918 163204
rect 16350 163192 16356 163204
rect 16408 163192 16414 163244
rect 360522 162648 360528 162700
rect 360580 162688 360586 162700
rect 418206 162688 418212 162700
rect 360580 162660 418212 162688
rect 360580 162648 360586 162660
rect 418206 162648 418212 162660
rect 418264 162648 418270 162700
rect 226294 162376 226300 162428
rect 226352 162416 226358 162428
rect 230986 162416 230992 162428
rect 226352 162388 230992 162416
rect 226352 162376 226358 162388
rect 230986 162376 230992 162388
rect 231044 162376 231050 162428
rect 131994 162104 132000 162156
rect 132052 162144 132058 162156
rect 138158 162144 138164 162156
rect 132052 162116 138164 162144
rect 132052 162104 132058 162116
rect 138158 162104 138164 162116
rect 138216 162104 138222 162156
rect 131902 162036 131908 162088
rect 131960 162076 131966 162088
rect 139630 162076 139636 162088
rect 131960 162048 139636 162076
rect 131960 162036 131966 162048
rect 139630 162036 139636 162048
rect 139688 162036 139694 162088
rect 178822 162036 178828 162088
rect 178880 162076 178886 162088
rect 181766 162076 181772 162088
rect 178880 162048 181772 162076
rect 178880 162036 178886 162048
rect 181766 162036 181772 162048
rect 181824 162036 181830 162088
rect 226294 162036 226300 162088
rect 226352 162076 226358 162088
rect 233470 162076 233476 162088
rect 226352 162048 233476 162076
rect 226352 162036 226358 162048
rect 233470 162036 233476 162048
rect 233528 162036 233534 162088
rect 266866 162036 266872 162088
rect 266924 162076 266930 162088
rect 274870 162076 274876 162088
rect 266924 162048 274876 162076
rect 266924 162036 266930 162048
rect 274870 162036 274876 162048
rect 274928 162036 274934 162088
rect 321698 162036 321704 162088
rect 321756 162076 321762 162088
rect 328414 162076 328420 162088
rect 321756 162048 328420 162076
rect 321756 162036 321762 162048
rect 328414 162036 328420 162048
rect 328472 162036 328478 162088
rect 77254 161968 77260 162020
rect 77312 162008 77318 162020
rect 87190 162008 87196 162020
rect 77312 161980 87196 162008
rect 77312 161968 77318 161980
rect 87190 161968 87196 161980
rect 87248 161968 87254 162020
rect 131994 161968 132000 162020
rect 132052 162008 132058 162020
rect 132270 162008 132276 162020
rect 132052 161980 132276 162008
rect 132052 161968 132058 161980
rect 132270 161968 132276 161980
rect 132328 161968 132334 162020
rect 85626 161900 85632 161952
rect 85684 161940 85690 161952
rect 87282 161940 87288 161952
rect 85684 161912 87288 161940
rect 85684 161900 85690 161912
rect 87282 161900 87288 161912
rect 87340 161900 87346 161952
rect 222430 161560 222436 161612
rect 222488 161560 222494 161612
rect 172842 161492 172848 161544
rect 172900 161532 172906 161544
rect 222448 161532 222476 161560
rect 172900 161504 222476 161532
rect 172900 161492 172906 161504
rect 320778 161288 320784 161340
rect 320836 161328 320842 161340
rect 327218 161328 327224 161340
rect 320836 161300 327224 161328
rect 320836 161288 320842 161300
rect 327218 161288 327224 161300
rect 327276 161288 327282 161340
rect 232918 160784 232924 160796
rect 231096 160756 232924 160784
rect 131350 160676 131356 160728
rect 131408 160716 131414 160728
rect 140458 160716 140464 160728
rect 131408 160688 140464 160716
rect 131408 160676 131414 160688
rect 140458 160676 140464 160688
rect 140516 160676 140522 160728
rect 131718 160608 131724 160660
rect 131776 160648 131782 160660
rect 139630 160648 139636 160660
rect 131776 160620 139636 160648
rect 131776 160608 131782 160620
rect 139630 160608 139636 160620
rect 139688 160608 139694 160660
rect 173946 160608 173952 160660
rect 174004 160648 174010 160660
rect 177534 160648 177540 160660
rect 174004 160620 177540 160648
rect 174004 160608 174010 160620
rect 177534 160608 177540 160620
rect 177592 160608 177598 160660
rect 179098 160608 179104 160660
rect 179156 160648 179162 160660
rect 182318 160648 182324 160660
rect 179156 160620 182324 160648
rect 179156 160608 179162 160620
rect 182318 160608 182324 160620
rect 182376 160608 182382 160660
rect 226386 160608 226392 160660
rect 226444 160648 226450 160660
rect 231096 160648 231124 160756
rect 232918 160744 232924 160756
rect 232976 160744 232982 160796
rect 266958 160744 266964 160796
rect 267016 160784 267022 160796
rect 267326 160784 267332 160796
rect 267016 160756 267332 160784
rect 267016 160744 267022 160756
rect 267326 160744 267332 160756
rect 267384 160744 267390 160796
rect 271285 160787 271343 160793
rect 271285 160753 271297 160787
rect 271331 160784 271343 160787
rect 274870 160784 274876 160796
rect 271331 160756 274876 160784
rect 271331 160753 271343 160756
rect 271285 160747 271343 160753
rect 274870 160744 274876 160756
rect 274928 160744 274934 160796
rect 266590 160676 266596 160728
rect 266648 160716 266654 160728
rect 274318 160716 274324 160728
rect 266648 160688 274324 160716
rect 266648 160676 266654 160688
rect 274318 160676 274324 160688
rect 274376 160676 274382 160728
rect 226444 160620 231124 160648
rect 226444 160608 226450 160620
rect 231354 160608 231360 160660
rect 231412 160648 231418 160660
rect 233470 160648 233476 160660
rect 231412 160620 233476 160648
rect 231412 160608 231418 160620
rect 233470 160608 233476 160620
rect 233528 160608 233534 160660
rect 267326 160608 267332 160660
rect 267384 160648 267390 160660
rect 271285 160651 271343 160657
rect 271285 160648 271297 160651
rect 267384 160620 271297 160648
rect 267384 160608 267390 160620
rect 271285 160617 271297 160620
rect 271331 160617 271343 160651
rect 271285 160611 271343 160617
rect 271374 160608 271380 160660
rect 271432 160648 271438 160660
rect 274870 160648 274876 160660
rect 271432 160620 274876 160648
rect 271432 160608 271438 160620
rect 274870 160608 274876 160620
rect 274928 160608 274934 160660
rect 77162 160540 77168 160592
rect 77220 160580 77226 160592
rect 87190 160580 87196 160592
rect 77220 160552 87196 160580
rect 77220 160540 77226 160552
rect 87190 160540 87196 160552
rect 87248 160540 87254 160592
rect 225558 159928 225564 159980
rect 225616 159968 225622 159980
rect 226294 159968 226300 159980
rect 225616 159940 226300 159968
rect 225616 159928 225622 159940
rect 226294 159928 226300 159940
rect 226352 159928 226358 159980
rect 173946 159316 173952 159368
rect 174004 159356 174010 159368
rect 180386 159356 180392 159368
rect 174004 159328 180392 159356
rect 174004 159316 174010 159328
rect 180386 159316 180392 159328
rect 180444 159316 180450 159368
rect 226294 159316 226300 159368
rect 226352 159356 226358 159368
rect 232734 159356 232740 159368
rect 226352 159328 232740 159356
rect 226352 159316 226358 159328
rect 232734 159316 232740 159328
rect 232792 159316 232798 159368
rect 79278 159248 79284 159300
rect 79336 159288 79342 159300
rect 79336 159260 85764 159288
rect 79336 159248 79342 159260
rect 85736 159152 85764 159260
rect 137606 159248 137612 159300
rect 137664 159288 137670 159300
rect 139630 159288 139636 159300
rect 137664 159260 139636 159288
rect 137664 159248 137670 159260
rect 139630 159248 139636 159260
rect 139688 159248 139694 159300
rect 178914 159248 178920 159300
rect 178972 159288 178978 159300
rect 182318 159288 182324 159300
rect 178972 159260 182324 159288
rect 178972 159248 178978 159260
rect 182318 159248 182324 159260
rect 182376 159248 182382 159300
rect 227214 159248 227220 159300
rect 227272 159288 227278 159300
rect 233470 159288 233476 159300
rect 227272 159260 233476 159288
rect 227272 159248 227278 159260
rect 233470 159248 233476 159260
rect 233528 159248 233534 159300
rect 266590 159248 266596 159300
rect 266648 159288 266654 159300
rect 274226 159288 274232 159300
rect 266648 159260 274232 159288
rect 266648 159248 266654 159260
rect 274226 159248 274232 159260
rect 274284 159248 274290 159300
rect 87282 159152 87288 159164
rect 85736 159124 87288 159152
rect 87282 159112 87288 159124
rect 87340 159112 87346 159164
rect 81670 159044 81676 159096
rect 81728 159084 81734 159096
rect 87190 159084 87196 159096
rect 81728 159056 87196 159084
rect 81728 159044 81734 159056
rect 87190 159044 87196 159056
rect 87248 159044 87254 159096
rect 361258 158500 361264 158552
rect 361316 158540 361322 158552
rect 415538 158540 415544 158552
rect 361316 158512 415544 158540
rect 361316 158500 361322 158512
rect 415538 158500 415544 158512
rect 415596 158500 415602 158552
rect 321606 158160 321612 158212
rect 321664 158200 321670 158212
rect 327218 158200 327224 158212
rect 321664 158172 327224 158200
rect 321664 158160 321670 158172
rect 327218 158160 327224 158172
rect 327276 158160 327282 158212
rect 321054 158024 321060 158076
rect 321112 158064 321118 158076
rect 327310 158064 327316 158076
rect 321112 158036 327316 158064
rect 321112 158024 321118 158036
rect 327310 158024 327316 158036
rect 327368 158024 327374 158076
rect 131350 157956 131356 158008
rect 131408 157996 131414 158008
rect 138894 157996 138900 158008
rect 131408 157968 138900 157996
rect 131408 157956 131414 157968
rect 138894 157956 138900 157968
rect 138952 157956 138958 158008
rect 173854 157956 173860 158008
rect 173912 157996 173918 158008
rect 173912 157968 176384 157996
rect 173912 157956 173918 157968
rect 79738 157888 79744 157940
rect 79796 157928 79802 157940
rect 87190 157928 87196 157940
rect 79796 157900 87196 157928
rect 79796 157888 79802 157900
rect 87190 157888 87196 157900
rect 87248 157888 87254 157940
rect 131626 157888 131632 157940
rect 131684 157928 131690 157940
rect 139630 157928 139636 157940
rect 131684 157900 139636 157928
rect 131684 157888 131690 157900
rect 139630 157888 139636 157900
rect 139688 157888 139694 157940
rect 173762 157888 173768 157940
rect 173820 157928 173826 157940
rect 176246 157928 176252 157940
rect 173820 157900 176252 157928
rect 173820 157888 173826 157900
rect 176246 157888 176252 157900
rect 176304 157888 176310 157940
rect 176356 157928 176384 157968
rect 226386 157956 226392 158008
rect 226444 157996 226450 158008
rect 228778 157996 228784 158008
rect 226444 157968 228784 157996
rect 226444 157956 226450 157968
rect 228778 157956 228784 157968
rect 228836 157956 228842 158008
rect 266590 157956 266596 158008
rect 266648 157996 266654 158008
rect 274410 157996 274416 158008
rect 266648 157968 274416 157996
rect 266648 157956 266654 157968
rect 274410 157956 274416 157968
rect 274468 157956 274474 158008
rect 182318 157928 182324 157940
rect 176356 157900 182324 157928
rect 182318 157888 182324 157900
rect 182376 157888 182382 157940
rect 227306 157888 227312 157940
rect 227364 157928 227370 157940
rect 233470 157928 233476 157940
rect 227364 157900 233476 157928
rect 227364 157888 227370 157900
rect 233470 157888 233476 157900
rect 233528 157888 233534 157940
rect 321606 157208 321612 157260
rect 321664 157248 321670 157260
rect 327218 157248 327224 157260
rect 321664 157220 327224 157248
rect 321664 157208 321670 157220
rect 327218 157208 327224 157220
rect 327276 157208 327282 157260
rect 222798 157140 222804 157192
rect 222856 157180 222862 157192
rect 233470 157180 233476 157192
rect 222856 157152 233476 157180
rect 222856 157140 222862 157152
rect 233470 157140 233476 157152
rect 233528 157140 233534 157192
rect 77254 156460 77260 156512
rect 77312 156500 77318 156512
rect 77312 156472 85120 156500
rect 77312 156460 77318 156472
rect 85092 156432 85120 156472
rect 173762 156460 173768 156512
rect 173820 156500 173826 156512
rect 181766 156500 181772 156512
rect 173820 156472 181772 156500
rect 173820 156460 173826 156472
rect 181766 156460 181772 156472
rect 181824 156460 181830 156512
rect 87190 156432 87196 156444
rect 85092 156404 87196 156432
rect 87190 156392 87196 156404
rect 87248 156392 87254 156444
rect 173578 156392 173584 156444
rect 173636 156432 173642 156444
rect 182318 156432 182324 156444
rect 173636 156404 182324 156432
rect 173636 156392 173642 156404
rect 182318 156392 182324 156404
rect 182376 156392 182382 156444
rect 267418 156392 267424 156444
rect 267476 156432 267482 156444
rect 274870 156432 274876 156444
rect 267476 156404 274876 156432
rect 267476 156392 267482 156404
rect 274870 156392 274876 156404
rect 274928 156392 274934 156444
rect 358590 156432 358596 156444
rect 358551 156404 358596 156432
rect 358590 156392 358596 156404
rect 358648 156392 358654 156444
rect 321606 155916 321612 155968
rect 321664 155956 321670 155968
rect 327218 155956 327224 155968
rect 321664 155928 327224 155956
rect 321664 155916 321670 155928
rect 327218 155916 327224 155928
rect 327276 155916 327282 155968
rect 173946 155100 173952 155152
rect 174004 155140 174010 155152
rect 182226 155140 182232 155152
rect 174004 155112 182232 155140
rect 174004 155100 174010 155112
rect 182226 155100 182232 155112
rect 182284 155100 182290 155152
rect 267786 155100 267792 155152
rect 267844 155140 267850 155152
rect 274962 155140 274968 155152
rect 267844 155112 274968 155140
rect 267844 155100 267850 155112
rect 274962 155100 274968 155112
rect 275020 155100 275026 155152
rect 321606 155100 321612 155152
rect 321664 155140 321670 155152
rect 321664 155112 321836 155140
rect 321664 155100 321670 155112
rect 79738 155032 79744 155084
rect 79796 155072 79802 155084
rect 87190 155072 87196 155084
rect 79796 155044 87196 155072
rect 79796 155032 79802 155044
rect 87190 155032 87196 155044
rect 87248 155032 87254 155084
rect 138158 155032 138164 155084
rect 138216 155072 138222 155084
rect 139722 155072 139728 155084
rect 138216 155044 139728 155072
rect 138216 155032 138222 155044
rect 139722 155032 139728 155044
rect 139780 155032 139786 155084
rect 174038 155032 174044 155084
rect 174096 155072 174102 155084
rect 179006 155072 179012 155084
rect 174096 155044 179012 155072
rect 174096 155032 174102 155044
rect 179006 155032 179012 155044
rect 179064 155032 179070 155084
rect 181122 155072 181128 155084
rect 179116 155044 181128 155072
rect 173394 154964 173400 155016
rect 173452 155004 173458 155016
rect 179116 155004 179144 155044
rect 181122 155032 181128 155044
rect 181180 155032 181186 155084
rect 230986 155032 230992 155084
rect 231044 155072 231050 155084
rect 234022 155072 234028 155084
rect 231044 155044 234028 155072
rect 231044 155032 231050 155044
rect 234022 155032 234028 155044
rect 234080 155032 234086 155084
rect 267694 155032 267700 155084
rect 267752 155072 267758 155084
rect 274870 155072 274876 155084
rect 267752 155044 274876 155072
rect 267752 155032 267758 155044
rect 274870 155032 274876 155044
rect 274928 155032 274934 155084
rect 321808 155072 321836 155112
rect 328414 155072 328420 155084
rect 321808 155044 328420 155072
rect 328414 155032 328420 155044
rect 328472 155032 328478 155084
rect 173452 154976 179144 155004
rect 173452 154964 173458 154976
rect 266590 154964 266596 155016
rect 266648 155004 266654 155016
rect 274502 155004 274508 155016
rect 266648 154976 274508 155004
rect 266648 154964 266654 154976
rect 274502 154964 274508 154976
rect 274560 154964 274566 155016
rect 267050 154896 267056 154948
rect 267108 154936 267114 154948
rect 267694 154936 267700 154948
rect 267108 154908 267700 154936
rect 267108 154896 267114 154908
rect 267694 154896 267700 154908
rect 267752 154896 267758 154948
rect 79738 154352 79744 154404
rect 79796 154392 79802 154404
rect 87190 154392 87196 154404
rect 79796 154364 87196 154392
rect 79796 154352 79802 154364
rect 87190 154352 87196 154364
rect 87248 154352 87254 154404
rect 172934 153876 172940 153928
rect 172992 153916 172998 153928
rect 178822 153916 178828 153928
rect 172992 153888 178828 153916
rect 172992 153876 172998 153888
rect 178822 153876 178828 153888
rect 178880 153876 178886 153928
rect 368526 153808 368532 153860
rect 368584 153848 368590 153860
rect 368986 153848 368992 153860
rect 368584 153820 368992 153848
rect 368584 153808 368590 153820
rect 368986 153808 368992 153820
rect 369044 153808 369050 153860
rect 320870 153740 320876 153792
rect 320928 153780 320934 153792
rect 328414 153780 328420 153792
rect 320928 153752 328420 153780
rect 320928 153740 320934 153752
rect 328414 153740 328420 153752
rect 328472 153740 328478 153792
rect 131534 153672 131540 153724
rect 131592 153712 131598 153724
rect 139630 153712 139636 153724
rect 131592 153684 139636 153712
rect 131592 153672 131598 153684
rect 139630 153672 139636 153684
rect 139688 153672 139694 153724
rect 173302 153672 173308 153724
rect 173360 153712 173366 153724
rect 181398 153712 181404 153724
rect 173360 153684 181404 153712
rect 173360 153672 173366 153684
rect 181398 153672 181404 153684
rect 181456 153672 181462 153724
rect 267142 153672 267148 153724
rect 267200 153712 267206 153724
rect 274962 153712 274968 153724
rect 267200 153684 274968 153712
rect 267200 153672 267206 153684
rect 274962 153672 274968 153684
rect 275020 153672 275026 153724
rect 427498 153672 427504 153724
rect 427556 153712 427562 153724
rect 429430 153712 429436 153724
rect 427556 153684 429436 153712
rect 427556 153672 427562 153684
rect 429430 153672 429436 153684
rect 429488 153672 429494 153724
rect 173486 153604 173492 153656
rect 173544 153644 173550 153656
rect 181950 153644 181956 153656
rect 173544 153616 181956 153644
rect 173544 153604 173550 153616
rect 181950 153604 181956 153616
rect 182008 153604 182014 153656
rect 267510 153604 267516 153656
rect 267568 153644 267574 153656
rect 274870 153644 274876 153656
rect 267568 153616 274876 153644
rect 267568 153604 267574 153616
rect 274870 153604 274876 153616
rect 274928 153604 274934 153656
rect 173210 153128 173216 153180
rect 173268 153168 173274 153180
rect 179098 153168 179104 153180
rect 173268 153140 179104 153168
rect 173268 153128 173274 153140
rect 179098 153128 179104 153140
rect 179156 153128 179162 153180
rect 79738 152992 79744 153044
rect 79796 153032 79802 153044
rect 87190 153032 87196 153044
rect 79796 153004 87196 153032
rect 79796 152992 79802 153004
rect 87190 152992 87196 153004
rect 87248 152992 87254 153044
rect 320502 152448 320508 152500
rect 320560 152488 320566 152500
rect 323170 152488 323176 152500
rect 320560 152460 323176 152488
rect 320560 152448 320566 152460
rect 323170 152448 323176 152460
rect 323228 152448 323234 152500
rect 85810 152380 85816 152432
rect 85868 152420 85874 152432
rect 87190 152420 87196 152432
rect 85868 152392 87196 152420
rect 85868 152380 85874 152392
rect 87190 152380 87196 152392
rect 87248 152380 87254 152432
rect 321606 152380 321612 152432
rect 321664 152420 321670 152432
rect 328414 152420 328420 152432
rect 321664 152392 328420 152420
rect 321664 152380 321670 152392
rect 328414 152380 328420 152392
rect 328472 152380 328478 152432
rect 174038 152312 174044 152364
rect 174096 152352 174102 152364
rect 182318 152352 182324 152364
rect 174096 152324 182324 152352
rect 174096 152312 174102 152324
rect 182318 152312 182324 152324
rect 182376 152312 182382 152364
rect 267878 152312 267884 152364
rect 267936 152352 267942 152364
rect 274870 152352 274876 152364
rect 267936 152324 274876 152352
rect 267936 152312 267942 152324
rect 274870 152312 274876 152324
rect 274928 152312 274934 152364
rect 368526 152312 368532 152364
rect 368584 152352 368590 152364
rect 368710 152352 368716 152364
rect 368584 152324 368716 152352
rect 368584 152312 368590 152324
rect 368710 152312 368716 152324
rect 368768 152312 368774 152364
rect 85902 151360 85908 151412
rect 85960 151400 85966 151412
rect 87466 151400 87472 151412
rect 85960 151372 87472 151400
rect 85960 151360 85966 151372
rect 87466 151360 87472 151372
rect 87524 151360 87530 151412
rect 320778 151360 320784 151412
rect 320836 151400 320842 151412
rect 323262 151400 323268 151412
rect 320836 151372 323268 151400
rect 320836 151360 320842 151372
rect 323262 151360 323268 151372
rect 323320 151360 323326 151412
rect 225558 150952 225564 151004
rect 225616 150992 225622 151004
rect 226202 150992 226208 151004
rect 225616 150964 226208 150992
rect 225616 150952 225622 150964
rect 226202 150952 226208 150964
rect 226260 150952 226266 151004
rect 173670 150884 173676 150936
rect 173728 150924 173734 150936
rect 182318 150924 182324 150936
rect 173728 150896 182324 150924
rect 173728 150884 173734 150896
rect 182318 150884 182324 150896
rect 182376 150884 182382 150936
rect 225650 150884 225656 150936
rect 225708 150924 225714 150936
rect 233470 150924 233476 150936
rect 225708 150896 233476 150924
rect 225708 150884 225714 150896
rect 233470 150884 233476 150896
rect 233528 150884 233534 150936
rect 267694 150884 267700 150936
rect 267752 150924 267758 150936
rect 274870 150924 274876 150936
rect 267752 150896 274876 150924
rect 267752 150884 267758 150896
rect 274870 150884 274876 150896
rect 274928 150884 274934 150936
rect 323170 150884 323176 150936
rect 323228 150924 323234 150936
rect 328414 150924 328420 150936
rect 323228 150896 328420 150924
rect 323228 150884 323234 150896
rect 328414 150884 328420 150896
rect 328472 150884 328478 150936
rect 177534 150816 177540 150868
rect 177592 150856 177598 150868
rect 182226 150856 182232 150868
rect 177592 150828 182232 150856
rect 177592 150816 177598 150828
rect 182226 150816 182232 150828
rect 182284 150816 182290 150868
rect 225558 150816 225564 150868
rect 225616 150856 225622 150868
rect 231354 150856 231360 150868
rect 225616 150828 231360 150856
rect 225616 150816 225622 150828
rect 231354 150816 231360 150828
rect 231412 150816 231418 150868
rect 266590 150816 266596 150868
rect 266648 150856 266654 150868
rect 271374 150856 271380 150868
rect 266648 150828 271380 150856
rect 266648 150816 266654 150828
rect 271374 150816 271380 150828
rect 271432 150816 271438 150868
rect 174038 150748 174044 150800
rect 174096 150788 174102 150800
rect 181030 150788 181036 150800
rect 174096 150760 181036 150788
rect 174096 150748 174102 150760
rect 181030 150748 181036 150760
rect 181088 150748 181094 150800
rect 181030 150612 181036 150664
rect 181088 150652 181094 150664
rect 181674 150652 181680 150664
rect 181088 150624 181680 150652
rect 181088 150612 181094 150624
rect 181674 150612 181680 150624
rect 181732 150612 181738 150664
rect 77254 149796 77260 149848
rect 77312 149836 77318 149848
rect 85810 149836 85816 149848
rect 77312 149808 85816 149836
rect 77312 149796 77318 149808
rect 85810 149796 85816 149808
rect 85868 149796 85874 149848
rect 321606 149728 321612 149780
rect 321664 149768 321670 149780
rect 327218 149768 327224 149780
rect 321664 149740 327224 149768
rect 321664 149728 321670 149740
rect 327218 149728 327224 149740
rect 327276 149728 327282 149780
rect 80106 149592 80112 149644
rect 80164 149632 80170 149644
rect 87190 149632 87196 149644
rect 80164 149604 87196 149632
rect 80164 149592 80170 149604
rect 87190 149592 87196 149604
rect 87248 149592 87254 149644
rect 321054 149592 321060 149644
rect 321112 149632 321118 149644
rect 323170 149632 323176 149644
rect 321112 149604 323176 149632
rect 321112 149592 321118 149604
rect 323170 149592 323176 149604
rect 323228 149592 323234 149644
rect 131810 149524 131816 149576
rect 131868 149564 131874 149576
rect 139630 149564 139636 149576
rect 131868 149536 139636 149564
rect 131868 149524 131874 149536
rect 139630 149524 139636 149536
rect 139688 149524 139694 149576
rect 176246 149524 176252 149576
rect 176304 149564 176310 149576
rect 182318 149564 182324 149576
rect 176304 149536 182324 149564
rect 176304 149524 176310 149536
rect 182318 149524 182324 149536
rect 182376 149524 182382 149576
rect 323262 149524 323268 149576
rect 323320 149564 323326 149576
rect 328414 149564 328420 149576
rect 323320 149536 328420 149564
rect 323320 149524 323326 149536
rect 328414 149524 328420 149536
rect 328472 149524 328478 149576
rect 131350 149456 131356 149508
rect 131408 149496 131414 149508
rect 137606 149496 137612 149508
rect 131408 149468 137612 149496
rect 131408 149456 131414 149468
rect 137606 149456 137612 149468
rect 137664 149456 137670 149508
rect 174038 149456 174044 149508
rect 174096 149496 174102 149508
rect 178914 149496 178920 149508
rect 174096 149468 178920 149496
rect 174096 149456 174102 149468
rect 178914 149456 178920 149468
rect 178972 149456 178978 149508
rect 225282 149388 225288 149440
rect 225340 149428 225346 149440
rect 227214 149428 227220 149440
rect 225340 149400 227220 149428
rect 225340 149388 225346 149400
rect 227214 149388 227220 149400
rect 227272 149388 227278 149440
rect 266590 149388 266596 149440
rect 266648 149428 266654 149440
rect 275698 149428 275704 149440
rect 266648 149400 275704 149428
rect 266648 149388 266654 149400
rect 275698 149388 275704 149400
rect 275756 149388 275762 149440
rect 12854 149320 12860 149372
rect 12912 149360 12918 149372
rect 16258 149360 16264 149372
rect 12912 149332 16264 149360
rect 12912 149320 12918 149332
rect 16258 149320 16264 149332
rect 16316 149320 16322 149372
rect 225190 148640 225196 148692
rect 225248 148680 225254 148692
rect 227306 148680 227312 148692
rect 225248 148652 227312 148680
rect 225248 148640 225254 148652
rect 227306 148640 227312 148652
rect 227364 148640 227370 148692
rect 78910 148436 78916 148488
rect 78968 148476 78974 148488
rect 85902 148476 85908 148488
rect 78968 148448 85908 148476
rect 78968 148436 78974 148448
rect 85902 148436 85908 148448
rect 85960 148436 85966 148488
rect 321606 148368 321612 148420
rect 321664 148408 321670 148420
rect 327862 148408 327868 148420
rect 321664 148380 327868 148408
rect 321664 148368 321670 148380
rect 327862 148368 327868 148380
rect 327920 148368 327926 148420
rect 174038 148164 174044 148216
rect 174096 148204 174102 148216
rect 180294 148204 180300 148216
rect 174096 148176 180300 148204
rect 174096 148164 174102 148176
rect 180294 148164 180300 148176
rect 180352 148164 180358 148216
rect 228778 148164 228784 148216
rect 228836 148204 228842 148216
rect 233470 148204 233476 148216
rect 228836 148176 233476 148204
rect 228836 148164 228842 148176
rect 233470 148164 233476 148176
rect 233528 148164 233534 148216
rect 266590 148164 266596 148216
rect 266648 148204 266654 148216
rect 274134 148204 274140 148216
rect 266648 148176 274140 148204
rect 266648 148164 266654 148176
rect 274134 148164 274140 148176
rect 274192 148164 274198 148216
rect 323170 148164 323176 148216
rect 323228 148204 323234 148216
rect 328414 148204 328420 148216
rect 323228 148176 328420 148204
rect 323228 148164 323234 148176
rect 328414 148164 328420 148176
rect 328472 148164 328478 148216
rect 78910 147688 78916 147740
rect 78968 147728 78974 147740
rect 87006 147728 87012 147740
rect 78968 147700 87012 147728
rect 78968 147688 78974 147700
rect 87006 147688 87012 147700
rect 87064 147688 87070 147740
rect 132270 146736 132276 146788
rect 132328 146776 132334 146788
rect 140550 146776 140556 146788
rect 132328 146748 140556 146776
rect 132328 146736 132334 146748
rect 140550 146736 140556 146748
rect 140608 146736 140614 146788
rect 226294 146736 226300 146788
rect 226352 146776 226358 146788
rect 233470 146776 233476 146788
rect 226352 146748 233476 146776
rect 226352 146736 226358 146748
rect 233470 146736 233476 146748
rect 233528 146736 233534 146788
rect 267878 146736 267884 146788
rect 267936 146776 267942 146788
rect 275514 146776 275520 146788
rect 267936 146748 275520 146776
rect 267936 146736 267942 146748
rect 275514 146736 275520 146748
rect 275572 146736 275578 146788
rect 79370 145376 79376 145428
rect 79428 145416 79434 145428
rect 87190 145416 87196 145428
rect 79428 145388 87196 145416
rect 79428 145376 79434 145388
rect 87190 145376 87196 145388
rect 87248 145376 87254 145428
rect 91698 145376 91704 145428
rect 91756 145416 91762 145428
rect 128130 145416 128136 145428
rect 91756 145388 128136 145416
rect 91756 145376 91762 145388
rect 128130 145376 128136 145388
rect 128188 145376 128194 145428
rect 132454 145376 132460 145428
rect 132512 145416 132518 145428
rect 140550 145416 140556 145428
rect 132512 145388 140556 145416
rect 132512 145376 132518 145388
rect 140550 145376 140556 145388
rect 140608 145376 140614 145428
rect 185630 145376 185636 145428
rect 185688 145416 185694 145428
rect 222154 145416 222160 145428
rect 185688 145388 222160 145416
rect 185688 145376 185694 145388
rect 222154 145376 222160 145388
rect 222212 145376 222218 145428
rect 226386 145376 226392 145428
rect 226444 145416 226450 145428
rect 233470 145416 233476 145428
rect 226444 145388 233476 145416
rect 226444 145376 226450 145388
rect 233470 145376 233476 145388
rect 233528 145376 233534 145428
rect 266774 145376 266780 145428
rect 266832 145416 266838 145428
rect 275606 145416 275612 145428
rect 266832 145388 275612 145416
rect 266832 145376 266838 145388
rect 275606 145376 275612 145388
rect 275664 145376 275670 145428
rect 279654 145376 279660 145428
rect 279712 145416 279718 145428
rect 322802 145416 322808 145428
rect 279712 145388 322808 145416
rect 279712 145376 279718 145388
rect 322802 145376 322808 145388
rect 322860 145376 322866 145428
rect 116078 144832 116084 144884
rect 116136 144872 116142 144884
rect 128038 144872 128044 144884
rect 116136 144844 128044 144872
rect 116136 144832 116142 144844
rect 128038 144832 128044 144844
rect 128096 144832 128102 144884
rect 292718 144832 292724 144884
rect 292776 144872 292782 144884
rect 312314 144872 312320 144884
rect 292776 144844 312320 144872
rect 292776 144832 292782 144844
rect 312314 144832 312320 144844
rect 312372 144832 312378 144884
rect 103658 144764 103664 144816
rect 103716 144804 103722 144816
rect 124266 144804 124272 144816
rect 103716 144776 124272 144804
rect 103716 144764 103722 144776
rect 124266 144764 124272 144776
rect 124324 144764 124330 144816
rect 171278 144764 171284 144816
rect 171336 144804 171342 144816
rect 189218 144804 189224 144816
rect 171336 144776 189224 144804
rect 171336 144764 171342 144776
rect 189218 144764 189224 144776
rect 189276 144764 189282 144816
rect 197498 144764 197504 144816
rect 197556 144804 197562 144816
rect 218290 144804 218296 144816
rect 197556 144776 218296 144804
rect 197556 144764 197562 144776
rect 218290 144764 218296 144776
rect 218348 144764 218354 144816
rect 280298 144764 280304 144816
rect 280356 144804 280362 144816
rect 308726 144804 308732 144816
rect 280356 144776 308732 144804
rect 280356 144764 280362 144776
rect 308726 144764 308732 144776
rect 308784 144764 308790 144816
rect 91238 144696 91244 144748
rect 91296 144736 91302 144748
rect 120678 144736 120684 144748
rect 91296 144708 120684 144736
rect 91296 144696 91302 144708
rect 120678 144696 120684 144708
rect 120736 144696 120742 144748
rect 185078 144696 185084 144748
rect 185136 144736 185142 144748
rect 214702 144736 214708 144748
rect 185136 144708 214708 144736
rect 185136 144696 185142 144708
rect 214702 144696 214708 144708
rect 214760 144696 214766 144748
rect 218934 144696 218940 144748
rect 218992 144736 218998 144748
rect 221970 144736 221976 144748
rect 218992 144708 221976 144736
rect 218992 144696 218998 144708
rect 221970 144696 221976 144708
rect 222028 144696 222034 144748
rect 290510 144696 290516 144748
rect 290568 144736 290574 144748
rect 326574 144736 326580 144748
rect 290568 144708 326580 144736
rect 290568 144696 290574 144708
rect 326574 144696 326580 144708
rect 326632 144696 326638 144748
rect 312774 144084 312780 144136
rect 312832 144124 312838 144136
rect 315994 144124 316000 144136
rect 312832 144096 316000 144124
rect 312832 144084 312838 144096
rect 315994 144084 316000 144096
rect 316052 144084 316058 144136
rect 132362 144016 132368 144068
rect 132420 144056 132426 144068
rect 140550 144056 140556 144068
rect 132420 144028 140556 144056
rect 132420 144016 132426 144028
rect 140550 144016 140556 144028
rect 140608 144016 140614 144068
rect 226478 144016 226484 144068
rect 226536 144056 226542 144068
rect 233470 144056 233476 144068
rect 226536 144028 233476 144056
rect 226536 144016 226542 144028
rect 233470 144016 233476 144028
rect 233528 144016 233534 144068
rect 321790 144016 321796 144068
rect 321848 144056 321854 144068
rect 327310 144056 327316 144068
rect 321848 144028 327316 144056
rect 321848 144016 321854 144028
rect 327310 144016 327316 144028
rect 327368 144016 327374 144068
rect 76061 143991 76119 143997
rect 76061 143957 76073 143991
rect 76107 143988 76119 143991
rect 87101 143991 87159 143997
rect 87101 143988 87113 143991
rect 76107 143960 87113 143988
rect 76107 143957 76119 143960
rect 76061 143951 76119 143957
rect 87101 143957 87113 143960
rect 87147 143957 87159 143991
rect 87101 143951 87159 143957
rect 95286 143920 95292 143932
rect 89876 143892 95292 143920
rect 87101 143855 87159 143861
rect 87101 143821 87113 143855
rect 87147 143852 87159 143855
rect 89876 143852 89904 143892
rect 95286 143880 95292 143892
rect 95344 143880 95350 143932
rect 87147 143824 89904 143852
rect 87147 143821 87159 143824
rect 87101 143815 87159 143821
rect 211022 143404 211028 143456
rect 211080 143444 211086 143456
rect 231354 143444 231360 143456
rect 211080 143416 231360 143444
rect 211080 143404 211086 143416
rect 231354 143404 231360 143416
rect 231412 143404 231418 143456
rect 76886 143336 76892 143388
rect 76944 143376 76950 143388
rect 88570 143376 88576 143388
rect 76944 143348 88576 143376
rect 76944 143336 76950 143348
rect 88570 143336 88576 143348
rect 88628 143336 88634 143388
rect 203754 143336 203760 143388
rect 203812 143376 203818 143388
rect 231170 143376 231176 143388
rect 203812 143348 231176 143376
rect 203812 143336 203818 143348
rect 231170 143336 231176 143348
rect 231228 143336 231234 143388
rect 294282 143336 294288 143388
rect 294340 143376 294346 143388
rect 325286 143376 325292 143388
rect 294340 143348 325292 143376
rect 294340 143336 294346 143348
rect 325286 143336 325292 143348
rect 325344 143336 325350 143388
rect 78910 143200 78916 143252
rect 78968 143240 78974 143252
rect 87098 143240 87104 143252
rect 78968 143212 87104 143240
rect 78968 143200 78974 143212
rect 87098 143200 87104 143212
rect 87156 143200 87162 143252
rect 200166 142288 200172 142300
rect 167984 142260 200172 142288
rect 167984 142232 168012 142260
rect 200166 142248 200172 142260
rect 200224 142248 200230 142300
rect 309373 142291 309431 142297
rect 261916 142260 296996 142288
rect 261916 142232 261944 142260
rect 167966 142180 167972 142232
rect 168024 142180 168030 142232
rect 168518 142180 168524 142232
rect 168576 142220 168582 142232
rect 196854 142220 196860 142232
rect 168576 142192 196860 142220
rect 168576 142180 168582 142192
rect 196854 142180 196860 142192
rect 196912 142180 196918 142232
rect 236874 142180 236880 142232
rect 236932 142220 236938 142232
rect 238990 142220 238996 142232
rect 236932 142192 238996 142220
rect 236932 142180 236938 142192
rect 238990 142180 238996 142192
rect 239048 142220 239054 142232
rect 239910 142220 239916 142232
rect 239048 142192 239916 142220
rect 239048 142180 239054 142192
rect 239910 142180 239916 142192
rect 239968 142180 239974 142232
rect 261898 142180 261904 142232
rect 261956 142180 261962 142232
rect 296968 142220 296996 142260
rect 309373 142257 309385 142291
rect 309419 142288 309431 142291
rect 318941 142291 318999 142297
rect 318941 142288 318953 142291
rect 309419 142260 318953 142288
rect 309419 142257 309431 142260
rect 309373 142251 309431 142257
rect 318941 142257 318953 142260
rect 318987 142257 318999 142291
rect 318941 142251 318999 142257
rect 302473 142223 302531 142229
rect 302473 142220 302485 142223
rect 296968 142192 302485 142220
rect 302473 142189 302485 142192
rect 302519 142189 302531 142223
rect 302473 142183 302531 142189
rect 318941 142155 318999 142161
rect 318941 142121 318953 142155
rect 318987 142152 318999 142155
rect 318987 142124 321652 142152
rect 318987 142121 318999 142124
rect 318941 142115 318999 142121
rect 76058 142084 76064 142096
rect 76019 142056 76064 142084
rect 76058 142044 76064 142056
rect 76116 142044 76122 142096
rect 302473 142087 302531 142093
rect 302473 142053 302485 142087
rect 302519 142084 302531 142087
rect 305046 142084 305052 142096
rect 302519 142056 305052 142084
rect 302519 142053 302531 142056
rect 302473 142047 302531 142053
rect 305046 142044 305052 142056
rect 305104 142084 305110 142096
rect 309373 142087 309431 142093
rect 309373 142084 309385 142087
rect 305104 142056 309385 142084
rect 305104 142044 305110 142056
rect 309373 142053 309385 142056
rect 309419 142053 309431 142087
rect 321624 142084 321652 142124
rect 324550 142084 324556 142096
rect 321624 142056 324556 142084
rect 309373 142047 309431 142053
rect 324550 142044 324556 142056
rect 324608 142044 324614 142096
rect 127578 141976 127584 142028
rect 127636 142016 127642 142028
rect 140366 142016 140372 142028
rect 127636 141988 140372 142016
rect 127636 141976 127642 141988
rect 140366 141976 140372 141988
rect 140424 141976 140430 142028
rect 173578 141976 173584 142028
rect 173636 142016 173642 142028
rect 219670 142016 219676 142028
rect 173636 141988 219676 142016
rect 173636 141976 173642 141988
rect 219670 141976 219676 141988
rect 219728 142016 219734 142028
rect 233470 142016 233476 142028
rect 219728 141988 233476 142016
rect 219728 141976 219734 141988
rect 233470 141976 233476 141988
rect 233528 141976 233534 142028
rect 267326 141976 267332 142028
rect 267384 142016 267390 142028
rect 316270 142016 316276 142028
rect 267384 141988 316276 142016
rect 267384 141976 267390 141988
rect 316270 141976 316276 141988
rect 316328 141976 316334 142028
rect 136870 141364 136876 141416
rect 136928 141404 136934 141416
rect 150394 141404 150400 141416
rect 136928 141376 150400 141404
rect 136928 141364 136934 141376
rect 150394 141364 150400 141376
rect 150452 141404 150458 141416
rect 167966 141404 167972 141416
rect 150452 141376 167972 141404
rect 150452 141364 150458 141376
rect 167966 141364 167972 141376
rect 168024 141364 168030 141416
rect 78910 141296 78916 141348
rect 78968 141336 78974 141348
rect 127210 141336 127216 141348
rect 78968 141308 127216 141336
rect 78968 141296 78974 141308
rect 127210 141296 127216 141308
rect 127268 141336 127274 141348
rect 127578 141336 127584 141348
rect 127268 141308 127584 141336
rect 127268 141296 127274 141308
rect 127578 141296 127584 141308
rect 127636 141296 127642 141348
rect 147450 141296 147456 141348
rect 147508 141336 147514 141348
rect 171278 141336 171284 141348
rect 147508 141308 171284 141336
rect 147508 141296 147514 141308
rect 171278 141296 171284 141308
rect 171336 141296 171342 141348
rect 231354 141296 231360 141348
rect 231412 141336 231418 141348
rect 246902 141336 246908 141348
rect 231412 141308 246908 141336
rect 231412 141296 231418 141308
rect 246902 141296 246908 141308
rect 246960 141336 246966 141348
rect 261898 141336 261904 141348
rect 246960 141308 261904 141336
rect 246960 141296 246966 141308
rect 261898 141296 261904 141308
rect 261956 141296 261962 141348
rect 316270 141296 316276 141348
rect 316328 141336 316334 141348
rect 327310 141336 327316 141348
rect 316328 141308 327316 141336
rect 316328 141296 316334 141308
rect 327310 141296 327316 141308
rect 327368 141296 327374 141348
rect 74126 141228 74132 141280
rect 74184 141268 74190 141280
rect 75414 141268 75420 141280
rect 74184 141240 75420 141268
rect 74184 141228 74190 141240
rect 75414 141228 75420 141240
rect 75472 141268 75478 141280
rect 113410 141268 113416 141280
rect 75472 141240 113416 141268
rect 75472 141228 75478 141240
rect 113410 141228 113416 141240
rect 113468 141268 113474 141280
rect 113870 141268 113876 141280
rect 113468 141240 113876 141268
rect 113468 141228 113474 141240
rect 113870 141228 113876 141240
rect 113928 141228 113934 141280
rect 231170 141228 231176 141280
rect 231228 141268 231234 141280
rect 231446 141268 231452 141280
rect 231228 141240 231452 141268
rect 231228 141228 231234 141240
rect 231446 141228 231452 141240
rect 231504 141228 231510 141280
rect 427314 140752 427320 140804
rect 427372 140792 427378 140804
rect 429522 140792 429528 140804
rect 427372 140764 429528 140792
rect 427372 140752 427378 140764
rect 429522 140752 429528 140764
rect 429580 140752 429586 140804
rect 113870 140616 113876 140668
rect 113928 140656 113934 140668
rect 137238 140656 137244 140668
rect 113928 140628 137244 140656
rect 113928 140616 113934 140628
rect 137238 140616 137244 140628
rect 137296 140616 137302 140668
rect 73942 140548 73948 140600
rect 74000 140588 74006 140600
rect 102370 140588 102376 140600
rect 74000 140560 102376 140588
rect 74000 140548 74006 140560
rect 102370 140548 102376 140560
rect 102428 140588 102434 140600
rect 137330 140588 137336 140600
rect 102428 140560 137336 140588
rect 102428 140548 102434 140560
rect 137330 140548 137336 140560
rect 137388 140548 137394 140600
rect 207250 140548 207256 140600
rect 207308 140588 207314 140600
rect 231078 140588 231084 140600
rect 207308 140560 231084 140588
rect 207308 140548 207314 140560
rect 231078 140548 231084 140560
rect 231136 140548 231142 140600
rect 301090 140548 301096 140600
rect 301148 140588 301154 140600
rect 325102 140588 325108 140600
rect 301148 140560 325108 140588
rect 301148 140548 301154 140560
rect 325102 140548 325108 140560
rect 325160 140548 325166 140600
rect 76058 140180 76064 140192
rect 76019 140152 76064 140180
rect 76058 140140 76064 140152
rect 76116 140140 76122 140192
rect 158769 139911 158827 139917
rect 158769 139877 158781 139911
rect 158815 139908 158827 139911
rect 164562 139908 164568 139920
rect 158815 139880 164568 139908
rect 158815 139877 158827 139880
rect 158769 139871 158827 139877
rect 164562 139868 164568 139880
rect 164620 139868 164626 139920
rect 251134 139868 251140 139920
rect 251192 139908 251198 139920
rect 253986 139908 253992 139920
rect 251192 139880 253992 139908
rect 251192 139868 251198 139880
rect 253986 139868 253992 139880
rect 254044 139868 254050 139920
rect 150578 139800 150584 139852
rect 150636 139840 150642 139852
rect 162262 139840 162268 139852
rect 150636 139812 162268 139840
rect 150636 139800 150642 139812
rect 162262 139800 162268 139812
rect 162320 139800 162326 139852
rect 239542 139800 239548 139852
rect 239600 139840 239606 139852
rect 322710 139840 322716 139852
rect 239600 139812 322716 139840
rect 239600 139800 239606 139812
rect 322710 139800 322716 139812
rect 322768 139800 322774 139852
rect 64834 139732 64840 139784
rect 64892 139772 64898 139784
rect 70446 139772 70452 139784
rect 64892 139744 70452 139772
rect 64892 139732 64898 139744
rect 70446 139732 70452 139744
rect 70504 139732 70510 139784
rect 156098 139732 156104 139784
rect 156156 139772 156162 139784
rect 157570 139772 157576 139784
rect 156156 139744 157576 139772
rect 156156 139732 156162 139744
rect 157570 139732 157576 139744
rect 157628 139732 157634 139784
rect 169990 139772 169996 139784
rect 157680 139744 169996 139772
rect 63638 139664 63644 139716
rect 63696 139704 63702 139716
rect 75230 139704 75236 139716
rect 63696 139676 75236 139704
rect 63696 139664 63702 139676
rect 75230 139664 75236 139676
rect 75288 139664 75294 139716
rect 151774 139664 151780 139716
rect 151832 139704 151838 139716
rect 157389 139707 157447 139713
rect 157389 139704 157401 139707
rect 151832 139676 157401 139704
rect 151832 139664 151838 139676
rect 157389 139673 157401 139676
rect 157435 139673 157447 139707
rect 157389 139667 157447 139673
rect 157478 139664 157484 139716
rect 157536 139704 157542 139716
rect 157680 139704 157708 139744
rect 169990 139732 169996 139744
rect 170048 139732 170054 139784
rect 241750 139732 241756 139784
rect 241808 139772 241814 139784
rect 244970 139772 244976 139784
rect 241808 139744 244976 139772
rect 241808 139732 241814 139744
rect 244970 139732 244976 139744
rect 245028 139732 245034 139784
rect 247086 139732 247092 139784
rect 247144 139772 247150 139784
rect 259230 139772 259236 139784
rect 247144 139744 259236 139772
rect 247144 139732 247150 139744
rect 259230 139732 259236 139744
rect 259288 139732 259294 139784
rect 157536 139676 157708 139704
rect 157536 139664 157542 139676
rect 160054 139664 160060 139716
rect 160112 139704 160118 139716
rect 162630 139704 162636 139716
rect 160112 139676 162636 139704
rect 160112 139664 160118 139676
rect 162630 139664 162636 139676
rect 162688 139664 162694 139716
rect 162725 139707 162783 139713
rect 162725 139673 162737 139707
rect 162771 139704 162783 139707
rect 169070 139704 169076 139716
rect 162771 139676 169076 139704
rect 162771 139673 162783 139676
rect 162725 139667 162783 139673
rect 169070 139664 169076 139676
rect 169128 139664 169134 139716
rect 244326 139664 244332 139716
rect 244384 139704 244390 139716
rect 256286 139704 256292 139716
rect 244384 139676 256292 139704
rect 244384 139664 244390 139676
rect 256286 139664 256292 139676
rect 256344 139664 256350 139716
rect 62258 139596 62264 139648
rect 62316 139636 62322 139648
rect 74218 139636 74224 139648
rect 62316 139608 74224 139636
rect 62316 139596 62322 139608
rect 74218 139596 74224 139608
rect 74276 139596 74282 139648
rect 156098 139596 156104 139648
rect 156156 139636 156162 139648
rect 157573 139639 157631 139645
rect 157573 139636 157585 139639
rect 156156 139608 157585 139636
rect 156156 139596 156162 139608
rect 157573 139605 157585 139608
rect 157619 139605 157631 139639
rect 157573 139599 157631 139605
rect 249202 139596 249208 139648
rect 249260 139636 249266 139648
rect 252054 139636 252060 139648
rect 249260 139608 252060 139636
rect 249260 139596 249266 139608
rect 252054 139596 252060 139608
rect 252112 139596 252118 139648
rect 264106 139636 264112 139648
rect 253176 139608 264112 139636
rect 60878 139528 60884 139580
rect 60936 139568 60942 139580
rect 73114 139568 73120 139580
rect 60936 139540 73120 139568
rect 60936 139528 60942 139540
rect 73114 139528 73120 139540
rect 73172 139528 73178 139580
rect 154258 139528 154264 139580
rect 154316 139568 154322 139580
rect 157294 139568 157300 139580
rect 154316 139540 157300 139568
rect 154316 139528 154322 139540
rect 157294 139528 157300 139540
rect 157352 139528 157358 139580
rect 157389 139571 157447 139577
rect 157389 139537 157401 139571
rect 157435 139568 157447 139571
rect 158769 139571 158827 139577
rect 158769 139568 158781 139571
rect 157435 139540 158781 139568
rect 157435 139537 157447 139540
rect 157389 139531 157447 139537
rect 158769 139537 158781 139540
rect 158815 139537 158827 139571
rect 158769 139531 158827 139537
rect 158858 139528 158864 139580
rect 158916 139568 158922 139580
rect 160974 139568 160980 139580
rect 158916 139540 160980 139568
rect 158916 139528 158922 139540
rect 160974 139528 160980 139540
rect 161032 139528 161038 139580
rect 161986 139528 161992 139580
rect 162044 139568 162050 139580
rect 162998 139568 163004 139580
rect 162044 139540 163004 139568
rect 162044 139528 162050 139540
rect 162998 139528 163004 139540
rect 163056 139528 163062 139580
rect 241474 139528 241480 139580
rect 241532 139568 241538 139580
rect 249662 139568 249668 139580
rect 241532 139540 249668 139568
rect 241532 139528 241538 139540
rect 249662 139528 249668 139540
rect 249720 139528 249726 139580
rect 249846 139528 249852 139580
rect 249904 139568 249910 139580
rect 253066 139568 253072 139580
rect 249904 139540 253072 139568
rect 249904 139528 249910 139540
rect 253066 139528 253072 139540
rect 253124 139528 253130 139580
rect 59498 139460 59504 139512
rect 59556 139500 59562 139512
rect 71090 139500 71096 139512
rect 59556 139472 71096 139500
rect 59556 139460 59562 139472
rect 71090 139460 71096 139472
rect 71148 139460 71154 139512
rect 77533 139503 77591 139509
rect 77533 139469 77545 139503
rect 77579 139500 77591 139503
rect 87101 139503 87159 139509
rect 87101 139500 87113 139503
rect 77579 139472 87113 139500
rect 77579 139469 77591 139472
rect 77533 139463 77591 139469
rect 87101 139469 87113 139472
rect 87147 139469 87159 139503
rect 116170 139500 116176 139512
rect 87101 139463 87159 139469
rect 109472 139472 116176 139500
rect 56738 139392 56744 139444
rect 56796 139432 56802 139444
rect 67962 139432 67968 139444
rect 56796 139404 67968 139432
rect 56796 139392 56802 139404
rect 67962 139392 67968 139404
rect 68020 139392 68026 139444
rect 109273 139435 109331 139441
rect 109273 139401 109285 139435
rect 109319 139432 109331 139435
rect 109472 139432 109500 139472
rect 116170 139460 116176 139472
rect 116228 139500 116234 139512
rect 118473 139503 118531 139509
rect 118473 139500 118485 139503
rect 116228 139472 118485 139500
rect 116228 139460 116234 139472
rect 118473 139469 118485 139472
rect 118519 139469 118531 139503
rect 118473 139463 118531 139469
rect 154718 139460 154724 139512
rect 154776 139500 154782 139512
rect 167322 139500 167328 139512
rect 154776 139472 167328 139500
rect 154776 139460 154782 139472
rect 167322 139460 167328 139472
rect 167380 139460 167386 139512
rect 109319 139404 109500 139432
rect 109319 139401 109331 139404
rect 109273 139395 109331 139401
rect 151866 139392 151872 139444
rect 151924 139432 151930 139444
rect 158033 139435 158091 139441
rect 158033 139432 158045 139435
rect 151924 139404 158045 139432
rect 151924 139392 151930 139404
rect 158033 139401 158045 139404
rect 158079 139401 158091 139435
rect 158033 139395 158091 139401
rect 158122 139392 158128 139444
rect 158180 139432 158186 139444
rect 160790 139432 160796 139444
rect 158180 139404 160796 139432
rect 158180 139392 158186 139404
rect 160790 139392 160796 139404
rect 160848 139392 160854 139444
rect 160882 139392 160888 139444
rect 160940 139432 160946 139444
rect 163458 139432 163464 139444
rect 160940 139404 163464 139432
rect 160940 139392 160946 139404
rect 163458 139392 163464 139404
rect 163516 139392 163522 139444
rect 251318 139392 251324 139444
rect 251376 139432 251382 139444
rect 253176 139432 253204 139608
rect 264106 139596 264112 139608
rect 264164 139596 264170 139648
rect 263094 139568 263100 139580
rect 251376 139404 253204 139432
rect 253268 139540 263100 139568
rect 251376 139392 251382 139404
rect 58118 139324 58124 139376
rect 58176 139364 58182 139376
rect 70078 139364 70084 139376
rect 58176 139336 70084 139364
rect 58176 139324 58182 139336
rect 70078 139324 70084 139336
rect 70136 139324 70142 139376
rect 75138 139324 75144 139376
rect 75196 139364 75202 139376
rect 77533 139367 77591 139373
rect 77533 139364 77545 139367
rect 75196 139336 77545 139364
rect 75196 139324 75202 139336
rect 77533 139333 77545 139336
rect 77579 139333 77591 139367
rect 109181 139367 109239 139373
rect 109181 139364 109193 139367
rect 77533 139327 77591 139333
rect 89968 139336 109193 139364
rect 55358 139256 55364 139308
rect 55416 139296 55422 139308
rect 66950 139296 66956 139308
rect 55416 139268 66956 139296
rect 55416 139256 55422 139268
rect 66950 139256 66956 139268
rect 67008 139256 67014 139308
rect 87101 139299 87159 139305
rect 87101 139265 87113 139299
rect 87147 139296 87159 139299
rect 89968 139296 89996 139336
rect 109181 139333 109193 139336
rect 109227 139333 109239 139367
rect 109181 139327 109239 139333
rect 124453 139367 124511 139373
rect 124453 139333 124465 139367
rect 124499 139364 124511 139367
rect 134113 139367 134171 139373
rect 134113 139364 134125 139367
rect 124499 139336 134125 139364
rect 124499 139333 124511 139336
rect 124453 139327 124511 139333
rect 134113 139333 134125 139336
rect 134159 139333 134171 139367
rect 134113 139327 134171 139333
rect 150486 139324 150492 139376
rect 150544 139364 150550 139376
rect 163274 139364 163280 139376
rect 150544 139336 163280 139364
rect 150544 139324 150550 139336
rect 163274 139324 163280 139336
rect 163332 139324 163338 139376
rect 249938 139324 249944 139376
rect 249996 139364 250002 139376
rect 253268 139364 253296 139540
rect 263094 139528 263100 139540
rect 263152 139528 263158 139580
rect 254081 139503 254139 139509
rect 254081 139469 254093 139503
rect 254127 139500 254139 139503
rect 261254 139500 261260 139512
rect 254127 139472 261260 139500
rect 254127 139469 254139 139472
rect 254081 139463 254139 139469
rect 261254 139460 261260 139472
rect 261312 139460 261318 139512
rect 253345 139435 253403 139441
rect 253345 139401 253357 139435
rect 253391 139432 253403 139435
rect 260150 139432 260156 139444
rect 253391 139404 260156 139432
rect 253391 139401 253403 139404
rect 253345 139395 253403 139401
rect 260150 139392 260156 139404
rect 260208 139392 260214 139444
rect 249996 139336 253296 139364
rect 253437 139367 253495 139373
rect 249996 139324 250002 139336
rect 253437 139333 253449 139367
rect 253483 139364 253495 139367
rect 258310 139364 258316 139376
rect 253483 139336 258316 139364
rect 253483 139333 253495 139336
rect 253437 139327 253495 139333
rect 258310 139324 258316 139336
rect 258368 139324 258374 139376
rect 87147 139268 89996 139296
rect 87147 139265 87159 139268
rect 87101 139259 87159 139265
rect 154626 139256 154632 139308
rect 154684 139296 154690 139308
rect 168058 139296 168064 139308
rect 154684 139268 168064 139296
rect 154684 139256 154690 139268
rect 168058 139256 168064 139268
rect 168116 139256 168122 139308
rect 244418 139256 244424 139308
rect 244476 139296 244482 139308
rect 257298 139296 257304 139308
rect 244476 139268 257304 139296
rect 244476 139256 244482 139268
rect 257298 139256 257304 139268
rect 257356 139256 257362 139308
rect 60786 139188 60792 139240
rect 60844 139228 60850 139240
rect 72102 139228 72108 139240
rect 60844 139200 72108 139228
rect 60844 139188 60850 139200
rect 72102 139188 72108 139200
rect 72160 139188 72166 139240
rect 144598 139188 144604 139240
rect 144656 139228 144662 139240
rect 170726 139228 170732 139240
rect 144656 139200 170732 139228
rect 144656 139188 144662 139200
rect 170726 139188 170732 139200
rect 170784 139188 170790 139240
rect 238622 139188 238628 139240
rect 238680 139228 238686 139240
rect 264474 139228 264480 139240
rect 238680 139200 264480 139228
rect 238680 139188 238686 139200
rect 264474 139188 264480 139200
rect 264532 139188 264538 139240
rect 333382 139188 333388 139240
rect 333440 139228 333446 139240
rect 334118 139228 334124 139240
rect 333440 139200 334124 139228
rect 333440 139188 333446 139200
rect 334118 139188 334124 139200
rect 334176 139188 334182 139240
rect 118473 139163 118531 139169
rect 118473 139129 118485 139163
rect 118519 139160 118531 139163
rect 124453 139163 124511 139169
rect 124453 139160 124465 139163
rect 118519 139132 124465 139160
rect 118519 139129 118531 139132
rect 118473 139123 118531 139129
rect 124453 139129 124465 139132
rect 124499 139129 124511 139163
rect 124453 139123 124511 139129
rect 143681 139163 143739 139169
rect 143681 139129 143693 139163
rect 143727 139160 143739 139163
rect 152694 139160 152700 139172
rect 143727 139132 152700 139160
rect 143727 139129 143739 139132
rect 143681 139123 143739 139129
rect 152694 139120 152700 139132
rect 152752 139120 152758 139172
rect 153338 139120 153344 139172
rect 153396 139160 153402 139172
rect 158033 139163 158091 139169
rect 153396 139132 157984 139160
rect 153396 139120 153402 139132
rect 63822 139052 63828 139104
rect 63880 139092 63886 139104
rect 68606 139092 68612 139104
rect 63880 139064 68612 139092
rect 63880 139052 63886 139064
rect 68606 139052 68612 139064
rect 68664 139052 68670 139104
rect 134113 139027 134171 139033
rect 134113 138993 134125 139027
rect 134159 139024 134171 139027
rect 136870 139024 136876 139036
rect 134159 138996 136876 139024
rect 134159 138993 134171 138996
rect 134113 138987 134171 138993
rect 136870 138984 136876 138996
rect 136928 139024 136934 139036
rect 143681 139027 143739 139033
rect 143681 139024 143693 139027
rect 136928 138996 143693 139024
rect 136928 138984 136934 138996
rect 143681 138993 143693 138996
rect 143727 138993 143739 139027
rect 157956 139024 157984 139132
rect 158033 139129 158045 139163
rect 158079 139160 158091 139163
rect 165206 139160 165212 139172
rect 158079 139132 165212 139160
rect 158079 139129 158091 139132
rect 158033 139123 158091 139129
rect 165206 139120 165212 139132
rect 165264 139120 165270 139172
rect 249846 139120 249852 139172
rect 249904 139160 249910 139172
rect 262082 139160 262088 139172
rect 249904 139132 262088 139160
rect 249904 139120 249910 139132
rect 262082 139120 262088 139132
rect 262140 139120 262146 139172
rect 248558 139052 248564 139104
rect 248616 139092 248622 139104
rect 253989 139095 254047 139101
rect 253989 139092 254001 139095
rect 248616 139064 254001 139092
rect 248616 139052 248622 139064
rect 253989 139061 254001 139064
rect 254035 139061 254047 139095
rect 253989 139055 254047 139061
rect 166126 139024 166132 139036
rect 157956 138996 166132 139024
rect 143681 138987 143739 138993
rect 166126 138984 166132 138996
rect 166184 138984 166190 139036
rect 247178 138984 247184 139036
rect 247236 139024 247242 139036
rect 253345 139027 253403 139033
rect 253345 139024 253357 139027
rect 247236 138996 253357 139024
rect 247236 138984 247242 138996
rect 253345 138993 253357 138996
rect 253391 138993 253403 139027
rect 253345 138987 253403 138993
rect 58670 138916 58676 138968
rect 58728 138956 58734 138968
rect 62994 138956 63000 138968
rect 58728 138928 63000 138956
rect 58728 138916 58734 138928
rect 62994 138916 63000 138928
rect 63052 138916 63058 138968
rect 64374 138916 64380 138968
rect 64432 138956 64438 138968
rect 68974 138956 68980 138968
rect 64432 138928 68980 138956
rect 64432 138916 64438 138928
rect 68974 138916 68980 138928
rect 69032 138916 69038 138968
rect 157570 138916 157576 138968
rect 157628 138956 157634 138968
rect 158214 138956 158220 138968
rect 157628 138928 158220 138956
rect 157628 138916 157634 138928
rect 158214 138916 158220 138928
rect 158272 138916 158278 138968
rect 245798 138916 245804 138968
rect 245856 138956 245862 138968
rect 253437 138959 253495 138965
rect 253437 138956 253449 138959
rect 245856 138928 253449 138956
rect 245856 138916 245862 138928
rect 253437 138925 253449 138928
rect 253483 138925 253495 138959
rect 253437 138919 253495 138925
rect 62810 138848 62816 138900
rect 62868 138888 62874 138900
rect 67686 138888 67692 138900
rect 62868 138860 67692 138888
rect 62868 138848 62874 138860
rect 67686 138848 67692 138860
rect 67744 138848 67750 138900
rect 157110 138848 157116 138900
rect 157168 138888 157174 138900
rect 159962 138888 159968 138900
rect 157168 138860 159968 138888
rect 157168 138848 157174 138860
rect 159962 138848 159968 138860
rect 160020 138848 160026 138900
rect 244970 138848 244976 138900
rect 245028 138888 245034 138900
rect 252238 138888 252244 138900
rect 245028 138860 252244 138888
rect 245028 138848 245034 138860
rect 252238 138848 252244 138860
rect 252296 138848 252302 138900
rect 341754 138848 341760 138900
rect 341812 138888 341818 138900
rect 341812 138860 342812 138888
rect 341812 138848 341818 138860
rect 59682 138780 59688 138832
rect 59740 138820 59746 138832
rect 63086 138820 63092 138832
rect 59740 138792 63092 138820
rect 59740 138780 59746 138792
rect 63086 138780 63092 138792
rect 63144 138780 63150 138832
rect 157573 138823 157631 138829
rect 157573 138789 157585 138823
rect 157619 138820 157631 138823
rect 162725 138823 162783 138829
rect 162725 138820 162737 138823
rect 157619 138792 162737 138820
rect 157619 138789 157631 138792
rect 157573 138783 157631 138789
rect 162725 138789 162737 138792
rect 162771 138789 162783 138823
rect 162725 138783 162783 138789
rect 242486 138780 242492 138832
rect 242544 138820 242550 138832
rect 249110 138820 249116 138832
rect 242544 138792 249116 138820
rect 242544 138780 242550 138792
rect 249110 138780 249116 138792
rect 249168 138780 249174 138832
rect 253894 138780 253900 138832
rect 253952 138820 253958 138832
rect 256654 138820 256660 138832
rect 253952 138792 256660 138820
rect 253952 138780 253958 138792
rect 256654 138780 256660 138792
rect 256712 138780 256718 138832
rect 338258 138780 338264 138832
rect 338316 138820 338322 138832
rect 342674 138820 342680 138832
rect 338316 138792 342680 138820
rect 338316 138780 338322 138792
rect 342674 138780 342680 138792
rect 342732 138780 342738 138832
rect 342784 138820 342812 138860
rect 345802 138820 345808 138832
rect 342784 138792 345808 138820
rect 345802 138780 345808 138792
rect 345860 138780 345866 138832
rect 61798 138712 61804 138764
rect 61856 138752 61862 138764
rect 65754 138752 65760 138764
rect 61856 138724 65760 138752
rect 61856 138712 61862 138724
rect 65754 138712 65760 138724
rect 65812 138712 65818 138764
rect 145242 138712 145248 138764
rect 145300 138752 145306 138764
rect 365214 138752 365220 138764
rect 145300 138724 365220 138752
rect 145300 138712 145306 138724
rect 365214 138712 365220 138724
rect 365272 138712 365278 138764
rect 60694 138644 60700 138696
rect 60752 138684 60758 138696
rect 63178 138684 63184 138696
rect 60752 138656 63184 138684
rect 60752 138644 60758 138656
rect 63178 138644 63184 138656
rect 63236 138644 63242 138696
rect 252146 138644 252152 138696
rect 252204 138684 252210 138696
rect 254170 138684 254176 138696
rect 252204 138656 254176 138684
rect 252204 138644 252210 138656
rect 254170 138644 254176 138656
rect 254228 138644 254234 138696
rect 256010 138644 256016 138696
rect 256068 138684 256074 138696
rect 258678 138684 258684 138696
rect 256068 138656 258684 138684
rect 256068 138644 256074 138656
rect 258678 138644 258684 138656
rect 258736 138644 258742 138696
rect 338166 138644 338172 138696
rect 338224 138684 338230 138696
rect 341662 138684 341668 138696
rect 338224 138656 341668 138684
rect 338224 138644 338230 138656
rect 341662 138644 341668 138656
rect 341720 138644 341726 138696
rect 341938 138644 341944 138696
rect 341996 138684 342002 138696
rect 344790 138684 344796 138696
rect 341996 138656 344796 138684
rect 341996 138644 342002 138656
rect 344790 138644 344796 138656
rect 344848 138644 344854 138696
rect 57658 138576 57664 138628
rect 57716 138616 57722 138628
rect 61614 138616 61620 138628
rect 57716 138588 61620 138616
rect 57716 138576 57722 138588
rect 61614 138576 61620 138588
rect 61672 138576 61678 138628
rect 65938 138576 65944 138628
rect 65996 138616 66002 138628
rect 70538 138616 70544 138628
rect 65996 138588 70544 138616
rect 65996 138576 66002 138588
rect 70538 138576 70544 138588
rect 70596 138576 70602 138628
rect 155178 138576 155184 138628
rect 155236 138616 155242 138628
rect 158030 138616 158036 138628
rect 155236 138588 158036 138616
rect 155236 138576 155242 138588
rect 158030 138576 158036 138588
rect 158088 138576 158094 138628
rect 252698 138576 252704 138628
rect 252756 138616 252762 138628
rect 254814 138616 254820 138628
rect 252756 138588 254820 138616
rect 252756 138576 252762 138588
rect 254814 138576 254820 138588
rect 254872 138576 254878 138628
rect 254998 138576 255004 138628
rect 255056 138616 255062 138628
rect 257482 138616 257488 138628
rect 255056 138588 257488 138616
rect 255056 138576 255062 138588
rect 257482 138576 257488 138588
rect 257540 138576 257546 138628
rect 334394 138576 334400 138628
rect 334452 138616 334458 138628
rect 335498 138616 335504 138628
rect 334452 138588 335504 138616
rect 334452 138576 334458 138588
rect 335498 138576 335504 138588
rect 335556 138576 335562 138628
rect 338534 138576 338540 138628
rect 338592 138616 338598 138628
rect 339638 138616 339644 138628
rect 338592 138588 339644 138616
rect 338592 138576 338598 138588
rect 339638 138576 339644 138588
rect 339696 138576 339702 138628
rect 341846 138576 341852 138628
rect 341904 138616 341910 138628
rect 343778 138616 343784 138628
rect 341904 138588 343784 138616
rect 341904 138576 341910 138588
rect 343778 138576 343784 138588
rect 343836 138576 343842 138628
rect 348654 138576 348660 138628
rect 348712 138616 348718 138628
rect 349942 138616 349948 138628
rect 348712 138588 349948 138616
rect 348712 138576 348718 138588
rect 349942 138576 349948 138588
rect 350000 138576 350006 138628
rect 284438 137828 284444 137880
rect 284496 137868 284502 137880
rect 324826 137868 324832 137880
rect 284496 137840 324832 137868
rect 284496 137828 284502 137840
rect 324826 137828 324832 137840
rect 324884 137828 324890 137880
rect 12854 137080 12860 137132
rect 12912 137120 12918 137132
rect 16074 137120 16080 137132
rect 12912 137092 16080 137120
rect 12912 137080 12918 137092
rect 16074 137080 16080 137092
rect 16132 137080 16138 137132
rect 137146 137080 137152 137132
rect 137204 137120 137210 137132
rect 137422 137120 137428 137132
rect 137204 137092 137428 137120
rect 137204 137080 137210 137092
rect 137422 137080 137428 137092
rect 137480 137080 137486 137132
rect 210010 136672 210016 136724
rect 210068 136712 210074 136724
rect 218934 136712 218940 136724
rect 210068 136684 218940 136712
rect 210068 136672 210074 136684
rect 218934 136672 218940 136684
rect 218992 136672 218998 136724
rect 346630 136468 346636 136520
rect 346688 136508 346694 136520
rect 347550 136508 347556 136520
rect 346688 136480 347556 136508
rect 346688 136468 346694 136480
rect 347550 136468 347556 136480
rect 347608 136468 347614 136520
rect 304034 136400 304040 136452
rect 304092 136440 304098 136452
rect 312774 136440 312780 136452
rect 304092 136412 312780 136440
rect 304092 136400 304098 136412
rect 312774 136400 312780 136412
rect 312832 136400 312838 136452
rect 291522 136264 291528 136316
rect 291580 136304 291586 136316
rect 292718 136304 292724 136316
rect 291580 136276 292724 136304
rect 291580 136264 291586 136276
rect 292718 136264 292724 136276
rect 292776 136264 292782 136316
rect 279102 136128 279108 136180
rect 279160 136168 279166 136180
rect 280298 136168 280304 136180
rect 279160 136140 280304 136168
rect 279160 136128 279166 136140
rect 280298 136128 280304 136140
rect 280356 136128 280362 136180
rect 324550 135788 324556 135840
rect 324608 135828 324614 135840
rect 346998 135828 347004 135840
rect 324608 135800 347004 135828
rect 324608 135788 324614 135800
rect 346998 135788 347004 135800
rect 347056 135828 347062 135840
rect 347056 135800 347964 135828
rect 347056 135788 347062 135800
rect 347936 135760 347964 135800
rect 359050 135760 359056 135772
rect 347936 135732 359056 135760
rect 359050 135720 359056 135732
rect 359108 135720 359114 135772
rect 286738 135040 286744 135092
rect 286796 135080 286802 135092
rect 324642 135080 324648 135092
rect 286796 135052 324648 135080
rect 286796 135040 286802 135052
rect 324642 135040 324648 135052
rect 324700 135040 324706 135092
rect 343870 135040 343876 135092
rect 343928 135080 343934 135092
rect 360798 135080 360804 135092
rect 343928 135052 360804 135080
rect 343928 135040 343934 135052
rect 360798 135040 360804 135052
rect 360856 135040 360862 135092
rect 324642 134428 324648 134480
rect 324700 134468 324706 134480
rect 343870 134468 343876 134480
rect 324700 134440 343876 134468
rect 324700 134428 324706 134440
rect 343870 134428 343876 134440
rect 343928 134428 343934 134480
rect 51494 134360 51500 134412
rect 51552 134400 51558 134412
rect 51586 134400 51592 134412
rect 51552 134372 51592 134400
rect 51552 134360 51558 134372
rect 51586 134360 51592 134372
rect 51644 134360 51650 134412
rect 343962 133680 343968 133732
rect 344020 133720 344026 133732
rect 360706 133720 360712 133732
rect 344020 133692 360712 133720
rect 344020 133680 344026 133692
rect 360706 133680 360712 133692
rect 360764 133680 360770 133732
rect 326574 133000 326580 133052
rect 326632 133040 326638 133052
rect 343962 133040 343968 133052
rect 326632 133012 343968 133040
rect 326632 133000 326638 133012
rect 343962 133000 343968 133012
rect 344020 133040 344026 133052
rect 344238 133040 344244 133052
rect 344020 133012 344244 133040
rect 344020 133000 344026 133012
rect 344238 133000 344244 133012
rect 344296 133000 344302 133052
rect 346078 132456 346084 132508
rect 346136 132496 346142 132508
rect 360430 132496 360436 132508
rect 346136 132468 360436 132496
rect 346136 132456 346142 132468
rect 360430 132456 360436 132468
rect 360488 132456 360494 132508
rect 354910 132388 354916 132440
rect 354968 132428 354974 132440
rect 355830 132428 355836 132440
rect 354968 132400 355836 132428
rect 354968 132388 354974 132400
rect 355830 132388 355836 132400
rect 355888 132388 355894 132440
rect 136870 132320 136876 132372
rect 136928 132360 136934 132372
rect 137330 132360 137336 132372
rect 136928 132332 137336 132360
rect 136928 132320 136934 132332
rect 137330 132320 137336 132332
rect 137388 132320 137394 132372
rect 343318 132320 343324 132372
rect 343376 132360 343382 132372
rect 360982 132360 360988 132372
rect 343376 132332 360988 132360
rect 343376 132320 343382 132332
rect 360982 132320 360988 132332
rect 361040 132320 361046 132372
rect 258954 132252 258960 132304
rect 259012 132292 259018 132304
rect 368894 132292 368900 132304
rect 259012 132264 368900 132292
rect 259012 132252 259018 132264
rect 368894 132252 368900 132264
rect 368952 132252 368958 132304
rect 324550 132184 324556 132236
rect 324608 132224 324614 132236
rect 324734 132224 324740 132236
rect 324608 132196 324740 132224
rect 324608 132184 324614 132196
rect 324734 132184 324740 132196
rect 324792 132184 324798 132236
rect 324826 131708 324832 131760
rect 324884 131748 324890 131760
rect 325470 131748 325476 131760
rect 324884 131720 325476 131748
rect 324884 131708 324890 131720
rect 325470 131708 325476 131720
rect 325528 131748 325534 131760
rect 343318 131748 343324 131760
rect 325528 131720 343324 131748
rect 325528 131708 325534 131720
rect 343318 131708 343324 131720
rect 343376 131708 343382 131760
rect 325102 131640 325108 131692
rect 325160 131680 325166 131692
rect 346078 131680 346084 131692
rect 325160 131652 346084 131680
rect 325160 131640 325166 131652
rect 346078 131640 346084 131652
rect 346136 131640 346142 131692
rect 56094 131572 56100 131624
rect 56152 131612 56158 131624
rect 56738 131612 56744 131624
rect 56152 131584 56744 131612
rect 56152 131572 56158 131584
rect 56738 131572 56744 131584
rect 56796 131572 56802 131624
rect 59682 131572 59688 131624
rect 59740 131612 59746 131624
rect 60786 131612 60792 131624
rect 59740 131584 60792 131612
rect 59740 131572 59746 131584
rect 60786 131572 60792 131584
rect 60844 131572 60850 131624
rect 155454 131572 155460 131624
rect 155512 131612 155518 131624
rect 156098 131612 156104 131624
rect 155512 131584 156104 131612
rect 155512 131572 155518 131584
rect 156098 131572 156104 131584
rect 156156 131572 156162 131624
rect 245338 131572 245344 131624
rect 245396 131612 245402 131624
rect 245798 131612 245804 131624
rect 245396 131584 245804 131612
rect 245396 131572 245402 131584
rect 245798 131572 245804 131584
rect 245856 131572 245862 131624
rect 248006 131572 248012 131624
rect 248064 131612 248070 131624
rect 248558 131612 248564 131624
rect 248064 131584 248564 131612
rect 248064 131572 248070 131584
rect 248558 131572 248564 131584
rect 248616 131572 248622 131624
rect 341662 131572 341668 131624
rect 341720 131612 341726 131624
rect 348010 131612 348016 131624
rect 341720 131584 348016 131612
rect 341720 131572 341726 131584
rect 348010 131572 348016 131584
rect 348068 131572 348074 131624
rect 339638 131504 339644 131556
rect 339696 131544 339702 131556
rect 350954 131544 350960 131556
rect 339696 131516 350960 131544
rect 339696 131504 339702 131516
rect 350954 131504 350960 131516
rect 351012 131504 351018 131556
rect 160974 131436 160980 131488
rect 161032 131476 161038 131488
rect 161710 131476 161716 131488
rect 161032 131448 161716 131476
rect 161032 131436 161038 131448
rect 161710 131436 161716 131448
rect 161768 131436 161774 131488
rect 341018 131436 341024 131488
rect 341076 131476 341082 131488
rect 352242 131476 352248 131488
rect 341076 131448 352248 131476
rect 341076 131436 341082 131448
rect 352242 131436 352248 131448
rect 352300 131436 352306 131488
rect 339546 131368 339552 131420
rect 339604 131408 339610 131420
rect 351598 131408 351604 131420
rect 339604 131380 351604 131408
rect 339604 131368 339610 131380
rect 351598 131368 351604 131380
rect 351656 131368 351662 131420
rect 338074 131300 338080 131352
rect 338132 131340 338138 131352
rect 350402 131340 350408 131352
rect 338132 131312 350408 131340
rect 338132 131300 338138 131312
rect 350402 131300 350408 131312
rect 350460 131300 350466 131352
rect 231354 131232 231360 131284
rect 231412 131272 231418 131284
rect 322618 131272 322624 131284
rect 231412 131244 322624 131272
rect 231412 131232 231418 131244
rect 322618 131232 322624 131244
rect 322676 131232 322682 131284
rect 335498 131232 335504 131284
rect 335556 131272 335562 131284
rect 348562 131272 348568 131284
rect 335556 131244 348568 131272
rect 335556 131232 335562 131244
rect 348562 131232 348568 131244
rect 348620 131232 348626 131284
rect 248466 131164 248472 131216
rect 248524 131204 248530 131216
rect 250950 131204 250956 131216
rect 248524 131176 250956 131204
rect 248524 131164 248530 131176
rect 250950 131164 250956 131176
rect 251008 131164 251014 131216
rect 336878 131164 336884 131216
rect 336936 131204 336942 131216
rect 349758 131204 349764 131216
rect 336936 131176 349764 131204
rect 336936 131164 336942 131176
rect 349758 131164 349764 131176
rect 349816 131164 349822 131216
rect 332738 131096 332744 131148
rect 332796 131136 332802 131148
rect 336789 131139 336847 131145
rect 336789 131136 336801 131139
rect 332796 131108 336801 131136
rect 332796 131096 332802 131108
rect 336789 131105 336801 131108
rect 336835 131105 336847 131139
rect 336789 131099 336847 131105
rect 341018 131096 341024 131148
rect 341076 131136 341082 131148
rect 346630 131136 346636 131148
rect 341076 131108 346636 131136
rect 341076 131096 341082 131108
rect 346630 131096 346636 131108
rect 346688 131096 346694 131148
rect 334118 131028 334124 131080
rect 334176 131068 334182 131080
rect 348010 131068 348016 131080
rect 334176 131040 348016 131068
rect 334176 131028 334182 131040
rect 348010 131028 348016 131040
rect 348068 131028 348074 131080
rect 335406 130960 335412 131012
rect 335464 131000 335470 131012
rect 349390 131000 349396 131012
rect 335464 130972 349396 131000
rect 335464 130960 335470 130972
rect 349390 130960 349396 130972
rect 349448 130960 349454 131012
rect 340558 130892 340564 130944
rect 340616 130932 340622 130944
rect 346722 130932 346728 130944
rect 340616 130904 346728 130932
rect 340616 130892 340622 130904
rect 346722 130892 346728 130904
rect 346780 130892 346786 130944
rect 360890 130932 360896 130944
rect 348764 130904 360896 130932
rect 342490 130864 342496 130876
rect 336712 130836 342496 130864
rect 63178 130688 63184 130740
rect 63236 130728 63242 130740
rect 65938 130728 65944 130740
rect 63236 130700 65944 130728
rect 63236 130688 63242 130700
rect 65938 130688 65944 130700
rect 65996 130688 66002 130740
rect 243590 130688 243596 130740
rect 243648 130728 243654 130740
rect 244326 130728 244332 130740
rect 243648 130700 244332 130728
rect 243648 130688 243654 130700
rect 244326 130688 244332 130700
rect 244384 130688 244390 130740
rect 250674 130688 250680 130740
rect 250732 130728 250738 130740
rect 251318 130728 251324 130740
rect 250732 130700 251324 130728
rect 250732 130688 250738 130700
rect 251318 130688 251324 130700
rect 251376 130688 251382 130740
rect 57014 130552 57020 130604
rect 57072 130592 57078 130604
rect 64374 130592 64380 130604
rect 57072 130564 64380 130592
rect 57072 130552 57078 130564
rect 64374 130552 64380 130564
rect 64432 130552 64438 130604
rect 63086 130484 63092 130536
rect 63144 130524 63150 130536
rect 65018 130524 65024 130536
rect 63144 130496 65024 130524
rect 63144 130484 63150 130496
rect 65018 130484 65024 130496
rect 65076 130484 65082 130536
rect 61614 130416 61620 130468
rect 61672 130456 61678 130468
rect 63270 130456 63276 130468
rect 61672 130428 63276 130456
rect 61672 130416 61678 130428
rect 63270 130416 63276 130428
rect 63328 130416 63334 130468
rect 246258 130416 246264 130468
rect 246316 130456 246322 130468
rect 247086 130456 247092 130468
rect 246316 130428 247092 130456
rect 246316 130416 246322 130428
rect 247086 130416 247092 130428
rect 247144 130416 247150 130468
rect 248926 130416 248932 130468
rect 248984 130456 248990 130468
rect 249846 130456 249852 130468
rect 248984 130428 249852 130456
rect 248984 130416 248990 130428
rect 249846 130416 249852 130428
rect 249904 130416 249910 130468
rect 325378 130416 325384 130468
rect 325436 130456 325442 130468
rect 336712 130456 336740 130836
rect 342490 130824 342496 130836
rect 342548 130864 342554 130876
rect 345253 130867 345311 130873
rect 345253 130864 345265 130867
rect 342548 130836 345265 130864
rect 342548 130824 342554 130836
rect 345253 130833 345265 130836
rect 345299 130833 345311 130867
rect 345253 130827 345311 130833
rect 342398 130756 342404 130808
rect 342456 130796 342462 130808
rect 348654 130796 348660 130808
rect 342456 130768 348660 130796
rect 342456 130756 342462 130768
rect 348654 130756 348660 130768
rect 348712 130756 348718 130808
rect 336789 130731 336847 130737
rect 336789 130697 336801 130731
rect 336835 130728 336847 130731
rect 347274 130728 347280 130740
rect 336835 130700 347280 130728
rect 336835 130697 336847 130700
rect 336789 130691 336847 130697
rect 347274 130688 347280 130700
rect 347332 130688 347338 130740
rect 345345 130663 345403 130669
rect 325436 130428 336740 130456
rect 337356 130632 345296 130660
rect 325436 130416 325442 130428
rect 62350 130348 62356 130400
rect 62408 130388 62414 130400
rect 63638 130388 63644 130400
rect 62408 130360 63644 130388
rect 62408 130348 62414 130360
rect 63638 130348 63644 130360
rect 63696 130348 63702 130400
rect 324734 130348 324740 130400
rect 324792 130388 324798 130400
rect 325286 130388 325292 130400
rect 324792 130360 325292 130388
rect 324792 130348 324798 130360
rect 325286 130348 325292 130360
rect 325344 130388 325350 130400
rect 337356 130388 337384 130632
rect 338718 130552 338724 130604
rect 338776 130592 338782 130604
rect 341846 130592 341852 130604
rect 338776 130564 341852 130592
rect 338776 130552 338782 130564
rect 341846 130552 341852 130564
rect 341904 130552 341910 130604
rect 339362 130484 339368 130536
rect 339420 130524 339426 130536
rect 341938 130524 341944 130536
rect 339420 130496 341944 130524
rect 339420 130484 339426 130496
rect 341938 130484 341944 130496
rect 341996 130484 342002 130536
rect 345158 130524 345164 130536
rect 345117 130496 345164 130524
rect 345158 130484 345164 130496
rect 345216 130524 345222 130536
rect 345268 130524 345296 130632
rect 345345 130629 345357 130663
rect 345391 130660 345403 130663
rect 348764 130660 348792 130904
rect 360890 130892 360896 130904
rect 360948 130892 360954 130944
rect 345391 130632 348792 130660
rect 345391 130629 345403 130632
rect 345345 130623 345403 130629
rect 345216 130496 345296 130524
rect 345216 130484 345250 130496
rect 345222 130456 345250 130484
rect 360338 130456 360344 130468
rect 345222 130428 360344 130456
rect 360338 130416 360344 130428
rect 360396 130416 360402 130468
rect 360522 130416 360528 130468
rect 360580 130416 360586 130468
rect 325344 130360 337384 130388
rect 325344 130348 325350 130360
rect 337522 130348 337528 130400
rect 337580 130388 337586 130400
rect 338166 130388 338172 130400
rect 337580 130360 338172 130388
rect 337580 130348 337586 130360
rect 338166 130348 338172 130360
rect 338224 130348 338230 130400
rect 339546 130348 339552 130400
rect 339604 130388 339610 130400
rect 341754 130388 341760 130400
rect 339604 130360 341760 130388
rect 339604 130348 339610 130360
rect 341754 130348 341760 130360
rect 341812 130348 341818 130400
rect 61430 130280 61436 130332
rect 61488 130320 61494 130332
rect 62258 130320 62264 130332
rect 61488 130292 62264 130320
rect 61488 130280 61494 130292
rect 62258 130280 62264 130292
rect 62316 130280 62322 130332
rect 62994 130280 63000 130332
rect 63052 130320 63058 130332
rect 64098 130320 64104 130332
rect 63052 130292 64104 130320
rect 63052 130280 63058 130292
rect 64098 130280 64104 130292
rect 64156 130280 64162 130332
rect 65754 130280 65760 130332
rect 65812 130320 65818 130332
rect 66766 130320 66772 130332
rect 65812 130292 66772 130320
rect 65812 130280 65818 130292
rect 66766 130280 66772 130292
rect 66824 130280 66830 130332
rect 149290 130280 149296 130332
rect 149348 130320 149354 130332
rect 150578 130320 150584 130332
rect 149348 130292 150584 130320
rect 149348 130280 149354 130292
rect 150578 130280 150584 130292
rect 150636 130280 150642 130332
rect 151038 130280 151044 130332
rect 151096 130320 151102 130332
rect 151774 130320 151780 130332
rect 151096 130292 151780 130320
rect 151096 130280 151102 130292
rect 151774 130280 151780 130292
rect 151832 130280 151838 130332
rect 153706 130280 153712 130332
rect 153764 130320 153770 130332
rect 154718 130320 154724 130332
rect 153764 130292 154724 130320
rect 153764 130280 153770 130292
rect 154718 130280 154724 130292
rect 154776 130280 154782 130332
rect 156374 130280 156380 130332
rect 156432 130320 156438 130332
rect 157478 130320 157484 130332
rect 156432 130292 157484 130320
rect 156432 130280 156438 130292
rect 157478 130280 157484 130292
rect 157536 130280 157542 130332
rect 158214 130280 158220 130332
rect 158272 130320 158278 130332
rect 159042 130320 159048 130332
rect 158272 130292 159048 130320
rect 158272 130280 158278 130292
rect 159042 130280 159048 130292
rect 159100 130280 159106 130332
rect 162998 130280 163004 130332
rect 163056 130320 163062 130332
rect 164378 130320 164384 130332
rect 163056 130292 164384 130320
rect 163056 130280 163062 130292
rect 164378 130280 164384 130292
rect 164436 130280 164442 130332
rect 254814 130280 254820 130332
rect 254872 130320 254878 130332
rect 255550 130320 255556 130332
rect 254872 130292 255556 130320
rect 254872 130280 254878 130292
rect 255550 130280 255556 130292
rect 255608 130280 255614 130332
rect 324642 130280 324648 130332
rect 324700 130320 324706 130332
rect 345710 130320 345716 130332
rect 324700 130292 345716 130320
rect 324700 130280 324706 130292
rect 345710 130280 345716 130292
rect 345768 130320 345774 130332
rect 360540 130320 360568 130416
rect 361074 130320 361080 130332
rect 345768 130292 361080 130320
rect 345768 130280 345774 130292
rect 361074 130280 361080 130292
rect 361132 130280 361138 130332
rect 231078 130212 231084 130264
rect 231136 130252 231142 130264
rect 246442 130252 246448 130264
rect 231136 130224 246448 130252
rect 231136 130212 231142 130224
rect 246442 130212 246448 130224
rect 246500 130212 246506 130264
rect 137054 127492 137060 127544
rect 137112 127532 137118 127544
rect 137422 127532 137428 127544
rect 137112 127504 137428 127532
rect 137112 127492 137118 127504
rect 137422 127492 137428 127504
rect 137480 127492 137486 127544
rect 84706 127424 84712 127476
rect 84764 127464 84770 127476
rect 85810 127464 85816 127476
rect 84764 127436 85816 127464
rect 84764 127424 84770 127436
rect 85810 127424 85816 127436
rect 85868 127424 85874 127476
rect 38798 126744 38804 126796
rect 38856 126784 38862 126796
rect 48458 126784 48464 126796
rect 38856 126756 48464 126784
rect 38856 126744 38862 126756
rect 48458 126744 48464 126756
rect 48516 126744 48522 126796
rect 357670 126744 357676 126796
rect 357728 126784 357734 126796
rect 405970 126784 405976 126796
rect 357728 126756 405976 126784
rect 357728 126744 357734 126756
rect 405970 126744 405976 126756
rect 406028 126744 406034 126796
rect 38246 126064 38252 126116
rect 38304 126104 38310 126116
rect 52598 126104 52604 126116
rect 38304 126076 52604 126104
rect 38304 126064 38310 126076
rect 52598 126064 52604 126076
rect 52656 126064 52662 126116
rect 356198 126064 356204 126116
rect 356256 126104 356262 126116
rect 405970 126104 405976 126116
rect 356256 126076 405976 126104
rect 356256 126064 356262 126076
rect 405970 126064 405976 126076
rect 406028 126064 406034 126116
rect 76886 125452 76892 125504
rect 76944 125492 76950 125504
rect 82682 125492 82688 125504
rect 76944 125464 82688 125492
rect 76944 125452 76950 125464
rect 82682 125452 82688 125464
rect 82740 125452 82746 125504
rect 169990 125384 169996 125436
rect 170048 125424 170054 125436
rect 170726 125424 170732 125436
rect 170048 125396 170732 125424
rect 170048 125384 170054 125396
rect 170726 125384 170732 125396
rect 170784 125424 170790 125436
rect 175510 125424 175516 125436
rect 170784 125396 175516 125424
rect 170784 125384 170790 125396
rect 175510 125384 175516 125396
rect 175568 125384 175574 125436
rect 263830 125248 263836 125300
rect 263888 125288 263894 125300
rect 264474 125288 264480 125300
rect 263888 125260 264480 125288
rect 263888 125248 263894 125260
rect 264474 125248 264480 125260
rect 264532 125288 264538 125300
rect 270362 125288 270368 125300
rect 264532 125260 270368 125288
rect 264532 125248 264538 125260
rect 270362 125248 270368 125260
rect 270420 125248 270426 125300
rect 76150 125044 76156 125096
rect 76208 125084 76214 125096
rect 76886 125084 76892 125096
rect 76208 125056 76892 125084
rect 76208 125044 76214 125056
rect 76886 125044 76892 125056
rect 76944 125044 76950 125096
rect 12670 123276 12676 123328
rect 12728 123316 12734 123328
rect 16166 123316 16172 123328
rect 12728 123288 16172 123316
rect 12728 123276 12734 123288
rect 16166 123276 16172 123288
rect 16224 123276 16230 123328
rect 38798 122596 38804 122648
rect 38856 122636 38862 122648
rect 54070 122636 54076 122648
rect 38856 122608 54076 122636
rect 38856 122596 38862 122608
rect 54070 122596 54076 122608
rect 54128 122596 54134 122648
rect 356290 122596 356296 122648
rect 356348 122636 356354 122648
rect 405970 122636 405976 122648
rect 356348 122608 405976 122636
rect 356348 122596 356354 122608
rect 405970 122596 405976 122608
rect 406028 122596 406034 122648
rect 137606 121984 137612 122036
rect 137664 122024 137670 122036
rect 144230 122024 144236 122036
rect 137664 121996 144236 122024
rect 137664 121984 137670 121996
rect 144230 121984 144236 121996
rect 144288 121984 144294 122036
rect 231446 121984 231452 122036
rect 231504 122024 231510 122036
rect 240370 122024 240376 122036
rect 231504 121996 240376 122024
rect 231504 121984 231510 121996
rect 240370 121984 240376 121996
rect 240428 121984 240434 122036
rect 325286 121984 325292 122036
rect 325344 122024 325350 122036
rect 334210 122024 334216 122036
rect 325344 121996 334216 122024
rect 325344 121984 325350 121996
rect 334210 121984 334216 121996
rect 334268 121984 334274 122036
rect 38798 120556 38804 120608
rect 38856 120596 38862 120608
rect 52598 120596 52604 120608
rect 38856 120568 52604 120596
rect 38856 120556 38862 120568
rect 52598 120556 52604 120568
rect 52656 120556 52662 120608
rect 356198 120556 356204 120608
rect 356256 120596 356262 120608
rect 405970 120596 405976 120608
rect 356256 120568 405976 120596
rect 356256 120556 356262 120568
rect 405970 120556 405976 120568
rect 406028 120556 406034 120608
rect 324550 119876 324556 119928
rect 324608 119916 324614 119928
rect 326574 119916 326580 119928
rect 324608 119888 326580 119916
rect 324608 119876 324614 119888
rect 326574 119876 326580 119888
rect 326632 119876 326638 119928
rect 262358 117904 262364 117956
rect 262416 117944 262422 117956
rect 269994 117944 270000 117956
rect 262416 117916 270000 117944
rect 262416 117904 262422 117916
rect 269994 117904 270000 117916
rect 270052 117904 270058 117956
rect 167874 117836 167880 117888
rect 167932 117876 167938 117888
rect 176246 117876 176252 117888
rect 167932 117848 176252 117876
rect 167932 117836 167938 117848
rect 176246 117836 176252 117848
rect 176304 117836 176310 117888
rect 38246 117088 38252 117140
rect 38304 117128 38310 117140
rect 54070 117128 54076 117140
rect 38304 117100 54076 117128
rect 38304 117088 38310 117100
rect 54070 117088 54076 117100
rect 54128 117088 54134 117140
rect 354910 117088 354916 117140
rect 354968 117128 354974 117140
rect 405970 117128 405976 117140
rect 354968 117100 405976 117128
rect 354968 117088 354974 117100
rect 405970 117088 405976 117100
rect 406028 117088 406034 117140
rect 427406 116408 427412 116460
rect 427464 116448 427470 116460
rect 429430 116448 429436 116460
rect 427464 116420 429436 116448
rect 427464 116408 427470 116420
rect 429430 116408 429436 116420
rect 429488 116408 429494 116460
rect 51589 115159 51647 115165
rect 51589 115125 51601 115159
rect 51635 115156 51647 115159
rect 51678 115156 51684 115168
rect 51635 115128 51684 115156
rect 51635 115125 51647 115128
rect 51589 115119 51647 115125
rect 51678 115116 51684 115128
rect 51736 115116 51742 115168
rect 38798 115048 38804 115100
rect 38856 115088 38862 115100
rect 52138 115088 52144 115100
rect 38856 115060 52144 115088
rect 38856 115048 38862 115060
rect 52138 115048 52144 115060
rect 52196 115048 52202 115100
rect 356198 115048 356204 115100
rect 356256 115088 356262 115100
rect 405970 115088 405976 115100
rect 356256 115060 405976 115088
rect 356256 115048 356262 115060
rect 405970 115048 405976 115060
rect 406028 115048 406034 115100
rect 51586 113728 51592 113740
rect 51547 113700 51592 113728
rect 51586 113688 51592 113700
rect 51644 113688 51650 113740
rect 38798 112940 38804 112992
rect 38856 112980 38862 112992
rect 51862 112980 51868 112992
rect 38856 112952 51868 112980
rect 38856 112940 38862 112952
rect 51862 112940 51868 112952
rect 51920 112940 51926 112992
rect 136870 112940 136876 112992
rect 136928 112980 136934 112992
rect 146622 112980 146628 112992
rect 136928 112952 146628 112980
rect 136928 112940 136934 112952
rect 146622 112940 146628 112952
rect 146680 112940 146686 112992
rect 355002 112940 355008 112992
rect 355060 112980 355066 112992
rect 405970 112980 405976 112992
rect 355060 112952 405976 112980
rect 355060 112940 355066 112952
rect 405970 112940 405976 112952
rect 406028 112940 406034 112992
rect 52598 111008 52604 111020
rect 48476 110980 52604 111008
rect 38246 110900 38252 110952
rect 38304 110940 38310 110952
rect 48476 110940 48504 110980
rect 52598 110968 52604 110980
rect 52656 110968 52662 111020
rect 427590 110968 427596 111020
rect 427648 111008 427654 111020
rect 428786 111008 428792 111020
rect 427648 110980 428792 111008
rect 427648 110968 427654 110980
rect 428786 110968 428792 110980
rect 428844 110968 428850 111020
rect 38304 110912 48504 110940
rect 38304 110900 38310 110912
rect 136870 110900 136876 110952
rect 136928 110940 136934 110952
rect 145334 110940 145340 110952
rect 136928 110912 145340 110940
rect 136928 110900 136934 110912
rect 145334 110900 145340 110912
rect 145392 110900 145398 110952
rect 356198 110900 356204 110952
rect 356256 110940 356262 110952
rect 406062 110940 406068 110952
rect 356256 110912 406068 110940
rect 356256 110900 356262 110912
rect 406062 110900 406068 110912
rect 406120 110900 406126 110952
rect 84706 109744 84712 109796
rect 84764 109784 84770 109796
rect 85810 109784 85816 109796
rect 84764 109756 85816 109784
rect 84764 109744 84770 109756
rect 85810 109744 85816 109756
rect 85868 109744 85874 109796
rect 231998 109540 232004 109592
rect 232056 109580 232062 109592
rect 238990 109580 238996 109592
rect 232056 109552 238996 109580
rect 232056 109540 232062 109552
rect 238990 109540 238996 109552
rect 239048 109580 239054 109592
rect 240094 109580 240100 109592
rect 239048 109552 240100 109580
rect 239048 109540 239054 109552
rect 240094 109540 240100 109552
rect 240152 109540 240158 109592
rect 74310 109472 74316 109524
rect 74368 109512 74374 109524
rect 82590 109512 82596 109524
rect 74368 109484 82596 109512
rect 74368 109472 74374 109484
rect 82590 109472 82596 109484
rect 82648 109472 82654 109524
rect 51586 108248 51592 108300
rect 51644 108288 51650 108300
rect 51681 108291 51739 108297
rect 51681 108288 51693 108291
rect 51644 108260 51693 108288
rect 51644 108248 51650 108260
rect 51681 108257 51693 108260
rect 51727 108257 51739 108291
rect 51681 108251 51739 108257
rect 137698 108180 137704 108232
rect 137756 108220 137762 108232
rect 143954 108220 143960 108232
rect 137756 108192 143960 108220
rect 137756 108180 137762 108192
rect 143954 108180 143960 108192
rect 144012 108180 144018 108232
rect 231538 108180 231544 108232
rect 231596 108220 231602 108232
rect 240830 108220 240836 108232
rect 231596 108192 240836 108220
rect 231596 108180 231602 108192
rect 240830 108180 240836 108192
rect 240888 108180 240894 108232
rect 325378 108180 325384 108232
rect 325436 108220 325442 108232
rect 334210 108220 334216 108232
rect 325436 108192 334216 108220
rect 325436 108180 325442 108192
rect 334210 108180 334216 108192
rect 334268 108180 334274 108232
rect 358314 108180 358320 108232
rect 358372 108180 358378 108232
rect 358332 108096 358360 108180
rect 358314 108044 358320 108096
rect 358372 108044 358378 108096
rect 38798 107432 38804 107484
rect 38856 107472 38862 107484
rect 51681 107475 51739 107481
rect 51681 107472 51693 107475
rect 38856 107444 51693 107472
rect 38856 107432 38862 107444
rect 51681 107441 51693 107444
rect 51727 107441 51739 107475
rect 51681 107435 51739 107441
rect 353530 107432 353536 107484
rect 353588 107472 353594 107484
rect 405970 107472 405976 107484
rect 353588 107444 405976 107472
rect 353588 107432 353594 107444
rect 405970 107432 405976 107444
rect 406028 107432 406034 107484
rect 13314 105460 13320 105512
rect 13372 105500 13378 105512
rect 18098 105500 18104 105512
rect 13372 105472 18104 105500
rect 13372 105460 13378 105472
rect 18098 105460 18104 105472
rect 18156 105460 18162 105512
rect 427590 105460 427596 105512
rect 427648 105500 427654 105512
rect 430074 105500 430080 105512
rect 427648 105472 430080 105500
rect 427648 105460 427654 105472
rect 430074 105460 430080 105472
rect 430132 105460 430138 105512
rect 38798 105392 38804 105444
rect 38856 105432 38862 105444
rect 52598 105432 52604 105444
rect 38856 105404 52604 105432
rect 38856 105392 38862 105404
rect 52598 105392 52604 105404
rect 52656 105392 52662 105444
rect 356198 105392 356204 105444
rect 356256 105432 356262 105444
rect 405970 105432 405976 105444
rect 356256 105404 405976 105432
rect 356256 105392 356262 105404
rect 405970 105392 405976 105404
rect 406028 105392 406034 105444
rect 358314 105364 358320 105376
rect 358275 105336 358320 105364
rect 358314 105324 358320 105336
rect 358372 105324 358378 105376
rect 51678 104072 51684 104084
rect 51639 104044 51684 104072
rect 51678 104032 51684 104044
rect 51736 104032 51742 104084
rect 427590 102672 427596 102724
rect 427648 102712 427654 102724
rect 429430 102712 429436 102724
rect 427648 102684 429436 102712
rect 427648 102672 427654 102684
rect 429430 102672 429436 102684
rect 429488 102672 429494 102724
rect 352702 101924 352708 101976
rect 352760 101964 352766 101976
rect 405970 101964 405976 101976
rect 352760 101936 405976 101964
rect 352760 101924 352766 101936
rect 405970 101924 405976 101936
rect 406028 101924 406034 101976
rect 50022 101516 50028 101568
rect 50080 101556 50086 101568
rect 51310 101556 51316 101568
rect 50080 101528 51316 101556
rect 50080 101516 50086 101528
rect 51310 101516 51316 101528
rect 51368 101516 51374 101568
rect 38614 101312 38620 101364
rect 38672 101352 38678 101364
rect 50022 101352 50028 101364
rect 38672 101324 50028 101352
rect 38672 101312 38678 101324
rect 50022 101312 50028 101324
rect 50080 101312 50086 101364
rect 38798 100564 38804 100616
rect 38856 100604 38862 100616
rect 52598 100604 52604 100616
rect 38856 100576 52604 100604
rect 38856 100564 38862 100576
rect 52598 100564 52604 100576
rect 52656 100564 52662 100616
rect 356198 100564 356204 100616
rect 356256 100604 356262 100616
rect 405970 100604 405976 100616
rect 356256 100576 405976 100604
rect 356256 100564 356262 100576
rect 405970 100564 405976 100576
rect 406028 100564 406034 100616
rect 13498 99884 13504 99936
rect 13556 99924 13562 99936
rect 17454 99924 17460 99936
rect 13556 99896 17460 99924
rect 13556 99884 13562 99896
rect 17454 99884 17460 99896
rect 17512 99884 17518 99936
rect 167874 98524 167880 98576
rect 167932 98564 167938 98576
rect 173394 98564 173400 98576
rect 167932 98536 173400 98564
rect 167932 98524 167938 98536
rect 173394 98524 173400 98536
rect 173452 98524 173458 98576
rect 261162 98524 261168 98576
rect 261220 98564 261226 98576
rect 267234 98564 267240 98576
rect 261220 98536 267240 98564
rect 261220 98524 261226 98536
rect 267234 98524 267240 98536
rect 267292 98524 267298 98576
rect 38798 97776 38804 97828
rect 38856 97816 38862 97828
rect 49930 97816 49936 97828
rect 38856 97788 49936 97816
rect 38856 97776 38862 97788
rect 49930 97776 49936 97788
rect 49988 97776 49994 97828
rect 352794 97776 352800 97828
rect 352852 97816 352858 97828
rect 405970 97816 405976 97828
rect 352852 97788 405976 97816
rect 352852 97776 352858 97788
rect 405970 97776 405976 97788
rect 406028 97776 406034 97828
rect 13130 95804 13136 95856
rect 13188 95844 13194 95856
rect 18098 95844 18104 95856
rect 13188 95816 18104 95844
rect 13188 95804 13194 95816
rect 18098 95804 18104 95816
rect 18156 95804 18162 95856
rect 52598 95844 52604 95856
rect 48476 95816 52604 95844
rect 38062 95736 38068 95788
rect 38120 95776 38126 95788
rect 48476 95776 48504 95816
rect 52598 95804 52604 95816
rect 52656 95804 52662 95856
rect 358314 95844 358320 95856
rect 358275 95816 358320 95844
rect 358314 95804 358320 95816
rect 358372 95804 358378 95856
rect 427222 95804 427228 95856
rect 427280 95844 427286 95856
rect 430166 95844 430172 95856
rect 427280 95816 430172 95844
rect 427280 95804 427286 95816
rect 430166 95804 430172 95816
rect 430224 95804 430230 95856
rect 38120 95748 48504 95776
rect 38120 95736 38126 95748
rect 356198 95736 356204 95788
rect 356256 95776 356262 95788
rect 405970 95776 405976 95788
rect 356256 95748 405976 95776
rect 356256 95736 356262 95748
rect 405970 95736 405976 95748
rect 406028 95736 406034 95788
rect 324550 95056 324556 95108
rect 324608 95096 324614 95108
rect 330070 95096 330076 95108
rect 324608 95068 330076 95096
rect 324608 95056 324614 95068
rect 330070 95056 330076 95068
rect 330128 95056 330134 95108
rect 231998 94988 232004 95040
rect 232056 95028 232062 95040
rect 236230 95028 236236 95040
rect 232056 95000 236236 95028
rect 232056 94988 232062 95000
rect 236230 94988 236236 95000
rect 236288 94988 236294 95040
rect 138158 94376 138164 94428
rect 138216 94416 138222 94428
rect 142390 94416 142396 94428
rect 138216 94388 142396 94416
rect 138216 94376 138222 94388
rect 142390 94376 142396 94388
rect 142448 94376 142454 94428
rect 235494 94376 235500 94428
rect 235552 94416 235558 94428
rect 240370 94416 240376 94428
rect 235552 94388 240376 94416
rect 235552 94376 235558 94388
rect 240370 94376 240376 94388
rect 240428 94376 240434 94428
rect 329334 94376 329340 94428
rect 329392 94416 329398 94428
rect 334210 94416 334216 94428
rect 329392 94388 334216 94416
rect 329392 94376 329398 94388
rect 334210 94376 334216 94388
rect 334268 94376 334274 94428
rect 73390 93696 73396 93748
rect 73448 93736 73454 93748
rect 73666 93736 73672 93748
rect 73448 93708 73672 93736
rect 73448 93696 73454 93708
rect 73666 93696 73672 93708
rect 73724 93696 73730 93748
rect 84798 93424 84804 93476
rect 84856 93464 84862 93476
rect 85810 93464 85816 93476
rect 84856 93436 85816 93464
rect 84856 93424 84862 93436
rect 85810 93424 85816 93436
rect 85868 93424 85874 93476
rect 267234 92948 267240 93000
rect 267292 92988 267298 93000
rect 270362 92988 270368 93000
rect 267292 92960 270368 92988
rect 267292 92948 267298 92960
rect 270362 92948 270368 92960
rect 270420 92948 270426 93000
rect 75414 92676 75420 92728
rect 75472 92716 75478 92728
rect 82682 92716 82688 92728
rect 75472 92688 82688 92716
rect 75472 92676 75478 92688
rect 82682 92676 82688 92688
rect 82740 92676 82746 92728
rect 173394 92540 173400 92592
rect 173452 92580 173458 92592
rect 175510 92580 175516 92592
rect 173452 92552 175516 92580
rect 173452 92540 173458 92552
rect 175510 92540 175516 92552
rect 175568 92540 175574 92592
rect 37602 92268 37608 92320
rect 37660 92308 37666 92320
rect 48550 92308 48556 92320
rect 37660 92280 48556 92308
rect 37660 92268 37666 92280
rect 48550 92268 48556 92280
rect 48608 92268 48614 92320
rect 352794 92268 352800 92320
rect 352852 92308 352858 92320
rect 405970 92308 405976 92320
rect 352852 92280 405976 92308
rect 352852 92268 352858 92280
rect 405970 92268 405976 92280
rect 406028 92268 406034 92320
rect 13406 91588 13412 91640
rect 13464 91628 13470 91640
rect 18098 91628 18104 91640
rect 13464 91600 18104 91628
rect 13464 91588 13470 91600
rect 18098 91588 18104 91600
rect 18156 91588 18162 91640
rect 73390 91452 73396 91504
rect 73448 91492 73454 91504
rect 76794 91492 76800 91504
rect 73448 91464 76800 91492
rect 73448 91452 73454 91464
rect 76794 91452 76800 91464
rect 76852 91452 76858 91504
rect 38798 90160 38804 90212
rect 38856 90200 38862 90212
rect 52598 90200 52604 90212
rect 38856 90172 52604 90200
rect 38856 90160 38862 90172
rect 52598 90160 52604 90172
rect 52656 90160 52662 90212
rect 356198 90160 356204 90212
rect 356256 90200 356262 90212
rect 405970 90200 405976 90212
rect 356256 90172 405976 90200
rect 356256 90160 356262 90172
rect 405970 90160 405976 90172
rect 406028 90160 406034 90212
rect 51497 89047 51555 89053
rect 51497 89013 51509 89047
rect 51543 89044 51555 89047
rect 51678 89044 51684 89056
rect 51543 89016 51684 89044
rect 51543 89013 51555 89016
rect 51497 89007 51555 89013
rect 51678 89004 51684 89016
rect 51736 89004 51742 89056
rect 358314 88868 358320 88920
rect 358372 88908 358378 88920
rect 358372 88880 358452 88908
rect 358372 88868 358378 88880
rect 358424 88716 358452 88880
rect 358406 88664 358412 88716
rect 358464 88664 358470 88716
rect 35949 87551 36007 87557
rect 35949 87517 35961 87551
rect 35995 87548 36007 87551
rect 45701 87551 45759 87557
rect 35995 87520 36176 87548
rect 35995 87517 36007 87520
rect 35949 87511 36007 87517
rect 23894 87440 23900 87492
rect 23952 87480 23958 87492
rect 36148 87489 36176 87520
rect 45701 87517 45713 87551
rect 45747 87548 45759 87551
rect 45747 87520 45928 87548
rect 45747 87517 45759 87520
rect 45701 87511 45759 87517
rect 45900 87489 45928 87520
rect 26473 87483 26531 87489
rect 26473 87480 26485 87483
rect 23952 87452 26485 87480
rect 23952 87440 23958 87452
rect 26473 87449 26485 87452
rect 26519 87449 26531 87483
rect 26473 87443 26531 87449
rect 36133 87483 36191 87489
rect 36133 87449 36145 87483
rect 36179 87449 36191 87483
rect 36133 87443 36191 87449
rect 45885 87483 45943 87489
rect 45885 87449 45897 87483
rect 45931 87449 45943 87483
rect 45885 87443 45943 87449
rect 65021 87483 65079 87489
rect 65021 87449 65033 87483
rect 65067 87480 65079 87483
rect 72010 87480 72016 87492
rect 65067 87452 72016 87480
rect 65067 87449 65079 87452
rect 65021 87443 65079 87449
rect 72010 87440 72016 87452
rect 72068 87440 72074 87492
rect 150394 87440 150400 87492
rect 150452 87480 150458 87492
rect 154074 87480 154080 87492
rect 150452 87452 154080 87480
rect 150452 87440 150458 87452
rect 154074 87440 154080 87452
rect 154132 87440 154138 87492
rect 154718 87440 154724 87492
rect 154776 87480 154782 87492
rect 172014 87480 172020 87492
rect 154776 87452 172020 87480
rect 154776 87440 154782 87452
rect 172014 87440 172020 87452
rect 172072 87440 172078 87492
rect 361074 87440 361080 87492
rect 361132 87480 361138 87492
rect 418206 87480 418212 87492
rect 361132 87452 418212 87480
rect 361132 87440 361138 87452
rect 418206 87440 418212 87452
rect 418264 87440 418270 87492
rect 36038 87372 36044 87424
rect 36096 87412 36102 87424
rect 45793 87415 45851 87421
rect 45793 87412 45805 87415
rect 36096 87384 45805 87412
rect 36096 87372 36102 87384
rect 45793 87381 45805 87384
rect 45839 87381 45851 87415
rect 45793 87375 45851 87381
rect 56097 87415 56155 87421
rect 56097 87381 56109 87415
rect 56143 87412 56155 87415
rect 73850 87412 73856 87424
rect 56143 87384 73856 87412
rect 56143 87381 56155 87384
rect 56097 87375 56155 87381
rect 73850 87372 73856 87384
rect 73908 87372 73914 87424
rect 160974 87372 160980 87424
rect 161032 87412 161038 87424
rect 163918 87412 163924 87424
rect 161032 87384 163924 87412
rect 161032 87372 161038 87384
rect 163918 87372 163924 87384
rect 163976 87372 163982 87424
rect 249018 87372 249024 87424
rect 249076 87412 249082 87424
rect 258954 87412 258960 87424
rect 249076 87384 258960 87412
rect 249076 87372 249082 87384
rect 258954 87372 258960 87384
rect 259012 87372 259018 87424
rect 359694 87372 359700 87424
rect 359752 87412 359758 87424
rect 360338 87412 360344 87424
rect 359752 87384 360344 87412
rect 359752 87372 359758 87384
rect 360338 87372 360344 87384
rect 360396 87412 360402 87424
rect 415538 87412 415544 87424
rect 360396 87384 415544 87412
rect 360396 87372 360402 87384
rect 415538 87372 415544 87384
rect 415596 87372 415602 87424
rect 29230 87304 29236 87356
rect 29288 87344 29294 87356
rect 73574 87344 73580 87356
rect 29288 87316 73580 87344
rect 29288 87304 29294 87316
rect 73574 87304 73580 87316
rect 73632 87304 73638 87356
rect 149750 87304 149756 87356
rect 149808 87344 149814 87356
rect 154166 87344 154172 87356
rect 149808 87316 154172 87344
rect 149808 87304 149814 87316
rect 154166 87304 154172 87316
rect 154224 87304 154230 87356
rect 343502 87304 343508 87356
rect 343560 87344 343566 87356
rect 348194 87344 348200 87356
rect 343560 87316 348200 87344
rect 343560 87304 343566 87316
rect 348194 87304 348200 87316
rect 348252 87304 348258 87356
rect 369998 87304 370004 87356
rect 370056 87344 370062 87356
rect 410202 87344 410208 87356
rect 370056 87316 410208 87344
rect 370056 87304 370062 87316
rect 410202 87304 410208 87316
rect 410260 87304 410266 87356
rect 31898 87236 31904 87288
rect 31956 87276 31962 87288
rect 73482 87276 73488 87288
rect 31956 87248 73488 87276
rect 31956 87236 31962 87248
rect 73482 87236 73488 87248
rect 73540 87236 73546 87288
rect 151038 87236 151044 87288
rect 151096 87276 151102 87288
rect 155454 87276 155460 87288
rect 151096 87248 155460 87276
rect 151096 87236 151102 87248
rect 155454 87236 155460 87248
rect 155512 87236 155518 87288
rect 244418 87236 244424 87288
rect 244476 87276 244482 87288
rect 254170 87276 254176 87288
rect 244476 87248 254176 87276
rect 244476 87236 244482 87248
rect 254170 87236 254176 87248
rect 254228 87236 254234 87288
rect 340926 87236 340932 87288
rect 340984 87276 340990 87288
rect 345250 87276 345256 87288
rect 340984 87248 345256 87276
rect 340984 87236 340990 87248
rect 345250 87236 345256 87248
rect 345308 87236 345314 87288
rect 34566 87168 34572 87220
rect 34624 87208 34630 87220
rect 73666 87208 73672 87220
rect 34624 87180 73672 87208
rect 34624 87168 34630 87180
rect 73666 87168 73672 87180
rect 73724 87168 73730 87220
rect 336878 87168 336884 87220
rect 336936 87208 336942 87220
rect 348746 87208 348752 87220
rect 336936 87180 348752 87208
rect 336936 87168 336942 87180
rect 348746 87168 348752 87180
rect 348804 87168 348810 87220
rect 21226 87100 21232 87152
rect 21284 87140 21290 87152
rect 34658 87140 34664 87152
rect 21284 87112 34664 87140
rect 21284 87100 21290 87112
rect 34658 87100 34664 87112
rect 34716 87100 34722 87152
rect 36133 87143 36191 87149
rect 36133 87109 36145 87143
rect 36179 87140 36191 87143
rect 45701 87143 45759 87149
rect 45701 87140 45713 87143
rect 36179 87112 45713 87140
rect 36179 87109 36191 87112
rect 36133 87103 36191 87109
rect 45701 87109 45713 87112
rect 45747 87109 45759 87143
rect 45701 87103 45759 87109
rect 45793 87143 45851 87149
rect 45793 87109 45805 87143
rect 45839 87140 45851 87143
rect 56097 87143 56155 87149
rect 56097 87140 56109 87143
rect 45839 87112 56109 87140
rect 45839 87109 45851 87112
rect 45793 87103 45851 87109
rect 56097 87109 56109 87112
rect 56143 87109 56155 87143
rect 56097 87103 56155 87109
rect 64374 87100 64380 87152
rect 64432 87140 64438 87152
rect 65938 87140 65944 87152
rect 64432 87112 65944 87140
rect 64432 87100 64438 87112
rect 65938 87100 65944 87112
rect 65996 87100 66002 87152
rect 149198 87100 149204 87152
rect 149256 87140 149262 87152
rect 157570 87140 157576 87152
rect 149256 87112 157576 87140
rect 149256 87100 149262 87112
rect 157570 87100 157576 87112
rect 157628 87100 157634 87152
rect 243038 87100 243044 87152
rect 243096 87140 243102 87152
rect 255090 87140 255096 87152
rect 243096 87112 255096 87140
rect 243096 87100 243102 87112
rect 255090 87100 255096 87112
rect 255148 87100 255154 87152
rect 338074 87100 338080 87152
rect 338132 87140 338138 87152
rect 349574 87140 349580 87152
rect 338132 87112 349580 87140
rect 338132 87100 338138 87112
rect 349574 87100 349580 87112
rect 349632 87100 349638 87152
rect 26562 87032 26568 87084
rect 26620 87072 26626 87084
rect 36038 87072 36044 87084
rect 26620 87044 36044 87072
rect 26620 87032 26626 87044
rect 36038 87032 36044 87044
rect 36096 87032 36102 87084
rect 45885 87075 45943 87081
rect 45885 87041 45897 87075
rect 45931 87072 45943 87075
rect 65021 87075 65079 87081
rect 65021 87072 65033 87075
rect 45931 87044 65033 87072
rect 45931 87041 45943 87044
rect 45885 87035 45943 87041
rect 65021 87041 65033 87044
rect 65067 87041 65079 87075
rect 65021 87035 65079 87041
rect 150578 87032 150584 87084
rect 150636 87072 150642 87084
rect 162078 87072 162084 87084
rect 150636 87044 162084 87072
rect 150636 87032 150642 87044
rect 162078 87032 162084 87044
rect 162136 87032 162142 87084
rect 339638 87032 339644 87084
rect 339696 87072 339702 87084
rect 351230 87072 351236 87084
rect 339696 87044 351236 87072
rect 339696 87032 339702 87044
rect 351230 87032 351236 87044
rect 351288 87032 351294 87084
rect 26473 87007 26531 87013
rect 26473 86973 26485 87007
rect 26519 87004 26531 87007
rect 35949 87007 36007 87013
rect 35949 87004 35961 87007
rect 26519 86976 35961 87004
rect 26519 86973 26531 86976
rect 26473 86967 26531 86973
rect 35949 86973 35961 86976
rect 35995 86973 36007 87007
rect 35949 86967 36007 86973
rect 59682 86964 59688 87016
rect 59740 87004 59746 87016
rect 67134 87004 67140 87016
rect 59740 86976 67140 87004
rect 59740 86964 59746 86976
rect 67134 86964 67140 86976
rect 67192 86964 67198 87016
rect 149198 86964 149204 87016
rect 149256 87004 149262 87016
rect 161434 87004 161440 87016
rect 149256 86976 161440 87004
rect 149256 86964 149262 86976
rect 161434 86964 161440 86976
rect 161492 86964 161498 87016
rect 241658 86964 241664 87016
rect 241716 87004 241722 87016
rect 254538 87004 254544 87016
rect 241716 86976 254544 87004
rect 241716 86964 241722 86976
rect 254538 86964 254544 86976
rect 254596 86964 254602 87016
rect 334118 86964 334124 87016
rect 334176 87004 334182 87016
rect 334176 86976 340420 87004
rect 334176 86964 334182 86976
rect 146438 86896 146444 86948
rect 146496 86936 146502 86948
rect 160238 86936 160244 86948
rect 146496 86908 160244 86936
rect 146496 86896 146502 86908
rect 160238 86896 160244 86908
rect 160296 86896 160302 86948
rect 244050 86896 244056 86948
rect 244108 86936 244114 86948
rect 252974 86936 252980 86948
rect 244108 86908 252980 86936
rect 244108 86896 244114 86908
rect 252974 86896 252980 86908
rect 253032 86896 253038 86948
rect 335406 86896 335412 86948
rect 335464 86936 335470 86948
rect 339917 86939 339975 86945
rect 339917 86936 339929 86939
rect 335464 86908 339929 86936
rect 335464 86896 335470 86908
rect 339917 86905 339929 86908
rect 339963 86905 339975 86939
rect 340392 86936 340420 86976
rect 341018 86964 341024 87016
rect 341076 87004 341082 87016
rect 352150 87004 352156 87016
rect 341076 86976 352156 87004
rect 341076 86964 341082 86976
rect 352150 86964 352156 86976
rect 352208 86964 352214 87016
rect 346170 86936 346176 86948
rect 340392 86908 346176 86936
rect 339917 86899 339975 86905
rect 346170 86896 346176 86908
rect 346228 86896 346234 86948
rect 57014 86828 57020 86880
rect 57072 86868 57078 86880
rect 67870 86868 67876 86880
rect 57072 86840 67876 86868
rect 57072 86828 57078 86840
rect 67870 86828 67876 86840
rect 67928 86828 67934 86880
rect 147818 86828 147824 86880
rect 147876 86868 147882 86880
rect 160882 86868 160888 86880
rect 147876 86840 160888 86868
rect 147876 86828 147882 86840
rect 160882 86828 160888 86840
rect 160940 86828 160946 86880
rect 240278 86828 240284 86880
rect 240336 86868 240342 86880
rect 254262 86868 254268 86880
rect 240336 86840 254268 86868
rect 240336 86828 240342 86840
rect 254262 86828 254268 86840
rect 254320 86828 254326 86880
rect 335498 86828 335504 86880
rect 335556 86868 335562 86880
rect 348010 86868 348016 86880
rect 335556 86840 348016 86868
rect 335556 86828 335562 86840
rect 348010 86828 348016 86840
rect 348068 86828 348074 86880
rect 56094 86760 56100 86812
rect 56152 86800 56158 86812
rect 66674 86800 66680 86812
rect 56152 86772 66680 86800
rect 56152 86760 56158 86772
rect 66674 86760 66680 86772
rect 66732 86760 66738 86812
rect 145058 86760 145064 86812
rect 145116 86800 145122 86812
rect 159594 86800 159600 86812
rect 145116 86772 159600 86800
rect 145116 86760 145122 86772
rect 159594 86760 159600 86772
rect 159652 86760 159658 86812
rect 238898 86760 238904 86812
rect 238956 86800 238962 86812
rect 253434 86800 253440 86812
rect 238956 86772 253440 86800
rect 238956 86760 238962 86772
rect 253434 86760 253440 86772
rect 253492 86760 253498 86812
rect 332738 86760 332744 86812
rect 332796 86800 332802 86812
rect 345342 86800 345348 86812
rect 332796 86772 345348 86800
rect 332796 86760 332802 86772
rect 345342 86760 345348 86772
rect 345400 86760 345406 86812
rect 339917 86735 339975 86741
rect 339917 86701 339929 86735
rect 339963 86732 339975 86735
rect 346998 86732 347004 86744
rect 339963 86704 347004 86732
rect 339963 86701 339975 86704
rect 339917 86695 339975 86701
rect 346998 86692 347004 86704
rect 347056 86692 347062 86744
rect 344330 86624 344336 86676
rect 344388 86664 344394 86676
rect 347274 86664 347280 86676
rect 344388 86636 347280 86664
rect 344388 86624 344394 86636
rect 347274 86624 347280 86636
rect 347332 86624 347338 86676
rect 257574 86488 257580 86540
rect 257632 86528 257638 86540
rect 258402 86528 258408 86540
rect 257632 86500 258408 86528
rect 257632 86488 257638 86500
rect 258402 86488 258408 86500
rect 258460 86488 258466 86540
rect 345066 86488 345072 86540
rect 345124 86528 345130 86540
rect 362454 86528 362460 86540
rect 345124 86500 362460 86528
rect 345124 86488 345130 86500
rect 362454 86488 362460 86500
rect 362512 86488 362518 86540
rect 252146 86216 252152 86268
rect 252204 86256 252210 86268
rect 255734 86256 255740 86268
rect 252204 86228 255740 86256
rect 252204 86216 252210 86228
rect 255734 86216 255740 86228
rect 255792 86216 255798 86268
rect 61614 86148 61620 86200
rect 61672 86188 61678 86200
rect 63270 86188 63276 86200
rect 61672 86160 63276 86188
rect 61672 86148 61678 86160
rect 63270 86148 63276 86160
rect 63328 86148 63334 86200
rect 67226 86148 67232 86200
rect 67284 86188 67290 86200
rect 68606 86188 68612 86200
rect 67284 86160 68612 86188
rect 67284 86148 67290 86160
rect 68606 86148 68612 86160
rect 68664 86148 68670 86200
rect 162354 86148 162360 86200
rect 162412 86188 162418 86200
rect 164562 86188 164568 86200
rect 162412 86160 164568 86188
rect 162412 86148 162418 86160
rect 164562 86148 164568 86160
rect 164620 86148 164626 86200
rect 245338 86148 245344 86200
rect 245396 86188 245402 86200
rect 252054 86188 252060 86200
rect 245396 86160 252060 86188
rect 245396 86148 245402 86160
rect 252054 86148 252060 86160
rect 252112 86148 252118 86200
rect 257666 86188 257672 86200
rect 256212 86160 257672 86188
rect 51494 86120 51500 86132
rect 51455 86092 51500 86120
rect 51494 86080 51500 86092
rect 51552 86080 51558 86132
rect 61430 86080 61436 86132
rect 61488 86120 61494 86132
rect 62258 86120 62264 86132
rect 61488 86092 62264 86120
rect 61488 86080 61494 86092
rect 62258 86080 62264 86092
rect 62316 86080 62322 86132
rect 62350 86080 62356 86132
rect 62408 86120 62414 86132
rect 63638 86120 63644 86132
rect 62408 86092 63644 86120
rect 62408 86080 62414 86092
rect 63638 86080 63644 86092
rect 63696 86080 63702 86132
rect 63730 86080 63736 86132
rect 63788 86120 63794 86132
rect 64742 86120 64748 86132
rect 63788 86092 64748 86120
rect 63788 86080 63794 86092
rect 64742 86080 64748 86092
rect 64800 86080 64806 86132
rect 65754 86080 65760 86132
rect 65812 86120 65818 86132
rect 66766 86120 66772 86132
rect 65812 86092 66772 86120
rect 65812 86080 65818 86092
rect 66766 86080 66772 86092
rect 66824 86080 66830 86132
rect 68514 86080 68520 86132
rect 68572 86120 68578 86132
rect 69434 86120 69440 86132
rect 68572 86092 69440 86120
rect 68572 86080 68578 86092
rect 69434 86080 69440 86092
rect 69492 86080 69498 86132
rect 152234 86080 152240 86132
rect 152292 86120 152298 86132
rect 153246 86120 153252 86132
rect 152292 86092 153252 86120
rect 152292 86080 152298 86092
rect 153246 86080 153252 86092
rect 153304 86080 153310 86132
rect 153430 86080 153436 86132
rect 153488 86120 153494 86132
rect 154718 86120 154724 86132
rect 153488 86092 154724 86120
rect 153488 86080 153494 86092
rect 154718 86080 154724 86092
rect 154776 86080 154782 86132
rect 162446 86080 162452 86132
rect 162504 86120 162510 86132
rect 163274 86120 163280 86132
rect 162504 86092 163280 86120
rect 162504 86080 162510 86092
rect 163274 86080 163280 86092
rect 163332 86080 163338 86132
rect 243498 86080 243504 86132
rect 243556 86120 243562 86132
rect 245154 86120 245160 86132
rect 243556 86092 245160 86120
rect 243556 86080 243562 86092
rect 245154 86080 245160 86092
rect 245212 86080 245218 86132
rect 246534 86080 246540 86132
rect 246592 86120 246598 86132
rect 247086 86120 247092 86132
rect 246592 86092 247092 86120
rect 246592 86080 246598 86092
rect 247086 86080 247092 86092
rect 247144 86080 247150 86132
rect 247730 86080 247736 86132
rect 247788 86120 247794 86132
rect 248558 86120 248564 86132
rect 247788 86092 248564 86120
rect 247788 86080 247794 86092
rect 248558 86080 248564 86092
rect 248616 86080 248622 86132
rect 256212 86064 256240 86160
rect 257666 86148 257672 86160
rect 257724 86148 257730 86200
rect 337614 86148 337620 86200
rect 337672 86188 337678 86200
rect 339086 86188 339092 86200
rect 337672 86160 339092 86188
rect 337672 86148 337678 86160
rect 339086 86148 339092 86160
rect 339144 86148 339150 86200
rect 341662 86148 341668 86200
rect 341720 86188 341726 86200
rect 344606 86188 344612 86200
rect 341720 86160 344612 86188
rect 341720 86148 341726 86160
rect 344606 86148 344612 86160
rect 344664 86148 344670 86200
rect 256286 86080 256292 86132
rect 256344 86120 256350 86132
rect 256930 86120 256936 86132
rect 256344 86092 256936 86120
rect 256344 86080 256350 86092
rect 256930 86080 256936 86092
rect 256988 86080 256994 86132
rect 338258 86080 338264 86132
rect 338316 86120 338322 86132
rect 338994 86120 339000 86132
rect 338316 86092 339000 86120
rect 338316 86080 338322 86092
rect 338994 86080 339000 86092
rect 339052 86080 339058 86132
rect 340098 86080 340104 86132
rect 340156 86120 340162 86132
rect 341754 86120 341760 86132
rect 340156 86092 341760 86120
rect 340156 86080 340162 86092
rect 341754 86080 341760 86092
rect 341812 86080 341818 86132
rect 342398 86080 342404 86132
rect 342456 86120 342462 86132
rect 344514 86120 344520 86132
rect 342456 86092 344520 86120
rect 342456 86080 342462 86092
rect 344514 86080 344520 86092
rect 344572 86080 344578 86132
rect 345894 86080 345900 86132
rect 345952 86120 345958 86132
rect 350402 86120 350408 86132
rect 345952 86092 350408 86120
rect 345952 86080 345958 86092
rect 350402 86080 350408 86092
rect 350460 86080 350466 86132
rect 66582 86012 66588 86064
rect 66640 86052 66646 86064
rect 67318 86052 67324 86064
rect 66640 86024 67324 86052
rect 66640 86012 66646 86024
rect 67318 86012 67324 86024
rect 67376 86012 67382 86064
rect 137882 86012 137888 86064
rect 137940 86052 137946 86064
rect 145794 86052 145800 86064
rect 137940 86024 145800 86052
rect 137940 86012 137946 86024
rect 145794 86012 145800 86024
rect 145852 86012 145858 86064
rect 256194 86012 256200 86064
rect 256252 86012 256258 86064
rect 324550 86012 324556 86064
rect 324608 86052 324614 86064
rect 329334 86052 329340 86064
rect 324608 86024 329340 86052
rect 324608 86012 324614 86024
rect 329334 86012 329340 86024
rect 329392 86012 329398 86064
rect 358406 86052 358412 86064
rect 358367 86024 358412 86052
rect 358406 86012 358412 86024
rect 358464 86012 358470 86064
rect 231078 85740 231084 85792
rect 231136 85780 231142 85792
rect 235494 85780 235500 85792
rect 231136 85752 235500 85780
rect 231136 85740 231142 85752
rect 235494 85740 235500 85752
rect 235552 85740 235558 85792
rect 354910 84040 354916 84092
rect 354968 84080 354974 84092
rect 355830 84080 355836 84092
rect 354968 84052 355836 84080
rect 354968 84040 354974 84052
rect 355830 84040 355836 84052
rect 355888 84040 355894 84092
rect 88478 81932 88484 81984
rect 88536 81972 88542 81984
rect 178730 81972 178736 81984
rect 88536 81944 178736 81972
rect 88536 81932 88542 81944
rect 178730 81932 178736 81944
rect 178788 81932 178794 81984
rect 182410 81932 182416 81984
rect 182468 81972 182474 81984
rect 276342 81972 276348 81984
rect 182468 81944 276348 81972
rect 182468 81932 182474 81944
rect 276342 81932 276348 81944
rect 276400 81932 276406 81984
rect 95746 81864 95752 81916
rect 95804 81904 95810 81916
rect 170634 81904 170640 81916
rect 95804 81876 170640 81904
rect 95804 81864 95810 81876
rect 170634 81864 170640 81876
rect 170692 81904 170698 81916
rect 189494 81904 189500 81916
rect 170692 81876 189500 81904
rect 170692 81864 170698 81876
rect 189494 81864 189500 81876
rect 189552 81904 189558 81916
rect 283150 81904 283156 81916
rect 189552 81876 283156 81904
rect 189552 81864 189558 81876
rect 283150 81864 283156 81876
rect 283208 81864 283214 81916
rect 102922 81796 102928 81848
rect 102980 81836 102986 81848
rect 176154 81836 176160 81848
rect 102980 81808 176160 81836
rect 102980 81796 102986 81808
rect 176154 81796 176160 81808
rect 176212 81836 176218 81848
rect 196670 81836 196676 81848
rect 176212 81808 196676 81836
rect 176212 81796 176218 81808
rect 196670 81796 196676 81808
rect 196728 81836 196734 81848
rect 290326 81836 290332 81848
rect 196728 81808 290332 81836
rect 196728 81796 196734 81808
rect 290326 81796 290332 81808
rect 290384 81796 290390 81848
rect 285818 81320 285824 81372
rect 285876 81360 285882 81372
rect 297502 81360 297508 81372
rect 285876 81332 297508 81360
rect 285876 81320 285882 81332
rect 297502 81320 297508 81332
rect 297560 81320 297566 81372
rect 96758 81252 96764 81304
rect 96816 81292 96822 81304
rect 109822 81292 109828 81304
rect 96816 81264 109828 81292
rect 96816 81252 96822 81264
rect 109822 81252 109828 81264
rect 109880 81252 109886 81304
rect 190598 81252 190604 81304
rect 190656 81292 190662 81304
rect 203754 81292 203760 81304
rect 190656 81264 203760 81292
rect 190656 81252 190662 81264
rect 203754 81252 203760 81264
rect 203812 81252 203818 81304
rect 276342 81252 276348 81304
rect 276400 81292 276406 81304
rect 428050 81292 428056 81304
rect 276400 81264 428056 81292
rect 276400 81252 276406 81264
rect 428050 81252 428056 81264
rect 428108 81252 428114 81304
rect 224454 80572 224460 80624
rect 224512 80612 224518 80624
rect 225190 80612 225196 80624
rect 224512 80584 225196 80612
rect 224512 80572 224518 80584
rect 225190 80572 225196 80584
rect 225248 80572 225254 80624
rect 318294 80572 318300 80624
rect 318352 80612 318358 80624
rect 319122 80612 319128 80624
rect 318352 80584 319128 80612
rect 318352 80572 318358 80584
rect 319122 80572 319128 80584
rect 319180 80572 319186 80624
rect 236230 79348 236236 79400
rect 236288 79388 236294 79400
rect 237242 79388 237248 79400
rect 236288 79360 237248 79388
rect 236288 79348 236294 79360
rect 237242 79348 237248 79360
rect 237300 79348 237306 79400
rect 60234 79144 60240 79196
rect 60292 79184 60298 79196
rect 64374 79184 64380 79196
rect 60292 79156 64380 79184
rect 60292 79144 60298 79156
rect 64374 79144 64380 79156
rect 64432 79144 64438 79196
rect 64469 79187 64527 79193
rect 64469 79153 64481 79187
rect 64515 79184 64527 79187
rect 66582 79184 66588 79196
rect 64515 79156 66588 79184
rect 64515 79153 64527 79156
rect 64469 79147 64527 79153
rect 66582 79144 66588 79156
rect 66640 79144 66646 79196
rect 75782 79144 75788 79196
rect 75840 79184 75846 79196
rect 76886 79184 76892 79196
rect 75840 79156 76892 79184
rect 75840 79144 75846 79156
rect 76886 79144 76892 79156
rect 76944 79144 76950 79196
rect 155454 79144 155460 79196
rect 155512 79184 155518 79196
rect 161710 79184 161716 79196
rect 155512 79156 161716 79184
rect 155512 79144 155518 79156
rect 161710 79144 161716 79156
rect 161768 79144 161774 79196
rect 245154 79144 245160 79196
rect 245212 79184 245218 79196
rect 251410 79184 251416 79196
rect 245212 79156 251416 79184
rect 245212 79144 245218 79156
rect 251410 79144 251416 79156
rect 251468 79144 251474 79196
rect 252054 79144 252060 79196
rect 252112 79184 252118 79196
rect 255550 79184 255556 79196
rect 252112 79156 255556 79184
rect 252112 79144 252118 79156
rect 255550 79144 255556 79156
rect 255608 79144 255614 79196
rect 333382 79144 333388 79196
rect 333440 79184 333446 79196
rect 334118 79184 334124 79196
rect 333440 79156 334124 79184
rect 333440 79144 333446 79156
rect 334118 79144 334124 79156
rect 334176 79144 334182 79196
rect 334394 79144 334400 79196
rect 334452 79184 334458 79196
rect 335406 79184 335412 79196
rect 334452 79156 335412 79184
rect 334452 79144 334458 79156
rect 335406 79144 335412 79156
rect 335464 79144 335470 79196
rect 339546 79144 339552 79196
rect 339604 79184 339610 79196
rect 343778 79184 343784 79196
rect 339604 79156 343784 79184
rect 339604 79144 339610 79156
rect 343778 79144 343784 79156
rect 343836 79144 343842 79196
rect 344514 79144 344520 79196
rect 344572 79184 344578 79196
rect 344572 79156 346952 79184
rect 344572 79144 344578 79156
rect 65478 79076 65484 79128
rect 65536 79116 65542 79128
rect 69342 79116 69348 79128
rect 65536 79088 69348 79116
rect 65536 79076 65542 79088
rect 69342 79076 69348 79088
rect 69400 79076 69406 79128
rect 154166 79076 154172 79128
rect 154224 79116 154230 79128
rect 158950 79116 158956 79128
rect 154224 79088 158956 79116
rect 154224 79076 154230 79088
rect 158950 79076 158956 79088
rect 159008 79076 159014 79128
rect 249018 79076 249024 79128
rect 249076 79116 249082 79128
rect 256194 79116 256200 79128
rect 249076 79088 256200 79116
rect 249076 79076 249082 79088
rect 256194 79076 256200 79088
rect 256252 79076 256258 79128
rect 338994 79076 339000 79128
rect 339052 79116 339058 79128
rect 342674 79116 342680 79128
rect 339052 79088 342680 79116
rect 339052 79076 339058 79088
rect 342674 79076 342680 79088
rect 342732 79076 342738 79128
rect 344606 79076 344612 79128
rect 344664 79116 344670 79128
rect 346814 79116 346820 79128
rect 344664 79088 346820 79116
rect 344664 79076 344670 79088
rect 346814 79076 346820 79088
rect 346872 79076 346878 79128
rect 346924 79116 346952 79156
rect 347274 79144 347280 79196
rect 347332 79184 347338 79196
rect 349942 79184 349948 79196
rect 347332 79156 349948 79184
rect 347332 79144 347338 79156
rect 349942 79144 349948 79156
rect 350000 79144 350006 79196
rect 347918 79116 347924 79128
rect 346924 79088 347924 79116
rect 347918 79076 347924 79088
rect 347976 79076 347982 79128
rect 57198 79008 57204 79060
rect 57256 79048 57262 79060
rect 61614 79048 61620 79060
rect 57256 79020 61620 79048
rect 57256 79008 57262 79020
rect 61614 79008 61620 79020
rect 61672 79008 61678 79060
rect 154718 79008 154724 79060
rect 154776 79048 154782 79060
rect 160974 79048 160980 79060
rect 154776 79020 160980 79048
rect 154776 79008 154782 79020
rect 160974 79008 160980 79020
rect 161032 79008 161038 79060
rect 337522 79008 337528 79060
rect 337580 79048 337586 79060
rect 338258 79048 338264 79060
rect 337580 79020 338264 79048
rect 337580 79008 337586 79020
rect 338258 79008 338264 79020
rect 338316 79008 338322 79060
rect 341754 79008 341760 79060
rect 341812 79048 341818 79060
rect 344790 79048 344796 79060
rect 341812 79020 344796 79048
rect 341812 79008 341818 79020
rect 344790 79008 344796 79020
rect 344848 79008 344854 79060
rect 62350 78940 62356 78992
rect 62408 78980 62414 78992
rect 64469 78983 64527 78989
rect 64469 78980 64481 78983
rect 62408 78952 64481 78980
rect 62408 78940 62414 78952
rect 64469 78949 64481 78952
rect 64515 78949 64527 78983
rect 151958 78980 151964 78992
rect 64469 78943 64527 78949
rect 151884 78952 151964 78980
rect 58118 78872 58124 78924
rect 58176 78912 58182 78924
rect 63917 78915 63975 78921
rect 63917 78912 63929 78915
rect 58176 78884 63929 78912
rect 58176 78872 58182 78884
rect 63917 78881 63929 78884
rect 63963 78881 63975 78915
rect 63917 78875 63975 78881
rect 64374 78872 64380 78924
rect 64432 78912 64438 78924
rect 68514 78912 68520 78924
rect 64432 78884 68520 78912
rect 64432 78872 64438 78884
rect 68514 78872 68520 78884
rect 68572 78872 68578 78924
rect 63638 78804 63644 78856
rect 63696 78844 63702 78856
rect 74770 78844 74776 78856
rect 63696 78816 74776 78844
rect 63696 78804 63702 78816
rect 74770 78804 74776 78816
rect 74828 78804 74834 78856
rect 62258 78736 62264 78788
rect 62316 78776 62322 78788
rect 67045 78779 67103 78785
rect 67045 78776 67057 78779
rect 62316 78748 67057 78776
rect 62316 78736 62322 78748
rect 67045 78745 67057 78748
rect 67091 78745 67103 78779
rect 67045 78739 67103 78745
rect 67134 78736 67140 78788
rect 67192 78776 67198 78788
rect 71642 78776 71648 78788
rect 67192 78748 71648 78776
rect 67192 78736 67198 78748
rect 71642 78736 71648 78748
rect 71700 78736 71706 78788
rect 151884 78776 151912 78952
rect 151958 78940 151964 78952
rect 152016 78940 152022 78992
rect 154074 78940 154080 78992
rect 154132 78980 154138 78992
rect 160330 78980 160336 78992
rect 154132 78952 160336 78980
rect 154132 78940 154138 78952
rect 160330 78940 160336 78952
rect 160388 78940 160394 78992
rect 244878 78940 244884 78992
rect 244936 78980 244942 78992
rect 252146 78980 252152 78992
rect 244936 78952 252152 78980
rect 244936 78940 244942 78952
rect 252146 78940 252152 78952
rect 252204 78940 252210 78992
rect 153338 78872 153344 78924
rect 153396 78912 153402 78924
rect 162446 78912 162452 78924
rect 153396 78884 162452 78912
rect 153396 78872 153402 78884
rect 162446 78872 162452 78884
rect 162504 78872 162510 78924
rect 247638 78872 247644 78924
rect 247696 78912 247702 78924
rect 256286 78912 256292 78924
rect 247696 78884 256292 78912
rect 247696 78872 247702 78884
rect 256286 78872 256292 78884
rect 256344 78872 256350 78924
rect 151958 78804 151964 78856
rect 152016 78844 152022 78856
rect 161802 78844 161808 78856
rect 152016 78816 161808 78844
rect 152016 78804 152022 78816
rect 161802 78804 161808 78816
rect 161860 78804 161866 78856
rect 246258 78804 246264 78856
rect 246316 78844 246322 78856
rect 255642 78844 255648 78856
rect 246316 78816 255648 78844
rect 246316 78804 246322 78816
rect 255642 78804 255648 78816
rect 255700 78804 255706 78856
rect 163090 78776 163096 78788
rect 151884 78748 163096 78776
rect 163090 78736 163096 78748
rect 163148 78736 163154 78788
rect 245798 78736 245804 78788
rect 245856 78776 245862 78788
rect 256930 78776 256936 78788
rect 245856 78748 256936 78776
rect 245856 78736 245862 78748
rect 256930 78736 256936 78748
rect 256988 78736 256994 78788
rect 60878 78668 60884 78720
rect 60936 78708 60942 78720
rect 72654 78708 72660 78720
rect 60936 78680 72660 78708
rect 60936 78668 60942 78680
rect 72654 78668 72660 78680
rect 72712 78668 72718 78720
rect 153246 78668 153252 78720
rect 153304 78708 153310 78720
rect 164562 78708 164568 78720
rect 153304 78680 164568 78708
rect 153304 78668 153310 78680
rect 164562 78668 164568 78680
rect 164620 78668 164626 78720
rect 247086 78668 247092 78720
rect 247144 78708 247150 78720
rect 258402 78708 258408 78720
rect 247144 78680 258408 78708
rect 247144 78668 247150 78680
rect 258402 78668 258408 78680
rect 258460 78668 258466 78720
rect 339086 78668 339092 78720
rect 339144 78708 339150 78720
rect 341662 78708 341668 78720
rect 339144 78680 341668 78708
rect 339144 78668 339150 78680
rect 341662 78668 341668 78680
rect 341720 78668 341726 78720
rect 59222 78600 59228 78652
rect 59280 78640 59286 78652
rect 63730 78640 63736 78652
rect 59280 78612 63736 78640
rect 59280 78600 59286 78612
rect 63730 78600 63736 78612
rect 63788 78600 63794 78652
rect 70630 78640 70636 78652
rect 63840 78612 70636 78640
rect 59498 78532 59504 78584
rect 59556 78572 59562 78584
rect 63840 78572 63868 78612
rect 70630 78600 70636 78612
rect 70688 78600 70694 78652
rect 153430 78600 153436 78652
rect 153488 78640 153494 78652
rect 165942 78640 165948 78652
rect 153488 78612 165948 78640
rect 153488 78600 153494 78612
rect 165942 78600 165948 78612
rect 166000 78600 166006 78652
rect 248558 78600 248564 78652
rect 248616 78640 248622 78652
rect 261070 78640 261076 78652
rect 248616 78612 261076 78640
rect 248616 78600 248622 78612
rect 261070 78600 261076 78612
rect 261128 78600 261134 78652
rect 338534 78600 338540 78652
rect 338592 78640 338598 78652
rect 345894 78640 345900 78652
rect 338592 78612 345900 78640
rect 338592 78600 338598 78612
rect 345894 78600 345900 78612
rect 345952 78600 345958 78652
rect 59556 78544 63868 78572
rect 63917 78575 63975 78581
rect 59556 78532 59562 78544
rect 63917 78541 63929 78575
rect 63963 78572 63975 78575
rect 69618 78572 69624 78584
rect 63963 78544 69624 78572
rect 63963 78541 63975 78544
rect 63917 78535 63975 78541
rect 69618 78532 69624 78544
rect 69676 78532 69682 78584
rect 154626 78532 154632 78584
rect 154684 78572 154690 78584
rect 167322 78572 167328 78584
rect 154684 78544 167328 78572
rect 154684 78532 154690 78544
rect 167322 78532 167328 78544
rect 167380 78532 167386 78584
rect 247178 78532 247184 78584
rect 247236 78572 247242 78584
rect 259690 78572 259696 78584
rect 247236 78544 259696 78572
rect 247236 78532 247242 78544
rect 259690 78532 259696 78544
rect 259748 78532 259754 78584
rect 55358 78464 55364 78516
rect 55416 78504 55422 78516
rect 66490 78504 66496 78516
rect 55416 78476 66496 78504
rect 55416 78464 55422 78476
rect 66490 78464 66496 78476
rect 66548 78464 66554 78516
rect 67045 78507 67103 78513
rect 67045 78473 67057 78507
rect 67091 78504 67103 78507
rect 73758 78504 73764 78516
rect 67091 78476 73764 78504
rect 67091 78473 67103 78476
rect 67045 78467 67103 78473
rect 73758 78464 73764 78476
rect 73816 78464 73822 78516
rect 154442 78464 154448 78516
rect 154500 78504 154506 78516
rect 168702 78504 168708 78516
rect 154500 78476 168708 78504
rect 154500 78464 154506 78476
rect 168702 78464 168708 78476
rect 168760 78464 168766 78516
rect 248466 78464 248472 78516
rect 248524 78504 248530 78516
rect 262450 78504 262456 78516
rect 248524 78476 262456 78504
rect 248524 78464 248530 78476
rect 262450 78464 262456 78476
rect 262508 78464 262514 78516
rect 63362 78396 63368 78448
rect 63420 78436 63426 78448
rect 67226 78436 67232 78448
rect 63420 78408 67232 78436
rect 63420 78396 63426 78408
rect 67226 78396 67232 78408
rect 67284 78396 67290 78448
rect 58210 78328 58216 78380
rect 58268 78368 58274 78380
rect 63822 78368 63828 78380
rect 58268 78340 63828 78368
rect 58268 78328 58274 78340
rect 63822 78328 63828 78340
rect 63880 78328 63886 78380
rect 156098 78328 156104 78380
rect 156156 78368 156162 78380
rect 162354 78368 162360 78380
rect 156156 78340 162360 78368
rect 156156 78328 156162 78340
rect 162354 78328 162360 78340
rect 162412 78328 162418 78380
rect 250398 78328 250404 78380
rect 250456 78368 250462 78380
rect 257574 78368 257580 78380
rect 250456 78340 257580 78368
rect 250456 78328 250462 78340
rect 257574 78328 257580 78340
rect 257632 78328 257638 78380
rect 61338 78056 61344 78108
rect 61396 78096 61402 78108
rect 65754 78096 65760 78108
rect 61396 78068 65760 78096
rect 61396 78056 61402 78068
rect 65754 78056 65760 78068
rect 65812 78056 65818 78108
rect 427406 77784 427412 77836
rect 427464 77824 427470 77836
rect 429522 77824 429528 77836
rect 427464 77796 429528 77824
rect 427464 77784 427470 77796
rect 429522 77784 429528 77796
rect 429580 77784 429586 77836
rect 88018 76424 88024 76476
rect 88076 76464 88082 76476
rect 88202 76464 88208 76476
rect 88076 76436 88208 76464
rect 88076 76424 88082 76436
rect 88202 76424 88208 76436
rect 88260 76424 88266 76476
rect 358409 76467 358467 76473
rect 358409 76433 358421 76467
rect 358455 76464 358467 76467
rect 358498 76464 358504 76476
rect 358455 76436 358504 76464
rect 358455 76433 358467 76436
rect 358409 76427 358467 76433
rect 358498 76424 358504 76436
rect 358556 76424 358562 76476
rect 79462 76356 79468 76408
rect 79520 76396 79526 76408
rect 123990 76396 123996 76408
rect 79520 76368 123996 76396
rect 79520 76356 79526 76368
rect 123990 76356 123996 76368
rect 124048 76396 124054 76408
rect 139630 76396 139636 76408
rect 124048 76368 139636 76396
rect 124048 76356 124054 76368
rect 139630 76356 139636 76368
rect 139688 76356 139694 76408
rect 173854 76356 173860 76408
rect 173912 76396 173918 76408
rect 218014 76396 218020 76408
rect 173912 76368 218020 76396
rect 173912 76356 173918 76368
rect 218014 76356 218020 76368
rect 218072 76396 218078 76408
rect 233470 76396 233476 76408
rect 218072 76368 233476 76396
rect 218072 76356 218078 76368
rect 233470 76356 233476 76368
rect 233528 76356 233534 76408
rect 266590 76356 266596 76408
rect 266648 76396 266654 76408
rect 312038 76396 312044 76408
rect 266648 76368 312044 76396
rect 266648 76356 266654 76368
rect 312038 76356 312044 76368
rect 312096 76396 312102 76408
rect 328414 76396 328420 76408
rect 312096 76368 328420 76396
rect 312096 76356 312102 76368
rect 328414 76356 328420 76368
rect 328472 76356 328478 76408
rect 80198 73704 80204 73756
rect 80256 73744 80262 73756
rect 87926 73744 87932 73756
rect 80256 73716 87932 73744
rect 80256 73704 80262 73716
rect 87926 73704 87932 73716
rect 87984 73704 87990 73756
rect 174038 73704 174044 73756
rect 174096 73744 174102 73756
rect 181030 73744 181036 73756
rect 174096 73716 181036 73744
rect 174096 73704 174102 73716
rect 181030 73704 181036 73716
rect 181088 73704 181094 73756
rect 226570 73704 226576 73756
rect 226628 73744 226634 73756
rect 233470 73744 233476 73756
rect 226628 73716 233476 73744
rect 226628 73704 226634 73716
rect 233470 73704 233476 73716
rect 233528 73704 233534 73756
rect 266590 73704 266596 73756
rect 266648 73744 266654 73756
rect 274870 73744 274876 73756
rect 266648 73716 274876 73744
rect 266648 73704 266654 73716
rect 274870 73704 274876 73716
rect 274928 73704 274934 73756
rect 304862 73704 304868 73756
rect 304920 73744 304926 73756
rect 305046 73744 305052 73756
rect 304920 73716 305052 73744
rect 304920 73704 304926 73716
rect 305046 73704 305052 73716
rect 305104 73704 305110 73756
rect 321790 73704 321796 73756
rect 321848 73744 321854 73756
rect 328322 73744 328328 73756
rect 321848 73716 328328 73744
rect 321848 73704 321854 73716
rect 328322 73704 328328 73716
rect 328380 73704 328386 73756
rect 110190 73432 110196 73484
rect 110248 73472 110254 73484
rect 116814 73472 116820 73484
rect 110248 73444 116820 73472
rect 110248 73432 110254 73444
rect 116814 73432 116820 73444
rect 116872 73432 116878 73484
rect 204122 72956 204128 73008
rect 204180 72996 204186 73008
rect 210930 72996 210936 73008
rect 204180 72968 210936 72996
rect 204180 72956 204186 72968
rect 210930 72956 210936 72968
rect 210988 72956 210994 73008
rect 217554 72956 217560 73008
rect 217612 72996 217618 73008
rect 224454 72996 224460 73008
rect 217612 72968 224460 72996
rect 217612 72956 217618 72968
rect 224454 72956 224460 72968
rect 224512 72956 224518 73008
rect 311210 72616 311216 72668
rect 311268 72656 311274 72668
rect 318294 72656 318300 72668
rect 311268 72628 318300 72656
rect 311268 72616 311274 72628
rect 318294 72616 318300 72628
rect 318352 72616 318358 72668
rect 79830 72344 79836 72396
rect 79888 72384 79894 72396
rect 85718 72384 85724 72396
rect 79888 72356 85724 72384
rect 79888 72344 79894 72356
rect 85718 72344 85724 72356
rect 85776 72344 85782 72396
rect 123530 72344 123536 72396
rect 123588 72384 123594 72396
rect 130982 72384 130988 72396
rect 123588 72356 130988 72384
rect 123588 72344 123594 72356
rect 130982 72344 130988 72356
rect 131040 72344 131046 72396
rect 172934 72344 172940 72396
rect 172992 72384 172998 72396
rect 180938 72384 180944 72396
rect 172992 72356 180944 72384
rect 172992 72344 172998 72356
rect 180938 72344 180944 72356
rect 180996 72344 181002 72396
rect 230158 72344 230164 72396
rect 230216 72384 230222 72396
rect 233470 72384 233476 72396
rect 230216 72356 233476 72384
rect 230216 72344 230222 72356
rect 233470 72344 233476 72356
rect 233528 72344 233534 72396
rect 266590 72344 266596 72396
rect 266648 72384 266654 72396
rect 274686 72384 274692 72396
rect 266648 72356 274692 72384
rect 266648 72344 266654 72356
rect 274686 72344 274692 72356
rect 274744 72344 274750 72396
rect 284530 72344 284536 72396
rect 284588 72384 284594 72396
rect 285818 72384 285824 72396
rect 284588 72356 285824 72384
rect 284588 72344 284594 72356
rect 285818 72344 285824 72356
rect 285876 72344 285882 72396
rect 297870 72344 297876 72396
rect 297928 72384 297934 72396
rect 304862 72384 304868 72396
rect 297928 72356 304868 72384
rect 297928 72344 297934 72356
rect 304862 72344 304868 72356
rect 304920 72344 304926 72396
rect 78910 70984 78916 71036
rect 78968 71024 78974 71036
rect 85626 71024 85632 71036
rect 78968 70996 85632 71024
rect 78968 70984 78974 70996
rect 85626 70984 85632 70996
rect 85684 70984 85690 71036
rect 174038 70984 174044 71036
rect 174096 71024 174102 71036
rect 178454 71024 178460 71036
rect 174096 70996 178460 71024
rect 174096 70984 174102 70996
rect 178454 70984 178460 70996
rect 178512 70984 178518 71036
rect 266590 70984 266596 71036
rect 266648 71024 266654 71036
rect 272018 71024 272024 71036
rect 266648 70996 272024 71024
rect 266648 70984 266654 70996
rect 272018 70984 272024 70996
rect 272076 70984 272082 71036
rect 132546 70916 132552 70968
rect 132604 70956 132610 70968
rect 139630 70956 139636 70968
rect 132604 70928 139636 70956
rect 132604 70916 132610 70928
rect 139630 70916 139636 70928
rect 139688 70916 139694 70968
rect 173302 70916 173308 70968
rect 173360 70956 173366 70968
rect 178270 70956 178276 70968
rect 173360 70928 178276 70956
rect 173360 70916 173366 70928
rect 178270 70916 178276 70928
rect 178328 70916 178334 70968
rect 230618 70916 230624 70968
rect 230676 70956 230682 70968
rect 233562 70956 233568 70968
rect 230676 70928 233568 70956
rect 230676 70916 230682 70928
rect 233562 70916 233568 70928
rect 233620 70916 233626 70968
rect 266682 70916 266688 70968
rect 266740 70956 266746 70968
rect 274778 70956 274784 70968
rect 266740 70928 274784 70956
rect 266740 70916 266746 70928
rect 274778 70916 274784 70928
rect 274836 70916 274842 70968
rect 321238 70916 321244 70968
rect 321296 70956 321302 70968
rect 328506 70956 328512 70968
rect 321296 70928 328512 70956
rect 321296 70916 321302 70928
rect 328506 70916 328512 70928
rect 328564 70916 328570 70968
rect 174038 69896 174044 69948
rect 174096 69936 174102 69948
rect 178362 69936 178368 69948
rect 174096 69908 178368 69936
rect 174096 69896 174102 69908
rect 178362 69896 178368 69908
rect 178420 69896 178426 69948
rect 358498 69664 358504 69676
rect 358424 69636 358504 69664
rect 80198 69556 80204 69608
rect 80256 69596 80262 69608
rect 87282 69596 87288 69608
rect 80256 69568 87288 69596
rect 80256 69556 80262 69568
rect 87282 69556 87288 69568
rect 87340 69556 87346 69608
rect 266590 69556 266596 69608
rect 266648 69596 266654 69608
rect 274962 69596 274968 69608
rect 266648 69568 274968 69596
rect 266648 69556 266654 69568
rect 274962 69556 274968 69568
rect 275020 69556 275026 69608
rect 358424 69540 358452 69636
rect 358498 69624 358504 69636
rect 358556 69624 358562 69676
rect 131350 69488 131356 69540
rect 131408 69528 131414 69540
rect 139722 69528 139728 69540
rect 131408 69500 139728 69528
rect 131408 69488 131414 69500
rect 139722 69488 139728 69500
rect 139780 69488 139786 69540
rect 225926 69488 225932 69540
rect 225984 69528 225990 69540
rect 230158 69528 230164 69540
rect 225984 69500 230164 69528
rect 225984 69488 225990 69500
rect 230158 69488 230164 69500
rect 230216 69488 230222 69540
rect 358406 69488 358412 69540
rect 358464 69488 358470 69540
rect 131810 69420 131816 69472
rect 131868 69460 131874 69472
rect 139538 69460 139544 69472
rect 131868 69432 139544 69460
rect 131868 69420 131874 69432
rect 139538 69420 139544 69432
rect 139596 69420 139602 69472
rect 321606 69080 321612 69132
rect 321664 69120 321670 69132
rect 327218 69120 327224 69132
rect 321664 69092 327224 69120
rect 321664 69080 321670 69092
rect 327218 69080 327224 69092
rect 327276 69080 327282 69132
rect 85718 68944 85724 68996
rect 85776 68984 85782 68996
rect 87650 68984 87656 68996
rect 85776 68956 87656 68984
rect 85776 68944 85782 68956
rect 87650 68944 87656 68956
rect 87708 68944 87714 68996
rect 79278 68196 79284 68248
rect 79336 68236 79342 68248
rect 85074 68236 85080 68248
rect 79336 68208 85080 68236
rect 79336 68196 79342 68208
rect 85074 68196 85080 68208
rect 85132 68196 85138 68248
rect 136778 68196 136784 68248
rect 136836 68236 136842 68248
rect 139630 68236 139636 68248
rect 136836 68208 139636 68236
rect 136836 68196 136842 68208
rect 139630 68196 139636 68208
rect 139688 68196 139694 68248
rect 172934 68196 172940 68248
rect 172992 68236 172998 68248
rect 180938 68236 180944 68248
rect 172992 68208 180944 68236
rect 172992 68196 172998 68208
rect 180938 68196 180944 68208
rect 180996 68196 181002 68248
rect 266590 68196 266596 68248
rect 266648 68236 266654 68248
rect 274686 68236 274692 68248
rect 266648 68208 274692 68236
rect 266648 68196 266654 68208
rect 274686 68196 274692 68208
rect 274744 68196 274750 68248
rect 85626 68128 85632 68180
rect 85684 68168 85690 68180
rect 87834 68168 87840 68180
rect 85684 68140 87840 68168
rect 85684 68128 85690 68140
rect 87834 68128 87840 68140
rect 87892 68128 87898 68180
rect 132362 68128 132368 68180
rect 132420 68168 132426 68180
rect 139906 68168 139912 68180
rect 132420 68140 139912 68168
rect 132420 68128 132426 68140
rect 139906 68128 139912 68140
rect 139964 68128 139970 68180
rect 178270 68128 178276 68180
rect 178328 68168 178334 68180
rect 181398 68168 181404 68180
rect 178328 68140 181404 68168
rect 178328 68128 178334 68140
rect 181398 68128 181404 68140
rect 181456 68128 181462 68180
rect 226294 68128 226300 68180
rect 226352 68168 226358 68180
rect 233470 68168 233476 68180
rect 226352 68140 233476 68168
rect 226352 68128 226358 68140
rect 233470 68128 233476 68140
rect 233528 68128 233534 68180
rect 79554 67516 79560 67568
rect 79612 67556 79618 67568
rect 129418 67556 129424 67568
rect 79612 67528 129424 67556
rect 79612 67516 79618 67528
rect 129418 67516 129424 67528
rect 129476 67516 129482 67568
rect 173394 67516 173400 67568
rect 173452 67556 173458 67568
rect 223442 67556 223448 67568
rect 173452 67528 223448 67556
rect 173452 67516 173458 67528
rect 223442 67516 223448 67528
rect 223500 67516 223506 67568
rect 267234 67516 267240 67568
rect 267292 67556 267298 67568
rect 317558 67556 317564 67568
rect 267292 67528 317564 67556
rect 267292 67516 267298 67528
rect 317558 67516 317564 67528
rect 317616 67516 317622 67568
rect 80198 67176 80204 67228
rect 80256 67216 80262 67228
rect 82774 67216 82780 67228
rect 80256 67188 82780 67216
rect 80256 67176 80262 67188
rect 82774 67176 82780 67188
rect 82832 67176 82838 67228
rect 321606 67040 321612 67092
rect 321664 67080 321670 67092
rect 327034 67080 327040 67092
rect 321664 67052 327040 67080
rect 321664 67040 321670 67052
rect 327034 67040 327040 67052
rect 327092 67040 327098 67092
rect 174038 66904 174044 66956
rect 174096 66944 174102 66956
rect 179098 66944 179104 66956
rect 174096 66916 179104 66944
rect 174096 66904 174102 66916
rect 179098 66904 179104 66916
rect 179156 66904 179162 66956
rect 135950 66836 135956 66888
rect 136008 66876 136014 66888
rect 139722 66876 139728 66888
rect 136008 66848 139728 66876
rect 136008 66836 136014 66848
rect 139722 66836 139728 66848
rect 139780 66836 139786 66888
rect 266682 66836 266688 66888
rect 266740 66876 266746 66888
rect 272662 66876 272668 66888
rect 266740 66848 272668 66876
rect 266740 66836 266746 66848
rect 272662 66836 272668 66848
rect 272720 66836 272726 66888
rect 80198 66768 80204 66820
rect 80256 66808 80262 66820
rect 87374 66808 87380 66820
rect 80256 66780 87380 66808
rect 80256 66768 80262 66780
rect 87374 66768 87380 66780
rect 87432 66768 87438 66820
rect 136134 66768 136140 66820
rect 136192 66808 136198 66820
rect 139630 66808 139636 66820
rect 136192 66780 139636 66808
rect 136192 66768 136198 66780
rect 139630 66768 139636 66780
rect 139688 66768 139694 66820
rect 173854 66768 173860 66820
rect 173912 66808 173918 66820
rect 181766 66808 181772 66820
rect 173912 66780 181772 66808
rect 173912 66768 173918 66780
rect 181766 66768 181772 66780
rect 181824 66768 181830 66820
rect 266590 66768 266596 66820
rect 266648 66808 266654 66820
rect 274226 66808 274232 66820
rect 266648 66780 274232 66808
rect 266648 66768 266654 66780
rect 274226 66768 274232 66780
rect 274284 66768 274290 66820
rect 80290 66700 80296 66752
rect 80348 66740 80354 66752
rect 87190 66740 87196 66752
rect 80348 66712 87196 66740
rect 80348 66700 80354 66712
rect 87190 66700 87196 66712
rect 87248 66700 87254 66752
rect 88202 66740 88208 66752
rect 88163 66712 88208 66740
rect 88202 66700 88208 66712
rect 88260 66700 88266 66752
rect 132362 66700 132368 66752
rect 132420 66740 132426 66752
rect 139814 66740 139820 66752
rect 132420 66712 139820 66740
rect 132420 66700 132426 66712
rect 139814 66700 139820 66712
rect 139872 66700 139878 66752
rect 226386 66700 226392 66752
rect 226444 66740 226450 66752
rect 233562 66740 233568 66752
rect 226444 66712 233568 66740
rect 226444 66700 226450 66712
rect 233562 66700 233568 66712
rect 233620 66700 233626 66752
rect 272018 66700 272024 66752
rect 272076 66740 272082 66752
rect 274870 66740 274876 66752
rect 272076 66712 274876 66740
rect 272076 66700 272082 66712
rect 274870 66700 274876 66712
rect 274928 66700 274934 66752
rect 317374 66700 317380 66752
rect 317432 66740 317438 66752
rect 317561 66743 317619 66749
rect 317561 66740 317573 66743
rect 317432 66712 317573 66740
rect 317432 66700 317438 66712
rect 317561 66709 317573 66712
rect 317607 66709 317619 66743
rect 317561 66703 317619 66709
rect 226294 66632 226300 66684
rect 226352 66672 226358 66684
rect 230618 66672 230624 66684
rect 226352 66644 230624 66672
rect 226352 66632 226358 66644
rect 230618 66632 230624 66644
rect 230676 66632 230682 66684
rect 178362 66428 178368 66480
rect 178420 66468 178426 66480
rect 182134 66468 182140 66480
rect 178420 66440 182140 66468
rect 178420 66428 178426 66440
rect 182134 66428 182140 66440
rect 182192 66428 182198 66480
rect 178454 66156 178460 66208
rect 178512 66196 178518 66208
rect 181950 66196 181956 66208
rect 178512 66168 181956 66196
rect 178512 66156 178518 66168
rect 181950 66156 181956 66168
rect 182008 66156 182014 66208
rect 321606 65952 321612 66004
rect 321664 65992 321670 66004
rect 327126 65992 327132 66004
rect 321664 65964 327132 65992
rect 321664 65952 321670 65964
rect 327126 65952 327132 65964
rect 327184 65952 327190 66004
rect 173854 65680 173860 65732
rect 173912 65720 173918 65732
rect 178822 65720 178828 65732
rect 173912 65692 178828 65720
rect 173912 65680 173918 65692
rect 178822 65680 178828 65692
rect 178880 65680 178886 65732
rect 80198 65408 80204 65460
rect 80256 65448 80262 65460
rect 87282 65448 87288 65460
rect 80256 65420 87288 65448
rect 80256 65408 80262 65420
rect 87282 65408 87288 65420
rect 87340 65408 87346 65460
rect 266590 65408 266596 65460
rect 266648 65448 266654 65460
rect 274778 65448 274784 65460
rect 266648 65420 274784 65448
rect 266648 65408 266654 65420
rect 274778 65408 274784 65420
rect 274836 65408 274842 65460
rect 82774 65340 82780 65392
rect 82832 65380 82838 65392
rect 87190 65380 87196 65392
rect 82832 65352 87196 65380
rect 82832 65340 82838 65352
rect 87190 65340 87196 65352
rect 87248 65340 87254 65392
rect 131350 65340 131356 65392
rect 131408 65380 131414 65392
rect 136778 65380 136784 65392
rect 131408 65352 136784 65380
rect 131408 65340 131414 65352
rect 136778 65340 136784 65352
rect 136836 65340 136842 65392
rect 225926 65340 225932 65392
rect 225984 65380 225990 65392
rect 233470 65380 233476 65392
rect 225984 65352 233476 65380
rect 225984 65340 225990 65352
rect 233470 65340 233476 65352
rect 233528 65340 233534 65392
rect 272662 65340 272668 65392
rect 272720 65380 272726 65392
rect 274870 65380 274876 65392
rect 272720 65352 274876 65380
rect 272720 65340 272726 65352
rect 274870 65340 274876 65352
rect 274928 65340 274934 65392
rect 85074 65272 85080 65324
rect 85132 65312 85138 65324
rect 87466 65312 87472 65324
rect 85132 65284 87472 65312
rect 85132 65272 85138 65284
rect 87466 65272 87472 65284
rect 87524 65272 87530 65324
rect 132178 65272 132184 65324
rect 132236 65312 132242 65324
rect 135950 65312 135956 65324
rect 132236 65284 135956 65312
rect 132236 65272 132242 65284
rect 135950 65272 135956 65284
rect 136008 65272 136014 65324
rect 226202 65272 226208 65324
rect 226260 65312 226266 65324
rect 233654 65312 233660 65324
rect 226260 65284 233660 65312
rect 226260 65272 226266 65284
rect 233654 65272 233660 65284
rect 233712 65272 233718 65324
rect 173486 64864 173492 64916
rect 173544 64904 173550 64916
rect 175878 64904 175884 64916
rect 173544 64876 175884 64904
rect 173544 64864 173550 64876
rect 175878 64864 175884 64876
rect 175936 64864 175942 64916
rect 321606 64592 321612 64644
rect 321664 64632 321670 64644
rect 327218 64632 327224 64644
rect 321664 64604 327224 64632
rect 321664 64592 321670 64604
rect 327218 64592 327224 64604
rect 327276 64592 327282 64644
rect 79462 64456 79468 64508
rect 79520 64496 79526 64508
rect 82406 64496 82412 64508
rect 79520 64468 82412 64496
rect 79520 64456 79526 64468
rect 82406 64456 82412 64468
rect 82464 64456 82470 64508
rect 229422 64320 229428 64372
rect 229480 64360 229486 64372
rect 233470 64360 233476 64372
rect 229480 64332 233476 64360
rect 229480 64320 229486 64332
rect 233470 64320 233476 64332
rect 233528 64320 233534 64372
rect 321606 64116 321612 64168
rect 321664 64156 321670 64168
rect 328230 64156 328236 64168
rect 321664 64128 328236 64156
rect 321664 64116 321670 64128
rect 328230 64116 328236 64128
rect 328288 64116 328294 64168
rect 266590 64048 266596 64100
rect 266648 64088 266654 64100
rect 273398 64088 273404 64100
rect 266648 64060 273404 64088
rect 266648 64048 266654 64060
rect 273398 64048 273404 64060
rect 273456 64048 273462 64100
rect 132362 63980 132368 64032
rect 132420 64020 132426 64032
rect 136134 64020 136140 64032
rect 132420 63992 136140 64020
rect 132420 63980 132426 63992
rect 136134 63980 136140 63992
rect 136192 63980 136198 64032
rect 179098 63980 179104 64032
rect 179156 64020 179162 64032
rect 182318 64020 182324 64032
rect 179156 63992 182324 64020
rect 179156 63980 179162 63992
rect 182318 63980 182324 63992
rect 182376 63980 182382 64032
rect 225742 63980 225748 64032
rect 225800 64020 225806 64032
rect 234206 64020 234212 64032
rect 225800 63992 234212 64020
rect 225800 63980 225806 63992
rect 234206 63980 234212 63992
rect 234264 63980 234270 64032
rect 320502 63640 320508 63692
rect 320560 63680 320566 63692
rect 326942 63680 326948 63692
rect 320560 63652 326948 63680
rect 320560 63640 320566 63652
rect 326942 63640 326948 63652
rect 327000 63640 327006 63692
rect 80198 62960 80204 63012
rect 80256 63000 80262 63012
rect 82590 63000 82596 63012
rect 80256 62972 82596 63000
rect 80256 62960 80262 62972
rect 82590 62960 82596 62972
rect 82648 62960 82654 63012
rect 80198 62688 80204 62740
rect 80256 62728 80262 62740
rect 85718 62728 85724 62740
rect 80256 62700 85724 62728
rect 80256 62688 80262 62700
rect 85718 62688 85724 62700
rect 85776 62688 85782 62740
rect 174038 62688 174044 62740
rect 174096 62728 174102 62740
rect 178270 62728 178276 62740
rect 174096 62700 178276 62728
rect 174096 62688 174102 62700
rect 178270 62688 178276 62700
rect 178328 62688 178334 62740
rect 266590 62688 266596 62740
rect 266648 62728 266654 62740
rect 272846 62728 272852 62740
rect 266648 62700 272852 62728
rect 266648 62688 266654 62700
rect 272846 62688 272852 62700
rect 272904 62688 272910 62740
rect 173486 62620 173492 62672
rect 173544 62660 173550 62672
rect 175602 62660 175608 62672
rect 173544 62632 175608 62660
rect 173544 62620 173550 62632
rect 175602 62620 175608 62632
rect 175660 62620 175666 62672
rect 230434 62620 230440 62672
rect 230492 62660 230498 62672
rect 233470 62660 233476 62672
rect 230492 62632 233476 62660
rect 230492 62620 230498 62632
rect 233470 62620 233476 62632
rect 233528 62620 233534 62672
rect 266682 62620 266688 62672
rect 266740 62660 266746 62672
rect 274870 62660 274876 62672
rect 266740 62632 274876 62660
rect 266740 62620 266746 62632
rect 274870 62620 274876 62632
rect 274928 62620 274934 62672
rect 82406 62552 82412 62604
rect 82464 62592 82470 62604
rect 87190 62592 87196 62604
rect 82464 62564 87196 62592
rect 82464 62552 82470 62564
rect 87190 62552 87196 62564
rect 87248 62552 87254 62604
rect 131718 62552 131724 62604
rect 131776 62592 131782 62604
rect 139630 62592 139636 62604
rect 131776 62564 139636 62592
rect 131776 62552 131782 62564
rect 139630 62552 139636 62564
rect 139688 62552 139694 62604
rect 175878 62552 175884 62604
rect 175936 62592 175942 62604
rect 181582 62592 181588 62604
rect 175936 62564 181588 62592
rect 175936 62552 175942 62564
rect 181582 62552 181588 62564
rect 181640 62552 181646 62604
rect 226294 62552 226300 62604
rect 226352 62592 226358 62604
rect 234390 62592 234396 62604
rect 226352 62564 234396 62592
rect 226352 62552 226358 62564
rect 234390 62552 234396 62564
rect 234448 62552 234454 62604
rect 273398 62552 273404 62604
rect 273456 62592 273462 62604
rect 274962 62592 274968 62604
rect 273456 62564 274968 62592
rect 273456 62552 273462 62564
rect 274962 62552 274968 62564
rect 275020 62552 275026 62604
rect 321054 62552 321060 62604
rect 321112 62592 321118 62604
rect 327126 62592 327132 62604
rect 321112 62564 327132 62592
rect 321112 62552 321118 62564
rect 327126 62552 327132 62564
rect 327184 62552 327190 62604
rect 131350 62484 131356 62536
rect 131408 62524 131414 62536
rect 139906 62524 139912 62536
rect 131408 62496 139912 62524
rect 131408 62484 131414 62496
rect 139906 62484 139912 62496
rect 139964 62484 139970 62536
rect 178822 62484 178828 62536
rect 178880 62524 178886 62536
rect 182318 62524 182324 62536
rect 178880 62496 182324 62524
rect 178880 62484 178886 62496
rect 182318 62484 182324 62496
rect 182376 62484 182382 62536
rect 173118 61600 173124 61652
rect 173176 61640 173182 61652
rect 175510 61640 175516 61652
rect 173176 61612 175516 61640
rect 173176 61600 173182 61612
rect 175510 61600 175516 61612
rect 175568 61600 175574 61652
rect 320686 61532 320692 61584
rect 320744 61572 320750 61584
rect 327310 61572 327316 61584
rect 320744 61544 327316 61572
rect 320744 61532 320750 61544
rect 327310 61532 327316 61544
rect 327368 61532 327374 61584
rect 226294 61396 226300 61448
rect 226352 61436 226358 61448
rect 229422 61436 229428 61448
rect 226352 61408 229428 61436
rect 226352 61396 226358 61408
rect 229422 61396 229428 61408
rect 229480 61396 229486 61448
rect 80198 61328 80204 61380
rect 80256 61368 80262 61380
rect 81670 61368 81676 61380
rect 80256 61340 81676 61368
rect 80256 61328 80262 61340
rect 81670 61328 81676 61340
rect 81728 61328 81734 61380
rect 230526 61260 230532 61312
rect 230584 61300 230590 61312
rect 233470 61300 233476 61312
rect 230584 61272 233476 61300
rect 230584 61260 230590 61272
rect 233470 61260 233476 61272
rect 233528 61260 233534 61312
rect 266590 61260 266596 61312
rect 266648 61300 266654 61312
rect 272754 61300 272760 61312
rect 266648 61272 272760 61300
rect 266648 61260 266654 61272
rect 272754 61260 272760 61272
rect 272812 61260 272818 61312
rect 82590 61192 82596 61244
rect 82648 61232 82654 61244
rect 87190 61232 87196 61244
rect 82648 61204 87196 61232
rect 82648 61192 82654 61204
rect 87190 61192 87196 61204
rect 87248 61192 87254 61244
rect 131350 61192 131356 61244
rect 131408 61232 131414 61244
rect 139722 61232 139728 61244
rect 131408 61204 139728 61232
rect 131408 61192 131414 61204
rect 139722 61192 139728 61204
rect 139780 61192 139786 61244
rect 175602 61192 175608 61244
rect 175660 61232 175666 61244
rect 181214 61232 181220 61244
rect 175660 61204 181220 61232
rect 175660 61192 175666 61204
rect 181214 61192 181220 61204
rect 181272 61192 181278 61244
rect 225742 61192 225748 61244
rect 225800 61232 225806 61244
rect 230434 61232 230440 61244
rect 225800 61204 230440 61232
rect 225800 61192 225806 61204
rect 230434 61192 230440 61204
rect 230492 61192 230498 61244
rect 173118 60512 173124 60564
rect 173176 60552 173182 60564
rect 175786 60552 175792 60564
rect 173176 60524 175792 60552
rect 173176 60512 173182 60524
rect 175786 60512 175792 60524
rect 175844 60512 175850 60564
rect 321054 60240 321060 60292
rect 321112 60280 321118 60292
rect 328414 60280 328420 60292
rect 321112 60252 328420 60280
rect 321112 60240 321118 60252
rect 328414 60240 328420 60252
rect 328472 60240 328478 60292
rect 80198 60104 80204 60156
rect 80256 60144 80262 60156
rect 81762 60144 81768 60156
rect 80256 60116 81768 60144
rect 80256 60104 80262 60116
rect 81762 60104 81768 60116
rect 81820 60104 81826 60156
rect 230618 59900 230624 59952
rect 230676 59940 230682 59952
rect 233470 59940 233476 59952
rect 230676 59912 233476 59940
rect 230676 59900 230682 59912
rect 233470 59900 233476 59912
rect 233528 59900 233534 59952
rect 266590 59900 266596 59952
rect 266648 59940 266654 59952
rect 272662 59940 272668 59952
rect 266648 59912 272668 59940
rect 266648 59900 266654 59912
rect 272662 59900 272668 59912
rect 272720 59900 272726 59952
rect 131350 59832 131356 59884
rect 131408 59872 131414 59884
rect 139814 59872 139820 59884
rect 131408 59844 139820 59872
rect 131408 59832 131414 59844
rect 139814 59832 139820 59844
rect 139872 59832 139878 59884
rect 175510 59832 175516 59884
rect 175568 59872 175574 59884
rect 181122 59872 181128 59884
rect 175568 59844 181128 59872
rect 175568 59832 175574 59844
rect 181122 59832 181128 59844
rect 181180 59832 181186 59884
rect 226294 59832 226300 59884
rect 226352 59872 226358 59884
rect 233562 59872 233568 59884
rect 226352 59844 233568 59872
rect 226352 59832 226358 59844
rect 233562 59832 233568 59844
rect 233620 59832 233626 59884
rect 272754 59832 272760 59884
rect 272812 59872 272818 59884
rect 275422 59872 275428 59884
rect 272812 59844 275428 59872
rect 272812 59832 272818 59844
rect 275422 59832 275428 59844
rect 275480 59832 275486 59884
rect 358406 59832 358412 59884
rect 358464 59872 358470 59884
rect 358590 59872 358596 59884
rect 358464 59844 358596 59872
rect 358464 59832 358470 59844
rect 358590 59832 358596 59844
rect 358648 59832 358654 59884
rect 131442 59764 131448 59816
rect 131500 59804 131506 59816
rect 139630 59804 139636 59816
rect 131500 59776 139636 59804
rect 131500 59764 131506 59776
rect 139630 59764 139636 59776
rect 139688 59764 139694 59816
rect 272846 59764 272852 59816
rect 272904 59804 272910 59816
rect 275698 59804 275704 59816
rect 272904 59776 275704 59804
rect 272904 59764 272910 59776
rect 275698 59764 275704 59776
rect 275756 59764 275762 59816
rect 85718 59696 85724 59748
rect 85776 59736 85782 59748
rect 87834 59736 87840 59748
rect 85776 59708 87840 59736
rect 85776 59696 85782 59708
rect 87834 59696 87840 59708
rect 87892 59696 87898 59748
rect 178270 59696 178276 59748
rect 178328 59736 178334 59748
rect 181030 59736 181036 59748
rect 178328 59708 181036 59736
rect 178328 59696 178334 59708
rect 181030 59696 181036 59708
rect 181088 59696 181094 59748
rect 81670 59492 81676 59544
rect 81728 59532 81734 59544
rect 87190 59532 87196 59544
rect 81728 59504 87196 59532
rect 81728 59492 81734 59504
rect 87190 59492 87196 59504
rect 87248 59492 87254 59544
rect 225742 59424 225748 59476
rect 225800 59464 225806 59476
rect 230526 59464 230532 59476
rect 225800 59436 230532 59464
rect 225800 59424 225806 59436
rect 230526 59424 230532 59436
rect 230584 59424 230590 59476
rect 173026 58744 173032 58796
rect 173084 58784 173090 58796
rect 175694 58784 175700 58796
rect 173084 58756 175700 58784
rect 173084 58744 173090 58756
rect 175694 58744 175700 58756
rect 175752 58744 175758 58796
rect 320502 58676 320508 58728
rect 320560 58716 320566 58728
rect 327218 58716 327224 58728
rect 320560 58688 327224 58716
rect 320560 58676 320566 58688
rect 327218 58676 327224 58688
rect 327276 58676 327282 58728
rect 79646 58608 79652 58660
rect 79704 58648 79710 58660
rect 82958 58648 82964 58660
rect 79704 58620 82964 58648
rect 79704 58608 79710 58620
rect 82958 58608 82964 58620
rect 83016 58608 83022 58660
rect 173578 58608 173584 58660
rect 173636 58648 173642 58660
rect 175602 58648 175608 58660
rect 173636 58620 175608 58648
rect 173636 58608 173642 58620
rect 175602 58608 175608 58620
rect 175660 58608 175666 58660
rect 267878 58608 267884 58660
rect 267936 58648 267942 58660
rect 272110 58648 272116 58660
rect 267936 58620 272116 58648
rect 267936 58608 267942 58620
rect 272110 58608 272116 58620
rect 272168 58608 272174 58660
rect 80198 58540 80204 58592
rect 80256 58580 80262 58592
rect 82406 58580 82412 58592
rect 80256 58552 82412 58580
rect 80256 58540 80262 58552
rect 82406 58540 82412 58552
rect 82464 58540 82470 58592
rect 267326 58540 267332 58592
rect 267384 58580 267390 58592
rect 272294 58580 272300 58592
rect 267384 58552 272300 58580
rect 267384 58540 267390 58552
rect 272294 58540 272300 58552
rect 272352 58540 272358 58592
rect 320410 58540 320416 58592
rect 320468 58580 320474 58592
rect 328322 58580 328328 58592
rect 320468 58552 328328 58580
rect 320468 58540 320474 58552
rect 328322 58540 328328 58552
rect 328380 58540 328386 58592
rect 81762 58472 81768 58524
rect 81820 58512 81826 58524
rect 87190 58512 87196 58524
rect 81820 58484 87196 58512
rect 81820 58472 81826 58484
rect 87190 58472 87196 58484
rect 87248 58472 87254 58524
rect 131350 58472 131356 58524
rect 131408 58512 131414 58524
rect 139722 58512 139728 58524
rect 131408 58484 139728 58512
rect 131408 58472 131414 58484
rect 139722 58472 139728 58484
rect 139780 58472 139786 58524
rect 175786 58472 175792 58524
rect 175844 58512 175850 58524
rect 181030 58512 181036 58524
rect 175844 58484 181036 58512
rect 175844 58472 175850 58484
rect 181030 58472 181036 58484
rect 181088 58472 181094 58524
rect 225558 58472 225564 58524
rect 225616 58512 225622 58524
rect 230618 58512 230624 58524
rect 225616 58484 230624 58512
rect 225616 58472 225622 58484
rect 230618 58472 230624 58484
rect 230676 58472 230682 58524
rect 272662 58472 272668 58524
rect 272720 58512 272726 58524
rect 275698 58512 275704 58524
rect 272720 58484 275704 58512
rect 272720 58472 272726 58484
rect 275698 58472 275704 58484
rect 275756 58472 275762 58524
rect 320410 57792 320416 57844
rect 320468 57832 320474 57844
rect 328414 57832 328420 57844
rect 320468 57804 328420 57832
rect 320468 57792 320474 57804
rect 328414 57792 328420 57804
rect 328472 57792 328478 57844
rect 267694 57384 267700 57436
rect 267752 57424 267758 57436
rect 272202 57424 272208 57436
rect 267752 57396 272208 57424
rect 267752 57384 267758 57396
rect 272202 57384 272208 57396
rect 272260 57384 272266 57436
rect 80198 57112 80204 57164
rect 80256 57152 80262 57164
rect 81854 57152 81860 57164
rect 80256 57124 81860 57152
rect 80256 57112 80262 57124
rect 81854 57112 81860 57124
rect 81912 57112 81918 57164
rect 88205 57155 88263 57161
rect 88205 57121 88217 57155
rect 88251 57152 88263 57155
rect 88294 57152 88300 57164
rect 88251 57124 88300 57152
rect 88251 57121 88263 57124
rect 88205 57115 88263 57121
rect 88294 57112 88300 57124
rect 88352 57112 88358 57164
rect 173302 57112 173308 57164
rect 173360 57152 173366 57164
rect 175510 57152 175516 57164
rect 173360 57124 175516 57152
rect 173360 57112 173366 57124
rect 175510 57112 175516 57124
rect 175568 57112 175574 57164
rect 317558 57152 317564 57164
rect 317519 57124 317564 57152
rect 317558 57112 317564 57124
rect 317616 57112 317622 57164
rect 82958 57044 82964 57096
rect 83016 57084 83022 57096
rect 87190 57084 87196 57096
rect 83016 57056 87196 57084
rect 83016 57044 83022 57056
rect 87190 57044 87196 57056
rect 87248 57044 87254 57096
rect 132178 57044 132184 57096
rect 132236 57084 132242 57096
rect 140366 57084 140372 57096
rect 132236 57056 140372 57084
rect 132236 57044 132242 57056
rect 140366 57044 140372 57056
rect 140424 57044 140430 57096
rect 226294 57044 226300 57096
rect 226352 57084 226358 57096
rect 233654 57084 233660 57096
rect 226352 57056 233660 57084
rect 226352 57044 226358 57056
rect 233654 57044 233660 57056
rect 233712 57044 233718 57096
rect 272294 57044 272300 57096
rect 272352 57084 272358 57096
rect 275698 57084 275704 57096
rect 272352 57056 275704 57084
rect 272352 57044 272358 57056
rect 275698 57044 275704 57056
rect 275756 57044 275762 57096
rect 82406 56976 82412 57028
rect 82464 57016 82470 57028
rect 87282 57016 87288 57028
rect 82464 56988 87288 57016
rect 82464 56976 82470 56988
rect 87282 56976 87288 56988
rect 87340 56976 87346 57028
rect 131350 56976 131356 57028
rect 131408 57016 131414 57028
rect 140458 57016 140464 57028
rect 131408 56988 140464 57016
rect 131408 56976 131414 56988
rect 140458 56976 140464 56988
rect 140516 56976 140522 57028
rect 225650 56976 225656 57028
rect 225708 57016 225714 57028
rect 233470 57016 233476 57028
rect 225708 56988 233476 57016
rect 225708 56976 225714 56988
rect 233470 56976 233476 56988
rect 233528 56976 233534 57028
rect 272110 56976 272116 57028
rect 272168 57016 272174 57028
rect 275238 57016 275244 57028
rect 272168 56988 275244 57016
rect 272168 56976 272174 56988
rect 275238 56976 275244 56988
rect 275296 56976 275302 57028
rect 175602 56568 175608 56620
rect 175660 56608 175666 56620
rect 181122 56608 181128 56620
rect 175660 56580 181128 56608
rect 175660 56568 175666 56580
rect 181122 56568 181128 56580
rect 181180 56568 181186 56620
rect 175694 56500 175700 56552
rect 175752 56540 175758 56552
rect 181030 56540 181036 56552
rect 175752 56512 181036 56540
rect 175752 56500 175758 56512
rect 181030 56500 181036 56512
rect 181088 56500 181094 56552
rect 320410 56500 320416 56552
rect 320468 56540 320474 56552
rect 327494 56540 327500 56552
rect 320468 56512 327500 56540
rect 320468 56500 320474 56512
rect 327494 56500 327500 56512
rect 327552 56500 327558 56552
rect 320502 56296 320508 56348
rect 320560 56336 320566 56348
rect 328598 56336 328604 56348
rect 320560 56308 328604 56336
rect 320560 56296 320566 56308
rect 328598 56296 328604 56308
rect 328656 56296 328662 56348
rect 173486 56024 173492 56076
rect 173544 56064 173550 56076
rect 175602 56064 175608 56076
rect 173544 56036 175608 56064
rect 173544 56024 173550 56036
rect 175602 56024 175608 56036
rect 175660 56024 175666 56076
rect 78910 55752 78916 55804
rect 78968 55792 78974 55804
rect 82958 55792 82964 55804
rect 78968 55764 82964 55792
rect 78968 55752 78974 55764
rect 82958 55752 82964 55764
rect 83016 55752 83022 55804
rect 136502 55752 136508 55804
rect 136560 55792 136566 55804
rect 140458 55792 140464 55804
rect 136560 55764 140464 55792
rect 136560 55752 136566 55764
rect 140458 55752 140464 55764
rect 140516 55752 140522 55804
rect 226478 55752 226484 55804
rect 226536 55792 226542 55804
rect 233470 55792 233476 55804
rect 226536 55764 233476 55792
rect 226536 55752 226542 55764
rect 233470 55752 233476 55764
rect 233528 55752 233534 55804
rect 267326 55752 267332 55804
rect 267384 55792 267390 55804
rect 272110 55792 272116 55804
rect 267384 55764 272116 55792
rect 267384 55752 267390 55764
rect 272110 55752 272116 55764
rect 272168 55752 272174 55804
rect 13130 55684 13136 55736
rect 13188 55724 13194 55736
rect 16350 55724 16356 55736
rect 13188 55696 16356 55724
rect 13188 55684 13194 55696
rect 16350 55684 16356 55696
rect 16408 55684 16414 55736
rect 81854 55684 81860 55736
rect 81912 55724 81918 55736
rect 87190 55724 87196 55736
rect 81912 55696 87196 55724
rect 81912 55684 81918 55696
rect 87190 55684 87196 55696
rect 87248 55684 87254 55736
rect 131350 55684 131356 55736
rect 131408 55724 131414 55736
rect 140274 55724 140280 55736
rect 131408 55696 140280 55724
rect 131408 55684 131414 55696
rect 140274 55684 140280 55696
rect 140332 55684 140338 55736
rect 175510 55684 175516 55736
rect 175568 55724 175574 55736
rect 181030 55724 181036 55736
rect 175568 55696 181036 55724
rect 175568 55684 175574 55696
rect 181030 55684 181036 55696
rect 181088 55684 181094 55736
rect 226386 55684 226392 55736
rect 226444 55724 226450 55736
rect 233562 55724 233568 55736
rect 226444 55696 233568 55724
rect 226444 55684 226450 55696
rect 233562 55684 233568 55696
rect 233620 55684 233626 55736
rect 272202 55684 272208 55736
rect 272260 55724 272266 55736
rect 275422 55724 275428 55736
rect 272260 55696 275428 55724
rect 272260 55684 272266 55696
rect 275422 55684 275428 55696
rect 275480 55684 275486 55736
rect 320410 55616 320416 55668
rect 320468 55656 320474 55668
rect 328414 55656 328420 55668
rect 320468 55628 328420 55656
rect 320468 55616 320474 55628
rect 328414 55616 328420 55628
rect 328472 55616 328478 55668
rect 129418 55004 129424 55056
rect 129476 55044 129482 55056
rect 140642 55044 140648 55056
rect 129476 55016 140648 55044
rect 129476 55004 129482 55016
rect 140642 55004 140648 55016
rect 140700 55004 140706 55056
rect 223442 55004 223448 55056
rect 223500 55044 223506 55056
rect 233470 55044 233476 55056
rect 223500 55016 233476 55044
rect 223500 55004 223506 55016
rect 233470 55004 233476 55016
rect 233528 55004 233534 55056
rect 317469 55047 317527 55053
rect 317469 55013 317481 55047
rect 317515 55044 317527 55047
rect 317558 55044 317564 55056
rect 317515 55016 317564 55044
rect 317515 55013 317527 55016
rect 317469 55007 317527 55013
rect 317558 55004 317564 55016
rect 317616 55044 317622 55056
rect 328506 55044 328512 55056
rect 317616 55016 328512 55044
rect 317616 55004 317622 55016
rect 328506 55004 328512 55016
rect 328564 55004 328570 55056
rect 80198 54392 80204 54444
rect 80256 54432 80262 54444
rect 80256 54404 87328 54432
rect 80256 54392 80262 54404
rect 82958 54256 82964 54308
rect 83016 54296 83022 54308
rect 87190 54296 87196 54308
rect 83016 54268 87196 54296
rect 83016 54256 83022 54268
rect 87190 54256 87196 54268
rect 87248 54256 87254 54308
rect 87300 54296 87328 54404
rect 134110 54392 134116 54444
rect 134168 54432 134174 54444
rect 140366 54432 140372 54444
rect 134168 54404 140372 54432
rect 134168 54392 134174 54404
rect 140366 54392 140372 54404
rect 140424 54392 140430 54444
rect 173578 54392 173584 54444
rect 173636 54432 173642 54444
rect 233470 54432 233476 54444
rect 173636 54404 181720 54432
rect 173636 54392 173642 54404
rect 131350 54324 131356 54376
rect 131408 54364 131414 54376
rect 136502 54364 136508 54376
rect 131408 54336 136508 54364
rect 131408 54324 131414 54336
rect 136502 54324 136508 54336
rect 136560 54324 136566 54376
rect 134110 54296 134116 54308
rect 87300 54268 134116 54296
rect 123548 54172 123576 54268
rect 134110 54256 134116 54268
rect 134168 54256 134174 54308
rect 181692 54296 181720 54404
rect 229348 54404 233476 54432
rect 229348 54296 229376 54404
rect 233470 54392 233476 54404
rect 233528 54392 233534 54444
rect 267878 54392 267884 54444
rect 267936 54432 267942 54444
rect 328414 54432 328420 54444
rect 267936 54404 275836 54432
rect 267936 54392 267942 54404
rect 272110 54324 272116 54376
rect 272168 54364 272174 54376
rect 275698 54364 275704 54376
rect 272168 54336 275704 54364
rect 272168 54324 272174 54336
rect 275698 54324 275704 54336
rect 275756 54324 275762 54376
rect 181692 54268 229376 54296
rect 275808 54296 275836 54404
rect 323832 54404 328420 54432
rect 323832 54296 323860 54404
rect 328414 54392 328420 54404
rect 328472 54392 328478 54444
rect 275808 54268 323860 54296
rect 175602 54188 175608 54240
rect 175660 54228 175666 54240
rect 181030 54228 181036 54240
rect 175660 54200 181036 54228
rect 175660 54188 175666 54200
rect 181030 54188 181036 54200
rect 181088 54188 181094 54240
rect 217572 54172 217600 54268
rect 311596 54172 311624 54268
rect 369170 54256 369176 54308
rect 369228 54296 369234 54308
rect 369538 54296 369544 54308
rect 369228 54268 369544 54296
rect 369228 54256 369234 54268
rect 369538 54256 369544 54268
rect 369596 54256 369602 54308
rect 320410 54188 320416 54240
rect 320468 54228 320474 54240
rect 327494 54228 327500 54240
rect 320468 54200 327500 54228
rect 320468 54188 320474 54200
rect 327494 54188 327500 54200
rect 327552 54188 327558 54240
rect 123530 54120 123536 54172
rect 123588 54120 123594 54172
rect 217554 54120 217560 54172
rect 217612 54120 217618 54172
rect 311578 54120 311584 54172
rect 311636 54120 311642 54172
rect 80198 53644 80204 53696
rect 80256 53684 80262 53696
rect 118654 53684 118660 53696
rect 80256 53656 118660 53684
rect 80256 53644 80262 53656
rect 118654 53644 118660 53656
rect 118712 53684 118718 53696
rect 140550 53684 140556 53696
rect 118712 53656 140556 53684
rect 118712 53644 118718 53656
rect 140550 53644 140556 53656
rect 140608 53644 140614 53696
rect 173578 53644 173584 53696
rect 173636 53684 173642 53696
rect 212494 53684 212500 53696
rect 173636 53656 212500 53684
rect 173636 53644 173642 53656
rect 212494 53644 212500 53656
rect 212552 53684 212558 53696
rect 233470 53684 233476 53696
rect 212552 53656 233476 53684
rect 212552 53644 212558 53656
rect 233470 53644 233476 53656
rect 233528 53644 233534 53696
rect 267878 53644 267884 53696
rect 267936 53684 267942 53696
rect 306610 53684 306616 53696
rect 267936 53656 306616 53684
rect 267936 53644 267942 53656
rect 306610 53644 306616 53656
rect 306668 53684 306674 53696
rect 328414 53684 328420 53696
rect 306668 53656 328420 53684
rect 306668 53644 306674 53656
rect 328414 53644 328420 53656
rect 328472 53644 328478 53696
rect 193453 53347 193511 53353
rect 193453 53313 193465 53347
rect 193499 53344 193511 53347
rect 203021 53347 203079 53353
rect 203021 53344 203033 53347
rect 193499 53316 203033 53344
rect 193499 53313 193511 53316
rect 193453 53307 193511 53313
rect 203021 53313 203033 53316
rect 203067 53313 203079 53347
rect 203021 53307 203079 53313
rect 205781 53347 205839 53353
rect 205781 53313 205793 53347
rect 205827 53344 205839 53347
rect 205827 53316 207940 53344
rect 205827 53313 205839 53316
rect 205781 53307 205839 53313
rect 207912 53288 207940 53316
rect 207894 53236 207900 53288
rect 207952 53276 207958 53288
rect 207952 53248 215484 53276
rect 207952 53236 207958 53248
rect 186737 53211 186795 53217
rect 186737 53177 186749 53211
rect 186783 53208 186795 53211
rect 193453 53211 193511 53217
rect 193453 53208 193465 53211
rect 186783 53180 193465 53208
rect 186783 53177 186795 53180
rect 186737 53171 186795 53177
rect 193453 53177 193465 53180
rect 193499 53177 193511 53211
rect 193453 53171 193511 53177
rect 203021 53143 203079 53149
rect 203021 53109 203033 53143
rect 203067 53140 203079 53143
rect 205781 53143 205839 53149
rect 205781 53140 205793 53143
rect 203067 53112 205793 53140
rect 203067 53109 203079 53112
rect 203021 53103 203079 53109
rect 205781 53109 205793 53112
rect 205827 53109 205839 53143
rect 205781 53103 205839 53109
rect 183701 53075 183759 53081
rect 183701 53041 183713 53075
rect 183747 53072 183759 53075
rect 186737 53075 186795 53081
rect 186737 53072 186749 53075
rect 183747 53044 186749 53072
rect 183747 53041 183759 53044
rect 183701 53035 183759 53041
rect 186737 53041 186749 53044
rect 186783 53041 186795 53075
rect 186737 53035 186795 53041
rect 80198 52964 80204 53016
rect 80256 53004 80262 53016
rect 113962 53004 113968 53016
rect 80256 52976 113968 53004
rect 80256 52964 80262 52976
rect 113962 52964 113968 52976
rect 114020 53004 114026 53016
rect 139998 53004 140004 53016
rect 114020 52976 140004 53004
rect 114020 52964 114026 52976
rect 139998 52964 140004 52976
rect 140056 52964 140062 53016
rect 171830 52964 171836 53016
rect 171888 53004 171894 53016
rect 174133 53007 174191 53013
rect 174133 53004 174145 53007
rect 171888 52976 174145 53004
rect 171888 52964 171894 52976
rect 174133 52973 174145 52976
rect 174179 52973 174191 53007
rect 215456 53004 215484 53248
rect 215456 52976 222384 53004
rect 174133 52967 174191 52973
rect 222356 52936 222384 52976
rect 267878 52964 267884 53016
rect 267936 53004 267942 53016
rect 301642 53004 301648 53016
rect 267936 52976 301648 53004
rect 267936 52964 267942 52976
rect 301642 52964 301648 52976
rect 301700 53004 301706 53016
rect 301700 52976 316960 53004
rect 301700 52964 301706 52976
rect 233470 52936 233476 52948
rect 222356 52908 233476 52936
rect 233470 52896 233476 52908
rect 233528 52896 233534 52948
rect 316932 52936 316960 52976
rect 328506 52936 328512 52948
rect 316932 52908 328512 52936
rect 328506 52896 328512 52908
rect 328564 52896 328570 52948
rect 174133 52871 174191 52877
rect 174133 52837 174145 52871
rect 174179 52868 174191 52871
rect 183701 52871 183759 52877
rect 183701 52868 183713 52871
rect 174179 52840 183713 52868
rect 174179 52837 174191 52840
rect 174133 52831 174191 52837
rect 183701 52837 183713 52840
rect 183747 52837 183759 52871
rect 183701 52831 183759 52837
rect 91238 51536 91244 51588
rect 91296 51576 91302 51588
rect 134754 51576 134760 51588
rect 91296 51548 134760 51576
rect 91296 51536 91302 51548
rect 134754 51536 134760 51548
rect 134812 51536 134818 51588
rect 187286 51536 187292 51588
rect 187344 51576 187350 51588
rect 232090 51576 232096 51588
rect 187344 51548 232096 51576
rect 187344 51536 187350 51548
rect 232090 51536 232096 51548
rect 232148 51536 232154 51588
rect 279010 51536 279016 51588
rect 279068 51576 279074 51588
rect 323814 51576 323820 51588
rect 279068 51548 323820 51576
rect 279068 51536 279074 51548
rect 323814 51536 323820 51548
rect 323872 51536 323878 51588
rect 88294 51468 88300 51520
rect 88352 51508 88358 51520
rect 93630 51508 93636 51520
rect 88352 51480 93636 51508
rect 88352 51468 88358 51480
rect 93630 51468 93636 51480
rect 93688 51468 93694 51520
rect 184986 51468 184992 51520
rect 185044 51508 185050 51520
rect 228686 51508 228692 51520
rect 185044 51480 228692 51508
rect 185044 51468 185050 51480
rect 228686 51468 228692 51480
rect 228744 51468 228750 51520
rect 312774 51468 312780 51520
rect 312832 51508 312838 51520
rect 314246 51508 314252 51520
rect 312832 51480 314252 51508
rect 312832 51468 312838 51480
rect 314246 51468 314252 51480
rect 314304 51468 314310 51520
rect 314798 51468 314804 51520
rect 314856 51508 314862 51520
rect 316638 51508 316644 51520
rect 314856 51480 316644 51508
rect 314856 51468 314862 51480
rect 316638 51468 316644 51480
rect 316696 51468 316702 51520
rect 220958 51400 220964 51452
rect 221016 51440 221022 51452
rect 222614 51440 222620 51452
rect 221016 51412 222620 51440
rect 221016 51400 221022 51412
rect 222614 51400 222620 51412
rect 222672 51400 222678 51452
rect 125094 51264 125100 51316
rect 125152 51304 125158 51316
rect 125922 51304 125928 51316
rect 125152 51276 125928 51304
rect 125152 51264 125158 51276
rect 125922 51264 125928 51276
rect 125980 51264 125986 51316
rect 111938 51128 111944 51180
rect 111996 51168 112002 51180
rect 121230 51168 121236 51180
rect 111996 51140 121236 51168
rect 111996 51128 112002 51140
rect 121230 51128 121236 51140
rect 121288 51128 121294 51180
rect 205778 51128 205784 51180
rect 205836 51168 205842 51180
rect 215530 51168 215536 51180
rect 205836 51140 215536 51168
rect 205836 51128 205842 51140
rect 215530 51128 215536 51140
rect 215588 51128 215594 51180
rect 299618 51128 299624 51180
rect 299676 51168 299682 51180
rect 309554 51168 309560 51180
rect 299676 51140 309560 51168
rect 299676 51128 299682 51140
rect 309554 51128 309560 51140
rect 309612 51128 309618 51180
rect 106418 51060 106424 51112
rect 106476 51100 106482 51112
rect 119114 51100 119120 51112
rect 106476 51072 119120 51100
rect 106476 51060 106482 51072
rect 119114 51060 119120 51072
rect 119172 51060 119178 51112
rect 200258 51060 200264 51112
rect 200316 51100 200322 51112
rect 213230 51100 213236 51112
rect 200316 51072 213236 51100
rect 200316 51060 200322 51072
rect 213230 51060 213236 51072
rect 213288 51060 213294 51112
rect 294098 51060 294104 51112
rect 294156 51100 294162 51112
rect 307254 51100 307260 51112
rect 294156 51072 307260 51100
rect 294156 51060 294162 51072
rect 307254 51060 307260 51072
rect 307312 51060 307318 51112
rect 102278 50992 102284 51044
rect 102336 51032 102342 51044
rect 116538 51032 116544 51044
rect 102336 51004 116544 51032
rect 102336 50992 102342 51004
rect 116538 50992 116544 51004
rect 116596 50992 116602 51044
rect 196118 50992 196124 51044
rect 196176 51032 196182 51044
rect 210838 51032 210844 51044
rect 196176 51004 210844 51032
rect 196176 50992 196182 51004
rect 210838 50992 210844 51004
rect 210896 50992 210902 51044
rect 289958 50992 289964 51044
rect 290016 51032 290022 51044
rect 304862 51032 304868 51044
rect 290016 51004 304868 51032
rect 290016 50992 290022 51004
rect 304862 50992 304868 51004
rect 304920 50992 304926 51044
rect 96761 50967 96819 50973
rect 96761 50933 96773 50967
rect 96807 50964 96819 50967
rect 114146 50964 114152 50976
rect 96807 50936 114152 50964
rect 96807 50933 96819 50936
rect 96761 50927 96819 50933
rect 114146 50924 114152 50936
rect 114204 50924 114210 50976
rect 170450 50924 170456 50976
rect 170508 50964 170514 50976
rect 189678 50964 189684 50976
rect 170508 50936 189684 50964
rect 170508 50924 170514 50936
rect 189678 50924 189684 50936
rect 189736 50924 189742 50976
rect 190598 50924 190604 50976
rect 190656 50964 190662 50976
rect 208446 50964 208452 50976
rect 190656 50936 208452 50964
rect 190656 50924 190662 50936
rect 208446 50924 208452 50936
rect 208504 50924 208510 50976
rect 218934 50924 218940 50976
rect 218992 50964 218998 50976
rect 220222 50964 220228 50976
rect 218992 50936 220228 50964
rect 218992 50924 218998 50936
rect 220222 50924 220228 50936
rect 220280 50924 220286 50976
rect 284438 50924 284444 50976
rect 284496 50964 284502 50976
rect 302470 50964 302476 50976
rect 284496 50936 302476 50964
rect 284496 50924 284502 50936
rect 302470 50924 302476 50936
rect 302528 50924 302534 50976
rect 91238 50856 91244 50908
rect 91296 50896 91302 50908
rect 112030 50896 112036 50908
rect 91296 50868 112036 50896
rect 91296 50856 91302 50868
rect 112030 50856 112036 50868
rect 112088 50856 112094 50908
rect 116078 50856 116084 50908
rect 116136 50896 116142 50908
rect 123622 50896 123628 50908
rect 116136 50868 123628 50896
rect 116136 50856 116142 50868
rect 123622 50856 123628 50868
rect 123680 50856 123686 50908
rect 185078 50856 185084 50908
rect 185136 50896 185142 50908
rect 206146 50896 206152 50908
rect 185136 50868 206152 50896
rect 185136 50856 185142 50868
rect 206146 50856 206152 50868
rect 206204 50856 206210 50908
rect 280298 50856 280304 50908
rect 280356 50896 280362 50908
rect 300170 50896 300176 50908
rect 280356 50868 300176 50896
rect 280356 50856 280362 50868
rect 300170 50856 300176 50868
rect 300228 50856 300234 50908
rect 305138 50856 305144 50908
rect 305196 50896 305202 50908
rect 311946 50896 311952 50908
rect 305196 50868 311952 50896
rect 305196 50856 305202 50868
rect 311946 50856 311952 50868
rect 312004 50856 312010 50908
rect 127118 50380 127124 50432
rect 127176 50420 127182 50432
rect 128682 50420 128688 50432
rect 127176 50392 128688 50420
rect 127176 50380 127182 50392
rect 128682 50380 128688 50392
rect 128740 50380 128746 50432
rect 211298 50380 211304 50432
rect 211356 50420 211362 50432
rect 217922 50420 217928 50432
rect 211356 50392 217928 50420
rect 211356 50380 211362 50392
rect 217922 50380 217928 50392
rect 217980 50380 217986 50432
rect 78910 50312 78916 50364
rect 78968 50352 78974 50364
rect 108626 50352 108632 50364
rect 78968 50324 108632 50352
rect 78968 50312 78974 50324
rect 108626 50312 108632 50324
rect 108684 50352 108690 50364
rect 140642 50352 140648 50364
rect 108684 50324 140648 50352
rect 108684 50312 108690 50324
rect 140642 50312 140648 50324
rect 140700 50312 140706 50364
rect 173302 50312 173308 50364
rect 173360 50352 173366 50364
rect 202558 50352 202564 50364
rect 173360 50324 202564 50352
rect 173360 50312 173366 50324
rect 202558 50312 202564 50324
rect 202616 50352 202622 50364
rect 233562 50352 233568 50364
rect 202616 50324 233568 50352
rect 202616 50312 202622 50324
rect 233562 50312 233568 50324
rect 233620 50312 233626 50364
rect 267510 50312 267516 50364
rect 267568 50352 267574 50364
rect 296582 50352 296588 50364
rect 267568 50324 296588 50352
rect 267568 50312 267574 50324
rect 296582 50312 296588 50324
rect 296640 50352 296646 50364
rect 327678 50352 327684 50364
rect 296640 50324 327684 50352
rect 296640 50312 296646 50324
rect 327678 50312 327684 50324
rect 327736 50312 327742 50364
rect 80198 50244 80204 50296
rect 80256 50284 80262 50296
rect 103566 50284 103572 50296
rect 80256 50256 103572 50284
rect 80256 50244 80262 50256
rect 103566 50244 103572 50256
rect 103624 50284 103630 50296
rect 140366 50284 140372 50296
rect 103624 50256 140372 50284
rect 103624 50244 103630 50256
rect 140366 50244 140372 50256
rect 140424 50244 140430 50296
rect 173578 50244 173584 50296
rect 173636 50284 173642 50296
rect 197498 50284 197504 50296
rect 173636 50256 197504 50284
rect 173636 50244 173642 50256
rect 197498 50244 197504 50256
rect 197556 50284 197562 50296
rect 233470 50284 233476 50296
rect 197556 50256 233476 50284
rect 197556 50244 197562 50256
rect 233470 50244 233476 50256
rect 233528 50244 233534 50296
rect 266774 50244 266780 50296
rect 266832 50284 266838 50296
rect 291522 50284 291528 50296
rect 266832 50256 291528 50284
rect 266832 50244 266838 50256
rect 291522 50244 291528 50256
rect 291580 50284 291586 50296
rect 328414 50284 328420 50296
rect 291580 50256 328420 50284
rect 291580 50244 291586 50256
rect 328414 50244 328420 50256
rect 328472 50244 328478 50296
rect 88386 49496 88392 49548
rect 88444 49536 88450 49548
rect 102370 49536 102376 49548
rect 88444 49508 102376 49536
rect 88444 49496 88450 49508
rect 102370 49496 102376 49508
rect 102428 49496 102434 49548
rect 182134 49496 182140 49548
rect 182192 49536 182198 49548
rect 194370 49536 194376 49548
rect 182192 49508 194376 49536
rect 182192 49496 182198 49508
rect 194370 49496 194376 49508
rect 194428 49496 194434 49548
rect 276158 49496 276164 49548
rect 276216 49536 276222 49548
rect 288394 49536 288400 49548
rect 276216 49508 288400 49536
rect 276216 49496 276222 49508
rect 288394 49496 288400 49508
rect 288452 49496 288458 49548
rect 80198 48884 80204 48936
rect 80256 48924 80262 48936
rect 98598 48924 98604 48936
rect 80256 48896 98604 48924
rect 80256 48884 80262 48896
rect 98598 48884 98604 48896
rect 98656 48924 98662 48936
rect 140550 48924 140556 48936
rect 98656 48896 140556 48924
rect 98656 48884 98662 48896
rect 140550 48884 140556 48896
rect 140608 48884 140614 48936
rect 172934 48884 172940 48936
rect 172992 48924 172998 48936
rect 192530 48924 192536 48936
rect 172992 48896 192536 48924
rect 172992 48884 172998 48896
rect 192530 48884 192536 48896
rect 192588 48924 192594 48936
rect 233470 48924 233476 48936
rect 192588 48896 233476 48924
rect 192588 48884 192594 48896
rect 233470 48884 233476 48896
rect 233528 48884 233534 48936
rect 267878 48884 267884 48936
rect 267936 48924 267942 48936
rect 286554 48924 286560 48936
rect 267936 48896 286560 48924
rect 267936 48884 267942 48896
rect 286554 48884 286560 48896
rect 286612 48924 286618 48936
rect 328414 48924 328420 48936
rect 286612 48896 328420 48924
rect 286612 48884 286618 48896
rect 328414 48884 328420 48896
rect 328472 48884 328478 48936
rect 96758 48516 96764 48528
rect 96719 48488 96764 48516
rect 96758 48476 96764 48488
rect 96816 48476 96822 48528
rect 181858 48136 181864 48188
rect 181916 48176 181922 48188
rect 182226 48176 182232 48188
rect 181916 48148 182232 48176
rect 181916 48136 181922 48148
rect 182226 48136 182232 48148
rect 182284 48176 182290 48188
rect 196670 48176 196676 48188
rect 182284 48148 196676 48176
rect 182284 48136 182290 48148
rect 196670 48136 196676 48148
rect 196728 48136 196734 48188
rect 232090 48136 232096 48188
rect 232148 48176 232154 48188
rect 238622 48176 238628 48188
rect 232148 48148 238628 48176
rect 232148 48136 232154 48148
rect 238622 48136 238628 48148
rect 238680 48176 238686 48188
rect 241106 48176 241112 48188
rect 238680 48148 241112 48176
rect 238680 48136 238686 48148
rect 241106 48136 241112 48148
rect 241164 48136 241170 48188
rect 276066 48136 276072 48188
rect 276124 48176 276130 48188
rect 293086 48176 293092 48188
rect 276124 48148 293092 48176
rect 276124 48136 276130 48148
rect 293086 48136 293092 48148
rect 293144 48136 293150 48188
rect 116173 47839 116231 47845
rect 116173 47805 116185 47839
rect 116219 47836 116231 47839
rect 125741 47839 125799 47845
rect 125741 47836 125753 47839
rect 116219 47808 125753 47836
rect 116219 47805 116231 47808
rect 116173 47799 116231 47805
rect 125741 47805 125753 47808
rect 125787 47805 125799 47839
rect 125741 47799 125799 47805
rect 125833 47839 125891 47845
rect 125833 47805 125845 47839
rect 125879 47836 125891 47839
rect 135401 47839 135459 47845
rect 135401 47836 135413 47839
rect 125879 47808 135413 47836
rect 125879 47805 125891 47808
rect 125833 47799 125891 47805
rect 135401 47805 135413 47808
rect 135447 47805 135459 47839
rect 135401 47799 135459 47805
rect 80198 47660 80204 47712
rect 80256 47700 80262 47712
rect 109365 47703 109423 47709
rect 80256 47672 85856 47700
rect 80256 47660 80262 47672
rect 85828 47632 85856 47672
rect 109365 47669 109377 47703
rect 109411 47700 109423 47703
rect 116173 47703 116231 47709
rect 116173 47700 116185 47703
rect 109411 47672 116185 47700
rect 109411 47669 109423 47672
rect 109365 47663 109423 47669
rect 116173 47669 116185 47672
rect 116219 47669 116231 47703
rect 116173 47663 116231 47669
rect 135401 47703 135459 47709
rect 135401 47669 135413 47703
rect 135447 47700 135459 47703
rect 139998 47700 140004 47712
rect 135447 47672 140004 47700
rect 135447 47669 135459 47672
rect 135401 47663 135459 47669
rect 139998 47660 140004 47672
rect 140056 47660 140062 47712
rect 105041 47635 105099 47641
rect 85828 47604 93768 47632
rect 93740 47576 93768 47604
rect 105041 47601 105053 47635
rect 105087 47632 105099 47635
rect 109181 47635 109239 47641
rect 109181 47632 109193 47635
rect 105087 47604 109193 47632
rect 105087 47601 105099 47604
rect 105041 47595 105099 47601
rect 109181 47601 109193 47604
rect 109227 47601 109239 47635
rect 109181 47595 109239 47601
rect 125833 47635 125891 47641
rect 125833 47601 125845 47635
rect 125879 47601 125891 47635
rect 125833 47595 125891 47601
rect 93722 47524 93728 47576
rect 93780 47564 93786 47576
rect 95473 47567 95531 47573
rect 95473 47564 95485 47567
rect 93780 47536 95485 47564
rect 93780 47524 93786 47536
rect 95473 47533 95485 47536
rect 95519 47533 95531 47567
rect 95473 47527 95531 47533
rect 125741 47567 125799 47573
rect 125741 47533 125753 47567
rect 125787 47564 125799 47567
rect 125848 47564 125876 47595
rect 125787 47536 125876 47564
rect 125787 47533 125799 47536
rect 125741 47527 125799 47533
rect 142850 47524 142856 47576
rect 142908 47564 142914 47576
rect 159502 47564 159508 47576
rect 142908 47536 159508 47564
rect 142908 47524 142914 47536
rect 159502 47524 159508 47536
rect 159560 47524 159566 47576
rect 100254 47456 100260 47508
rect 100312 47496 100318 47508
rect 100438 47496 100444 47508
rect 100312 47468 100444 47496
rect 100312 47456 100318 47468
rect 100438 47456 100444 47468
rect 100496 47496 100502 47508
rect 125833 47499 125891 47505
rect 125833 47496 125845 47499
rect 100496 47468 125845 47496
rect 100496 47456 100502 47468
rect 125833 47465 125845 47468
rect 125879 47465 125891 47499
rect 125833 47459 125891 47465
rect 126017 47499 126075 47505
rect 126017 47465 126029 47499
rect 126063 47496 126075 47499
rect 156834 47496 156840 47508
rect 126063 47468 156840 47496
rect 126063 47465 126075 47468
rect 126017 47459 126075 47465
rect 156834 47456 156840 47468
rect 156892 47496 156898 47508
rect 167690 47496 167696 47508
rect 156892 47468 167696 47496
rect 156892 47456 156898 47468
rect 167690 47456 167696 47468
rect 167748 47456 167754 47508
rect 173302 47456 173308 47508
rect 173360 47496 173366 47508
rect 187562 47496 187568 47508
rect 173360 47468 187568 47496
rect 173360 47456 173366 47468
rect 187562 47456 187568 47468
rect 187620 47496 187626 47508
rect 233470 47496 233476 47508
rect 187620 47468 233476 47496
rect 187620 47456 187626 47468
rect 233470 47456 233476 47468
rect 233528 47456 233534 47508
rect 267878 47456 267884 47508
rect 267936 47496 267942 47508
rect 281586 47496 281592 47508
rect 267936 47468 281592 47496
rect 267936 47456 267942 47468
rect 281586 47456 281592 47468
rect 281644 47496 281650 47508
rect 327862 47496 327868 47508
rect 281644 47468 327868 47496
rect 281644 47456 281650 47468
rect 327862 47456 327868 47468
rect 327920 47456 327926 47508
rect 60694 47388 60700 47440
rect 60752 47428 60758 47440
rect 74218 47428 74224 47440
rect 60752 47400 74224 47428
rect 60752 47388 60758 47400
rect 74218 47388 74224 47400
rect 74276 47388 74282 47440
rect 95473 47431 95531 47437
rect 95473 47397 95485 47431
rect 95519 47428 95531 47431
rect 105041 47431 105099 47437
rect 105041 47428 105053 47431
rect 95519 47400 105053 47428
rect 95519 47397 95531 47400
rect 95473 47391 95531 47397
rect 105041 47397 105053 47400
rect 105087 47397 105099 47431
rect 105041 47391 105099 47397
rect 295478 47388 295484 47440
rect 295536 47428 295542 47440
rect 353622 47428 353628 47440
rect 295536 47400 353628 47428
rect 295536 47388 295542 47400
rect 353622 47388 353628 47400
rect 353680 47428 353686 47440
rect 419770 47428 419776 47440
rect 353680 47400 419776 47428
rect 353680 47388 353686 47400
rect 419770 47388 419776 47400
rect 419828 47388 419834 47440
rect 286002 47320 286008 47372
rect 286060 47360 286066 47372
rect 338350 47360 338356 47372
rect 286060 47332 338356 47360
rect 286060 47320 286066 47332
rect 338350 47320 338356 47332
rect 338408 47320 338414 47372
rect 74678 46776 74684 46828
rect 74736 46816 74742 46828
rect 88110 46816 88116 46828
rect 74736 46788 88116 46816
rect 74736 46776 74742 46788
rect 88110 46776 88116 46788
rect 88168 46776 88174 46828
rect 88018 46708 88024 46760
rect 88076 46748 88082 46760
rect 100254 46748 100260 46760
rect 88076 46720 100260 46748
rect 88076 46708 88082 46720
rect 100254 46708 100260 46720
rect 100312 46708 100318 46760
rect 275974 46708 275980 46760
rect 276032 46748 276038 46760
rect 295478 46748 295484 46760
rect 276032 46720 295484 46748
rect 276032 46708 276038 46720
rect 295478 46708 295484 46720
rect 295536 46708 295542 46760
rect 338350 46640 338356 46692
rect 338408 46680 338414 46692
rect 339638 46680 339644 46692
rect 338408 46652 339644 46680
rect 338408 46640 338414 46652
rect 339638 46640 339644 46652
rect 339696 46640 339702 46692
rect 73114 46164 73120 46216
rect 73172 46204 73178 46216
rect 88202 46204 88208 46216
rect 73172 46176 88208 46204
rect 73172 46164 73178 46176
rect 88202 46164 88208 46176
rect 88260 46204 88266 46216
rect 106602 46204 106608 46216
rect 88260 46176 106608 46204
rect 88260 46164 88266 46176
rect 106602 46164 106608 46176
rect 106660 46164 106666 46216
rect 74218 46096 74224 46148
rect 74276 46136 74282 46148
rect 88018 46136 88024 46148
rect 74276 46108 88024 46136
rect 74276 46096 74282 46108
rect 88018 46096 88024 46108
rect 88076 46096 88082 46148
rect 88110 46096 88116 46148
rect 88168 46136 88174 46148
rect 109454 46136 109460 46148
rect 88168 46108 109460 46136
rect 88168 46096 88174 46108
rect 109454 46096 109460 46108
rect 109512 46096 109518 46148
rect 317466 46136 317472 46148
rect 317427 46108 317472 46136
rect 317466 46096 317472 46108
rect 317524 46096 317530 46148
rect 167230 46028 167236 46080
rect 167288 46068 167294 46080
rect 169714 46068 169720 46080
rect 167288 46040 169720 46068
rect 167288 46028 167294 46040
rect 169714 46028 169720 46040
rect 169772 46028 169778 46080
rect 289961 46071 290019 46077
rect 289961 46037 289973 46071
rect 290007 46068 290019 46071
rect 298238 46068 298244 46080
rect 290007 46040 298244 46068
rect 290007 46037 290019 46040
rect 289961 46031 290019 46037
rect 298238 46028 298244 46040
rect 298296 46028 298302 46080
rect 350126 46028 350132 46080
rect 350184 46068 350190 46080
rect 361074 46068 361080 46080
rect 350184 46040 361080 46068
rect 350184 46028 350190 46040
rect 361074 46028 361080 46040
rect 361132 46028 361138 46080
rect 53702 45960 53708 46012
rect 53760 46000 53766 46012
rect 95470 46000 95476 46012
rect 53760 45972 95476 46000
rect 53760 45960 53766 45972
rect 95470 45960 95476 45972
rect 95528 45960 95534 46012
rect 144690 45960 144696 46012
rect 144748 46000 144754 46012
rect 369722 46000 369728 46012
rect 144748 45972 369728 46000
rect 144748 45960 144754 45972
rect 369722 45960 369728 45972
rect 369780 45960 369786 46012
rect 57198 45892 57204 45944
rect 57256 45932 57262 45944
rect 98046 45932 98052 45944
rect 57256 45904 98052 45932
rect 57256 45892 57262 45904
rect 98046 45892 98052 45904
rect 98104 45932 98110 45944
rect 153430 45932 153436 45944
rect 98104 45904 153436 45932
rect 98104 45892 98110 45904
rect 153430 45892 153436 45904
rect 153488 45892 153494 45944
rect 238622 45892 238628 45944
rect 238680 45932 238686 45944
rect 322526 45932 322532 45944
rect 238680 45904 322532 45932
rect 238680 45892 238686 45904
rect 322526 45892 322532 45904
rect 322584 45892 322590 45944
rect 332646 45892 332652 45944
rect 332704 45932 332710 45944
rect 369814 45932 369820 45944
rect 332704 45904 369820 45932
rect 332704 45892 332710 45904
rect 369814 45892 369820 45904
rect 369872 45892 369878 45944
rect 95470 45824 95476 45876
rect 95528 45864 95534 45876
rect 95746 45864 95752 45876
rect 95528 45836 95752 45864
rect 95528 45824 95534 45836
rect 95746 45824 95752 45836
rect 95804 45864 95810 45876
rect 150578 45864 150584 45876
rect 95804 45836 150584 45864
rect 95804 45824 95810 45836
rect 150578 45824 150584 45836
rect 150636 45864 150642 45876
rect 170174 45864 170180 45876
rect 150636 45836 170180 45864
rect 150636 45824 150642 45836
rect 170174 45824 170180 45836
rect 170232 45824 170238 45876
rect 250950 45824 250956 45876
rect 251008 45864 251014 45876
rect 275514 45864 275520 45876
rect 251008 45836 275520 45864
rect 251008 45824 251014 45836
rect 275514 45824 275520 45836
rect 275572 45864 275578 45876
rect 276158 45864 276164 45876
rect 275572 45836 276164 45864
rect 275572 45824 275578 45836
rect 276158 45824 276164 45836
rect 276216 45824 276222 45876
rect 298333 45867 298391 45873
rect 298333 45833 298345 45867
rect 298379 45864 298391 45867
rect 357118 45864 357124 45876
rect 298379 45836 357124 45864
rect 298379 45833 298391 45836
rect 298333 45827 298391 45833
rect 357118 45824 357124 45836
rect 357176 45824 357182 45876
rect 253986 45756 253992 45808
rect 254044 45796 254050 45808
rect 262542 45796 262548 45808
rect 254044 45768 262548 45796
rect 254044 45756 254050 45768
rect 262542 45756 262548 45768
rect 262600 45796 262606 45808
rect 263094 45796 263100 45808
rect 262600 45768 263100 45796
rect 262600 45756 262606 45768
rect 263094 45756 263100 45768
rect 263152 45756 263158 45808
rect 284346 45756 284352 45808
rect 284404 45796 284410 45808
rect 336142 45796 336148 45808
rect 284404 45768 336148 45796
rect 284404 45756 284410 45768
rect 336142 45756 336148 45768
rect 336200 45756 336206 45808
rect 347918 45756 347924 45808
rect 347976 45796 347982 45808
rect 359694 45796 359700 45808
rect 347976 45768 359700 45796
rect 347976 45756 347982 45768
rect 359694 45756 359700 45768
rect 359752 45756 359758 45808
rect 50206 45688 50212 45740
rect 50264 45728 50270 45740
rect 369170 45728 369176 45740
rect 50264 45700 369176 45728
rect 50264 45688 50270 45700
rect 369170 45688 369176 45700
rect 369228 45688 369234 45740
rect 298333 45663 298391 45669
rect 298333 45660 298345 45663
rect 298256 45632 298345 45660
rect 298256 45601 298284 45632
rect 298333 45629 298345 45632
rect 298379 45629 298391 45663
rect 298333 45623 298391 45629
rect 283153 45595 283211 45601
rect 283153 45561 283165 45595
rect 283199 45592 283211 45595
rect 289961 45595 290019 45601
rect 289961 45592 289973 45595
rect 283199 45564 289973 45592
rect 283199 45561 283211 45564
rect 283153 45555 283211 45561
rect 289961 45561 289973 45564
rect 290007 45561 290019 45595
rect 289961 45555 290019 45561
rect 298241 45595 298299 45601
rect 298241 45561 298253 45595
rect 298287 45561 298299 45595
rect 298241 45555 298299 45561
rect 278553 45527 278611 45533
rect 278553 45493 278565 45527
rect 278599 45524 278611 45527
rect 283061 45527 283119 45533
rect 283061 45524 283073 45527
rect 278599 45496 283073 45524
rect 278599 45493 278611 45496
rect 278553 45487 278611 45493
rect 283061 45493 283073 45496
rect 283107 45493 283119 45527
rect 283061 45487 283119 45493
rect 169530 45348 169536 45400
rect 169588 45388 169594 45400
rect 181950 45388 181956 45400
rect 169588 45360 181956 45388
rect 169588 45348 169594 45360
rect 181950 45348 181956 45360
rect 182008 45348 182014 45400
rect 182042 45348 182048 45400
rect 182100 45388 182106 45400
rect 201454 45388 201460 45400
rect 182100 45360 201460 45388
rect 182100 45348 182106 45360
rect 201454 45348 201460 45360
rect 201512 45348 201518 45400
rect 276066 45348 276072 45400
rect 276124 45388 276130 45400
rect 290694 45388 290700 45400
rect 276124 45360 290700 45388
rect 276124 45348 276130 45360
rect 290694 45348 290700 45360
rect 290752 45388 290758 45400
rect 324550 45388 324556 45400
rect 290752 45360 324556 45388
rect 290752 45348 290758 45360
rect 324550 45348 324556 45360
rect 324608 45388 324614 45400
rect 346630 45388 346636 45400
rect 324608 45360 346636 45388
rect 324608 45348 324614 45360
rect 346630 45348 346636 45360
rect 346688 45388 346694 45400
rect 347918 45388 347924 45400
rect 346688 45360 347924 45388
rect 346688 45348 346694 45360
rect 347918 45348 347924 45360
rect 347976 45348 347982 45400
rect 357118 45348 357124 45400
rect 357176 45388 357182 45400
rect 376990 45388 376996 45400
rect 357176 45360 376996 45388
rect 357176 45348 357182 45360
rect 376990 45348 376996 45360
rect 377048 45388 377054 45400
rect 422530 45388 422536 45400
rect 377048 45360 422536 45388
rect 377048 45348 377054 45360
rect 422530 45348 422536 45360
rect 422588 45348 422594 45400
rect 262818 45280 262824 45332
rect 262876 45320 262882 45332
rect 275882 45320 275888 45332
rect 262876 45292 275888 45320
rect 262876 45280 262882 45292
rect 275882 45280 275888 45292
rect 275940 45320 275946 45332
rect 278553 45323 278611 45329
rect 278553 45320 278565 45323
rect 275940 45292 278565 45320
rect 275940 45280 275946 45292
rect 278553 45289 278565 45292
rect 278599 45289 278611 45323
rect 278553 45283 278611 45289
rect 317101 44847 317159 44853
rect 317101 44813 317113 44847
rect 317147 44844 317159 44847
rect 317466 44844 317472 44856
rect 317147 44816 317472 44844
rect 317147 44813 317159 44816
rect 317101 44807 317159 44813
rect 317466 44804 317472 44816
rect 317524 44804 317530 44856
rect 169714 44736 169720 44788
rect 169772 44776 169778 44788
rect 182042 44776 182048 44788
rect 169772 44748 182048 44776
rect 169772 44736 169778 44748
rect 182042 44736 182048 44748
rect 182100 44736 182106 44788
rect 263094 44736 263100 44788
rect 263152 44776 263158 44788
rect 276066 44776 276072 44788
rect 263152 44748 276072 44776
rect 263152 44736 263158 44748
rect 276066 44736 276072 44748
rect 276124 44736 276130 44788
rect 12854 42560 12860 42612
rect 12912 42600 12918 42612
rect 16258 42600 16264 42612
rect 12912 42572 16264 42600
rect 12912 42560 12918 42572
rect 16258 42560 16264 42572
rect 16316 42560 16322 42612
rect 358406 40628 358412 40640
rect 358367 40600 358412 40628
rect 358406 40588 358412 40600
rect 358464 40588 358470 40640
rect 317098 37840 317104 37852
rect 317059 37812 317104 37840
rect 317098 37800 317104 37812
rect 317156 37800 317162 37852
rect 358406 37840 358412 37852
rect 358367 37812 358412 37840
rect 358406 37800 358412 37812
rect 358464 37800 358470 37852
rect 101358 37732 101364 37784
rect 101416 37772 101422 37784
rect 102278 37772 102284 37784
rect 101416 37744 102284 37772
rect 101416 37732 101422 37744
rect 102278 37732 102284 37744
rect 102336 37732 102342 37784
rect 210010 37732 210016 37784
rect 210068 37772 210074 37784
rect 211298 37772 211304 37784
rect 210068 37744 211304 37772
rect 210068 37732 210074 37744
rect 211298 37732 211304 37744
rect 211356 37732 211362 37784
rect 215070 37732 215076 37784
rect 215128 37772 215134 37784
rect 218934 37772 218940 37784
rect 215128 37744 218940 37772
rect 215128 37732 215134 37744
rect 218934 37732 218940 37744
rect 218992 37732 218998 37784
rect 220038 37732 220044 37784
rect 220096 37772 220102 37784
rect 220958 37772 220964 37784
rect 220096 37744 220964 37772
rect 220096 37732 220102 37744
rect 220958 37732 220964 37744
rect 221016 37732 221022 37784
rect 289038 37732 289044 37784
rect 289096 37772 289102 37784
rect 289958 37772 289964 37784
rect 289096 37744 289964 37772
rect 289096 37732 289102 37744
rect 289958 37732 289964 37744
rect 290016 37732 290022 37784
rect 304034 37732 304040 37784
rect 304092 37772 304098 37784
rect 305138 37772 305144 37784
rect 304092 37744 305144 37772
rect 304092 37732 304098 37744
rect 305138 37732 305144 37744
rect 305196 37732 305202 37784
rect 96390 37460 96396 37512
rect 96448 37500 96454 37512
rect 96758 37500 96764 37512
rect 96448 37472 96764 37500
rect 96448 37460 96454 37472
rect 96758 37460 96764 37472
rect 96816 37460 96822 37512
rect 195014 37392 195020 37444
rect 195072 37432 195078 37444
rect 196118 37432 196124 37444
rect 195072 37404 196124 37432
rect 195072 37392 195078 37404
rect 196118 37392 196124 37404
rect 196176 37392 196182 37444
rect 279102 37324 279108 37376
rect 279160 37364 279166 37376
rect 280298 37364 280304 37376
rect 279160 37336 280304 37364
rect 279160 37324 279166 37336
rect 280298 37324 280304 37336
rect 280356 37324 280362 37376
rect 121414 37120 121420 37172
rect 121472 37160 121478 37172
rect 125094 37160 125100 37172
rect 121472 37132 125100 37160
rect 121472 37120 121478 37132
rect 125094 37120 125100 37132
rect 125152 37120 125158 37172
rect 314062 37120 314068 37172
rect 314120 37160 314126 37172
rect 314798 37160 314804 37172
rect 314120 37132 314804 37160
rect 314120 37120 314126 37132
rect 314798 37120 314804 37132
rect 314856 37120 314862 37172
rect 309094 36712 309100 36764
rect 309152 36752 309158 36764
rect 312774 36752 312780 36764
rect 309152 36724 312780 36752
rect 309152 36712 309158 36724
rect 312774 36712 312780 36724
rect 312832 36712 312838 36764
rect 111386 36644 111392 36696
rect 111444 36684 111450 36696
rect 111938 36684 111944 36696
rect 111444 36656 111944 36684
rect 111444 36644 111450 36656
rect 111938 36644 111944 36656
rect 111996 36644 112002 36696
rect 126382 36576 126388 36628
rect 126440 36616 126446 36628
rect 127118 36616 127124 36628
rect 126440 36588 127124 36616
rect 126440 36576 126446 36588
rect 127118 36576 127124 36588
rect 127176 36576 127182 36628
rect 276158 33040 276164 33092
rect 276216 33080 276222 33092
rect 369630 33080 369636 33092
rect 276216 33052 369636 33080
rect 276216 33040 276222 33052
rect 369630 33040 369636 33052
rect 369688 33040 369694 33092
rect 182318 32972 182324 33024
rect 182376 33012 182382 33024
rect 369446 33012 369452 33024
rect 182376 32984 369452 33012
rect 182376 32972 182382 32984
rect 369446 32972 369452 32984
rect 369504 32972 369510 33024
rect 88478 32904 88484 32956
rect 88536 32944 88542 32956
rect 369170 32944 369176 32956
rect 88536 32916 369176 32944
rect 88536 32904 88542 32916
rect 369170 32904 369176 32916
rect 369228 32904 369234 32956
rect 12670 29436 12676 29488
rect 12728 29476 12734 29488
rect 16166 29476 16172 29488
rect 12728 29448 16172 29476
rect 12728 29436 12734 29448
rect 16166 29436 16172 29448
rect 16224 29436 16230 29488
rect 358222 28116 358228 28128
rect 358183 28088 358228 28116
rect 358222 28076 358228 28088
rect 358280 28076 358286 28128
rect 427498 28076 427504 28128
rect 427556 28116 427562 28128
rect 429798 28116 429804 28128
rect 427556 28088 429804 28116
rect 427556 28076 427562 28088
rect 429798 28076 429804 28088
rect 429856 28076 429862 28128
rect 358225 18531 358283 18537
rect 358225 18497 358237 18531
rect 358271 18528 358283 18531
rect 358314 18528 358320 18540
rect 358271 18500 358320 18528
rect 358271 18497 358283 18500
rect 358225 18491 358283 18497
rect 358314 18488 358320 18500
rect 358372 18488 358378 18540
rect 185170 17060 185176 17112
rect 185228 17100 185234 17112
rect 186366 17100 186372 17112
rect 185228 17072 186372 17100
rect 185228 17060 185234 17072
rect 186366 17060 186372 17072
rect 186424 17060 186430 17112
rect 191334 17060 191340 17112
rect 191392 17100 191398 17112
rect 192070 17100 192076 17112
rect 191392 17072 192076 17100
rect 191392 17060 191398 17072
rect 192070 17060 192076 17072
rect 192128 17060 192134 17112
rect 196118 17060 196124 17112
rect 196176 17100 196182 17112
rect 196302 17100 196308 17112
rect 196176 17072 196308 17100
rect 196176 17060 196182 17072
rect 196302 17060 196308 17072
rect 196360 17060 196366 17112
rect 92618 16788 92624 16840
rect 92676 16828 92682 16840
rect 105130 16828 105136 16840
rect 92676 16800 105136 16828
rect 92676 16788 92682 16800
rect 105130 16788 105136 16800
rect 105188 16788 105194 16840
rect 80750 16720 80756 16772
rect 80808 16760 80814 16772
rect 102370 16760 102376 16772
rect 80808 16732 102376 16760
rect 80808 16720 80814 16732
rect 102370 16720 102376 16732
rect 102428 16720 102434 16772
rect 285358 16720 285364 16772
rect 285416 16760 285422 16772
rect 299710 16760 299716 16772
rect 285416 16732 299716 16760
rect 285416 16720 285422 16732
rect 299710 16720 299716 16732
rect 299768 16720 299774 16772
rect 67870 16652 67876 16704
rect 67928 16692 67934 16704
rect 107062 16692 107068 16704
rect 67928 16664 107068 16692
rect 67928 16652 67934 16664
rect 107062 16652 107068 16664
rect 107120 16652 107126 16704
rect 170910 16652 170916 16704
rect 170968 16692 170974 16704
rect 201362 16692 201368 16704
rect 170968 16664 201368 16692
rect 170968 16652 170974 16664
rect 201362 16652 201368 16664
rect 201420 16652 201426 16704
rect 273950 16652 273956 16704
rect 274008 16692 274014 16704
rect 295386 16692 295392 16704
rect 274008 16664 295392 16692
rect 274008 16652 274014 16664
rect 295386 16652 295392 16664
rect 295444 16652 295450 16704
rect 54990 16584 54996 16636
rect 55048 16624 55054 16636
rect 112030 16624 112036 16636
rect 55048 16596 112036 16624
rect 55048 16584 55054 16596
rect 112030 16584 112036 16596
rect 112088 16584 112094 16636
rect 158030 16584 158036 16636
rect 158088 16624 158094 16636
rect 206330 16624 206336 16636
rect 158088 16596 206336 16624
rect 158088 16584 158094 16596
rect 206330 16584 206336 16596
rect 206388 16584 206394 16636
rect 261070 16584 261076 16636
rect 261128 16624 261134 16636
rect 300354 16624 300360 16636
rect 261128 16596 300360 16624
rect 261128 16584 261134 16596
rect 300354 16584 300360 16596
rect 300412 16584 300418 16636
rect 29230 16516 29236 16568
rect 29288 16556 29294 16568
rect 122058 16556 122064 16568
rect 29288 16528 122064 16556
rect 29288 16516 29294 16528
rect 122058 16516 122064 16528
rect 122116 16516 122122 16568
rect 145150 16516 145156 16568
rect 145208 16556 145214 16568
rect 211298 16556 211304 16568
rect 145208 16528 211304 16556
rect 145208 16516 145214 16528
rect 211298 16516 211304 16528
rect 211356 16516 211362 16568
rect 248190 16516 248196 16568
rect 248248 16556 248254 16568
rect 305322 16556 305328 16568
rect 248248 16528 305328 16556
rect 248248 16516 248254 16528
rect 305322 16516 305328 16528
rect 305380 16516 305386 16568
rect 42110 16448 42116 16500
rect 42168 16488 42174 16500
rect 116998 16488 117004 16500
rect 42168 16460 117004 16488
rect 42168 16448 42174 16460
rect 116998 16448 117004 16460
rect 117056 16448 117062 16500
rect 119390 16448 119396 16500
rect 119448 16488 119454 16500
rect 221326 16488 221332 16500
rect 119448 16460 221332 16488
rect 119448 16448 119454 16460
rect 221326 16448 221332 16460
rect 221384 16448 221390 16500
rect 235310 16448 235316 16500
rect 235368 16488 235374 16500
rect 310382 16488 310388 16500
rect 235368 16460 310388 16488
rect 235368 16448 235374 16460
rect 310382 16448 310388 16460
rect 310440 16448 310446 16500
rect 16350 16380 16356 16432
rect 16408 16420 16414 16432
rect 127210 16420 127216 16432
rect 16408 16392 127216 16420
rect 16408 16380 16414 16392
rect 127210 16380 127216 16392
rect 127268 16380 127274 16432
rect 132270 16380 132276 16432
rect 132328 16420 132334 16432
rect 216358 16420 216364 16432
rect 132328 16392 216364 16420
rect 132328 16380 132334 16392
rect 216358 16380 216364 16392
rect 216416 16380 216422 16432
rect 222430 16380 222436 16432
rect 222488 16420 222494 16432
rect 315350 16420 315356 16432
rect 222488 16392 315356 16420
rect 222488 16380 222494 16392
rect 315350 16380 315356 16392
rect 315408 16380 315414 16432
rect 13038 15564 13044 15616
rect 13096 15604 13102 15616
rect 16074 15604 16080 15616
rect 13096 15576 16080 15604
rect 13096 15564 13102 15576
rect 16074 15564 16080 15576
rect 16132 15564 16138 15616
rect 427314 15428 427320 15480
rect 427372 15468 427378 15480
rect 429430 15468 429436 15480
rect 427372 15440 429436 15468
rect 427372 15428 427378 15440
rect 429430 15428 429436 15440
rect 429488 15428 429494 15480
rect 351230 12912 351236 12964
rect 351288 12952 351294 12964
rect 358314 12952 358320 12964
rect 351288 12924 358320 12952
rect 351288 12912 351294 12924
rect 358314 12912 358320 12924
rect 358372 12912 358378 12964
rect 286830 12436 286836 12488
rect 286888 12476 286894 12488
rect 290050 12476 290056 12488
rect 286888 12448 290056 12476
rect 286888 12436 286894 12448
rect 290050 12436 290056 12448
rect 290108 12436 290114 12488
rect 280390 12368 280396 12420
rect 280448 12408 280454 12420
rect 312590 12408 312596 12420
rect 280448 12380 312596 12408
rect 280448 12368 280454 12380
rect 312590 12368 312596 12380
rect 312648 12368 312654 12420
rect 105130 12300 105136 12352
rect 105188 12340 105194 12352
rect 106510 12340 106516 12352
rect 105188 12312 106516 12340
rect 105188 12300 105194 12312
rect 106510 12300 106516 12312
rect 106568 12300 106574 12352
rect 183790 12300 183796 12352
rect 183848 12340 183854 12352
rect 196118 12340 196124 12352
rect 183848 12312 196124 12340
rect 183848 12300 183854 12312
rect 196118 12300 196124 12312
rect 196176 12300 196182 12352
rect 265854 12300 265860 12352
rect 265912 12340 265918 12352
rect 402750 12340 402756 12352
rect 265912 12312 402756 12340
rect 265912 12300 265918 12312
rect 402750 12300 402756 12312
rect 402808 12300 402814 12352
rect 93630 12232 93636 12284
rect 93688 12272 93694 12284
rect 96850 12272 96856 12284
rect 93688 12244 96856 12272
rect 93688 12232 93694 12244
rect 96850 12232 96856 12244
rect 96908 12232 96914 12284
rect 185170 12232 185176 12284
rect 185228 12272 185234 12284
rect 209550 12272 209556 12284
rect 185228 12244 209556 12272
rect 185228 12232 185234 12244
rect 209550 12232 209556 12244
rect 209608 12232 209614 12284
rect 228594 12232 228600 12284
rect 228652 12272 228658 12284
rect 415630 12272 415636 12284
rect 228652 12244 415636 12272
rect 228652 12232 228658 12244
rect 415630 12232 415636 12244
rect 415688 12232 415694 12284
rect 192070 12096 192076 12148
rect 192128 12136 192134 12148
rect 196670 12136 196676 12148
rect 192128 12108 196676 12136
rect 192128 12096 192134 12108
rect 196670 12096 196676 12108
rect 196728 12096 196734 12148
rect 385178 12096 385184 12148
rect 385236 12136 385242 12148
rect 389870 12136 389876 12148
rect 385236 12108 389876 12136
rect 385236 12096 385242 12108
rect 389870 12096 389876 12108
rect 389928 12096 389934 12148
rect 324550 9376 324556 9428
rect 324608 9416 324614 9428
rect 325470 9416 325476 9428
rect 324608 9388 325476 9416
rect 324608 9376 324614 9388
rect 325470 9376 325476 9388
rect 325528 9376 325534 9428
rect 428050 9376 428056 9428
rect 428108 9416 428114 9428
rect 428510 9416 428516 9428
rect 428108 9388 428516 9416
rect 428108 9376 428114 9388
rect 428510 9376 428516 9388
rect 428568 9376 428574 9428
<< via1 >>
rect 249024 395183 249076 395192
rect 249024 395149 249033 395183
rect 249033 395149 249067 395183
rect 249067 395149 249076 395183
rect 249024 395140 249076 395149
rect 88576 393780 88628 393832
rect 89588 393780 89640 393832
rect 106516 393780 106568 393832
rect 107252 393780 107304 393832
rect 124456 393780 124508 393832
rect 125008 393780 125060 393832
rect 212776 393780 212828 393832
rect 213512 393780 213564 393832
rect 355192 393780 355244 393832
rect 358596 393780 358648 393832
rect 70636 393644 70688 393696
rect 71832 393644 71884 393696
rect 337528 393372 337580 393424
rect 358504 393372 358556 393424
rect 304592 393304 304644 393356
rect 408368 393304 408420 393356
rect 299440 393236 299492 393288
rect 426032 393236 426084 393288
rect 106332 393168 106384 393220
rect 372948 393168 373000 393220
rect 91336 393100 91388 393152
rect 390612 393100 390664 393152
rect 18196 392760 18248 392812
rect 18748 392760 18800 392812
rect 314620 389700 314672 389752
rect 429436 389700 429488 389752
rect 70636 389292 70688 389344
rect 111300 389292 111352 389344
rect 54076 389224 54128 389276
rect 116268 389224 116320 389276
rect 124456 389224 124508 389276
rect 142672 389224 142724 389276
rect 194836 389224 194888 389276
rect 195848 389224 195900 389276
rect 283984 389224 284036 389276
rect 106516 389156 106568 389208
rect 205324 389156 205376 389208
rect 36136 389088 36188 389140
rect 121328 389088 121380 389140
rect 178092 389088 178144 389140
rect 288952 389088 289004 389140
rect 88576 389020 88628 389072
rect 210292 389020 210344 389072
rect 212776 389020 212828 389072
rect 279016 389020 279068 389072
rect 18196 388952 18248 389004
rect 126296 388952 126348 389004
rect 160428 388952 160480 389004
rect 294196 388952 294248 389004
rect 200356 388884 200408 388936
rect 96304 388544 96356 388596
rect 127860 388544 127912 388596
rect 185360 388544 185412 388596
rect 228600 388544 228652 388596
rect 13412 388476 13464 388528
rect 101272 388476 101324 388528
rect 190328 388476 190380 388528
rect 265860 388476 265912 388528
rect 13504 388408 13556 388460
rect 215352 388408 215404 388460
rect 220320 388408 220372 388460
rect 315632 388408 315684 388460
rect 13596 388340 13648 388392
rect 309008 388340 309060 388392
rect 249116 385552 249168 385604
rect 226484 382764 226536 382816
rect 227220 382764 227272 382816
rect 230900 382764 230952 382816
rect 315816 378616 315868 378668
rect 429436 378616 429488 378668
rect 248932 375896 248984 375948
rect 249024 375896 249076 375948
rect 226484 375148 226536 375200
rect 228784 375148 228836 375200
rect 248932 375148 248984 375200
rect 266596 373176 266648 373228
rect 266780 373176 266832 373228
rect 131816 371748 131868 371800
rect 134760 371748 134812 371800
rect 225840 371748 225892 371800
rect 229980 371748 230032 371800
rect 320324 371748 320376 371800
rect 362460 371748 362512 371800
rect 186280 368620 186332 368672
rect 191524 368620 191576 368672
rect 209004 368552 209056 368604
rect 210016 368552 210068 368604
rect 277544 368280 277596 368332
rect 280396 368280 280448 368332
rect 89864 367668 89916 367720
rect 92532 367668 92584 367720
rect 90048 367600 90100 367652
rect 91428 367600 91480 367652
rect 95016 367600 95068 367652
rect 96856 367600 96908 367652
rect 99984 367600 100036 367652
rect 100904 367600 100956 367652
rect 105044 367600 105096 367652
rect 106608 367600 106660 367652
rect 110012 367600 110064 367652
rect 112036 367600 112088 367652
rect 114980 367600 115032 367652
rect 116176 367600 116228 367652
rect 120040 367600 120092 367652
rect 121696 367600 121748 367652
rect 184072 367600 184124 367652
rect 185176 367600 185228 367652
rect 185268 367600 185320 367652
rect 186556 367600 186608 367652
rect 199068 367600 199120 367652
rect 200264 367600 200316 367652
rect 204036 367600 204088 367652
rect 205876 367600 205928 367652
rect 214064 367600 214116 367652
rect 215536 367600 215588 367652
rect 278372 367600 278424 367652
rect 279660 367600 279712 367652
rect 282972 367600 283024 367652
rect 283800 367600 283852 367652
rect 293368 367600 293420 367652
rect 294288 367600 294340 367652
rect 298244 367600 298296 367652
rect 299716 367600 299768 367652
rect 303304 367600 303356 367652
rect 305236 367600 305288 367652
rect 308364 367600 308416 367652
rect 309284 367600 309336 367652
rect 127860 366172 127912 366224
rect 429436 366172 429488 366224
rect 266596 363520 266648 363572
rect 266780 363520 266832 363572
rect 116176 363452 116228 363504
rect 117004 363452 117056 363504
rect 210016 363452 210068 363504
rect 211028 363452 211080 363504
rect 67692 359848 67744 359900
rect 75972 359848 76024 359900
rect 53708 359780 53760 359832
rect 76984 359780 77036 359832
rect 50212 359712 50264 359764
rect 76800 359712 76852 359764
rect 64196 359644 64248 359696
rect 75696 359644 75748 359696
rect 60700 359576 60752 359628
rect 75788 359576 75840 359628
rect 57204 359508 57256 359560
rect 76064 359508 76116 359560
rect 71188 359372 71240 359424
rect 75880 359372 75932 359424
rect 185176 358624 185228 358676
rect 186004 358624 186056 358676
rect 80204 357876 80256 357928
rect 127216 357876 127268 357928
rect 139636 357876 139688 357928
rect 174044 357876 174096 357928
rect 221056 357876 221108 357928
rect 233476 357876 233528 357928
rect 267332 357876 267384 357928
rect 314896 357876 314948 357928
rect 328420 357876 328472 357928
rect 75696 357536 75748 357588
rect 76432 357536 76484 357588
rect 75788 357468 75840 357520
rect 76156 357468 76208 357520
rect 74776 357400 74828 357452
rect 76892 357400 76944 357452
rect 80204 356516 80256 356568
rect 121788 356516 121840 356568
rect 139636 356516 139688 356568
rect 173492 356516 173544 356568
rect 215628 356516 215680 356568
rect 233476 356516 233528 356568
rect 266596 356516 266648 356568
rect 266780 356516 266832 356568
rect 267884 356516 267936 356568
rect 309376 356516 309428 356568
rect 328328 356516 328380 356568
rect 80204 355156 80256 355208
rect 117556 355156 117608 355208
rect 139636 355156 139688 355208
rect 174044 355156 174096 355208
rect 211396 355156 211448 355208
rect 233476 355156 233528 355208
rect 266780 355156 266832 355208
rect 266872 355156 266924 355208
rect 267884 355156 267936 355208
rect 305328 355156 305380 355208
rect 328420 355156 328472 355208
rect 79284 355088 79336 355140
rect 112128 355088 112180 355140
rect 139728 355088 139780 355140
rect 173768 355088 173820 355140
rect 205968 355088 206020 355140
rect 233568 355088 233620 355140
rect 267424 355088 267476 355140
rect 299808 355088 299860 355140
rect 328512 355088 328564 355140
rect 100904 355020 100956 355072
rect 102376 355020 102428 355072
rect 125744 355020 125796 355072
rect 127216 355020 127268 355072
rect 194744 355020 194796 355072
rect 196308 355020 196360 355072
rect 279660 355020 279712 355072
rect 280396 355020 280448 355072
rect 283800 355020 283852 355072
rect 285364 355020 285416 355072
rect 288584 355020 288636 355072
rect 290332 355020 290384 355072
rect 309284 355020 309336 355072
rect 310388 355020 310440 355072
rect 313424 355020 313476 355072
rect 315356 355020 315408 355072
rect 76064 354000 76116 354052
rect 189224 354000 189276 354052
rect 191340 354000 191392 354052
rect 200264 354000 200316 354052
rect 201368 354000 201420 354052
rect 76248 353864 76300 353916
rect 219584 353864 219636 353916
rect 221332 353864 221384 353916
rect 78916 353796 78968 353848
rect 106516 353796 106568 353848
rect 139636 353796 139688 353848
rect 174044 353796 174096 353848
rect 200356 353796 200408 353848
rect 233476 353796 233528 353848
rect 267884 353796 267936 353848
rect 294196 353796 294248 353848
rect 328052 353796 328104 353848
rect 80204 352368 80256 352420
rect 102652 352368 102704 352420
rect 139636 352368 139688 352420
rect 174044 352368 174096 352420
rect 196216 352368 196268 352420
rect 233476 352368 233528 352420
rect 267884 352368 267936 352420
rect 290056 352368 290108 352420
rect 328512 352368 328564 352420
rect 97316 352003 97368 352012
rect 97316 351969 97325 352003
rect 97325 351969 97359 352003
rect 97359 351969 97368 352003
rect 97316 351960 97368 351969
rect 186280 351867 186332 351876
rect 186280 351833 186289 351867
rect 186289 351833 186323 351867
rect 186323 351833 186332 351867
rect 186280 351824 186332 351833
rect 284996 351595 285048 351604
rect 284996 351561 285005 351595
rect 285005 351561 285039 351595
rect 285039 351561 285048 351595
rect 284996 351552 285048 351561
rect 226300 351280 226352 351332
rect 231636 351280 231688 351332
rect 131816 351076 131868 351128
rect 137428 351076 137480 351128
rect 320600 351076 320652 351128
rect 327224 351076 327276 351128
rect 79100 351008 79152 351060
rect 89864 351008 89916 351060
rect 139636 351008 139688 351060
rect 173768 351008 173820 351060
rect 185268 351008 185320 351060
rect 233568 351008 233620 351060
rect 267516 351008 267568 351060
rect 277544 351008 277596 351060
rect 327868 351008 327920 351060
rect 174044 350940 174096 350992
rect 233476 350940 233528 350992
rect 80204 350328 80256 350380
rect 139728 350328 139780 350380
rect 267700 350328 267752 350380
rect 327500 350328 327552 350380
rect 131816 349716 131868 349768
rect 137520 349716 137572 349768
rect 226392 349716 226444 349768
rect 231176 349716 231228 349768
rect 321612 349716 321664 349768
rect 327132 349716 327184 349768
rect 80204 349648 80256 349700
rect 87196 349648 87248 349700
rect 137428 349648 137480 349700
rect 139636 349648 139688 349700
rect 231636 349648 231688 349700
rect 233476 349648 233528 349700
rect 267884 349648 267936 349700
rect 274784 349648 274836 349700
rect 173032 349036 173084 349088
rect 180852 349036 180904 349088
rect 321612 348424 321664 348476
rect 327040 348424 327092 348476
rect 131908 348356 131960 348408
rect 137428 348356 137480 348408
rect 226392 348356 226444 348408
rect 233292 348356 233344 348408
rect 131816 348288 131868 348340
rect 137612 348288 137664 348340
rect 226484 348288 226536 348340
rect 233384 348288 233436 348340
rect 320692 348288 320744 348340
rect 327224 348288 327276 348340
rect 80204 348220 80256 348272
rect 87472 348220 87524 348272
rect 137520 348220 137572 348272
rect 139636 348220 139688 348272
rect 231176 348220 231228 348272
rect 233476 348220 233528 348272
rect 267884 348220 267936 348272
rect 274968 348220 275020 348272
rect 172940 347948 172992 348000
rect 180944 347948 180996 348000
rect 132184 346928 132236 346980
rect 139820 346928 139872 346980
rect 226392 346928 226444 346980
rect 228416 346928 228468 346980
rect 321060 346928 321112 346980
rect 323176 346928 323228 346980
rect 80204 346860 80256 346912
rect 87288 346860 87340 346912
rect 137428 346860 137480 346912
rect 139636 346860 139688 346912
rect 174044 346860 174096 346912
rect 182324 346860 182376 346912
rect 267884 346860 267936 346912
rect 274876 346860 274928 346912
rect 79284 346792 79336 346844
rect 87380 346792 87432 346844
rect 137612 346792 137664 346844
rect 139728 346792 139780 346844
rect 173768 346792 173820 346844
rect 182140 346792 182192 346844
rect 267424 346792 267476 346844
rect 275060 346792 275112 346844
rect 321612 345704 321664 345756
rect 326948 345704 327000 345756
rect 131816 345636 131868 345688
rect 134116 345636 134168 345688
rect 172848 345636 172900 345688
rect 181588 345636 181640 345688
rect 226300 345636 226352 345688
rect 227956 345636 228008 345688
rect 79652 345568 79704 345620
rect 87196 345568 87248 345620
rect 131908 345568 131960 345620
rect 139636 345568 139688 345620
rect 172940 345568 172992 345620
rect 182324 345568 182376 345620
rect 226392 345568 226444 345620
rect 234580 345568 234632 345620
rect 270736 345568 270788 345620
rect 274876 345568 274928 345620
rect 320508 345568 320560 345620
rect 323268 345568 323320 345620
rect 228416 345500 228468 345552
rect 233476 345500 233528 345552
rect 267884 345500 267936 345552
rect 275152 345500 275204 345552
rect 323176 345500 323228 345552
rect 328052 345500 328104 345552
rect 80204 344752 80256 344804
rect 87104 344752 87156 344804
rect 172756 344752 172808 344804
rect 180944 344752 180996 344804
rect 85816 344616 85868 344668
rect 87380 344616 87432 344668
rect 320968 344480 321020 344532
rect 323268 344480 323320 344532
rect 131816 344208 131868 344260
rect 139820 344208 139872 344260
rect 226484 344208 226536 344260
rect 234488 344208 234540 344260
rect 321612 344208 321664 344260
rect 327408 344208 327460 344260
rect 132368 344140 132420 344192
rect 139728 344140 139780 344192
rect 173124 344140 173176 344192
rect 182324 344140 182376 344192
rect 226392 344140 226444 344192
rect 234396 344140 234448 344192
rect 76064 344072 76116 344124
rect 76156 344072 76208 344124
rect 227956 344072 228008 344124
rect 233476 344072 233528 344124
rect 266688 344072 266740 344124
rect 274968 344072 275020 344124
rect 323176 344072 323228 344124
rect 328512 344072 328564 344124
rect 76156 343732 76208 343784
rect 321612 342848 321664 342900
rect 327224 342848 327276 342900
rect 131816 342780 131868 342832
rect 137520 342780 137572 342832
rect 173952 342780 174004 342832
rect 181404 342780 181456 342832
rect 226392 342780 226444 342832
rect 230532 342780 230584 342832
rect 80204 342712 80256 342764
rect 88116 342712 88168 342764
rect 134116 342712 134168 342764
rect 139636 342712 139688 342764
rect 172756 342712 172808 342764
rect 180944 342712 180996 342764
rect 267608 342712 267660 342764
rect 274876 342712 274928 342764
rect 323268 342712 323320 342764
rect 328052 342712 328104 342764
rect 267884 342644 267936 342696
rect 270736 342644 270788 342696
rect 80204 342100 80256 342152
rect 85816 342100 85868 342152
rect 131908 341488 131960 341540
rect 135404 341488 135456 341540
rect 173768 341488 173820 341540
rect 182324 341488 182376 341540
rect 226484 341488 226536 341540
rect 232004 341488 232056 341540
rect 321060 341488 321112 341540
rect 327132 341488 327184 341540
rect 131816 341420 131868 341472
rect 135312 341420 135364 341472
rect 174044 341420 174096 341472
rect 181404 341420 181456 341472
rect 226392 341420 226444 341472
rect 231820 341420 231872 341472
rect 321612 341420 321664 341472
rect 327040 341420 327092 341472
rect 80204 341352 80256 341404
rect 88484 341352 88536 341404
rect 267884 341352 267936 341404
rect 275060 341352 275112 341404
rect 131816 340060 131868 340112
rect 139544 340060 139596 340112
rect 173860 340060 173912 340112
rect 181404 340060 181456 340112
rect 226392 340060 226444 340112
rect 233568 340060 233620 340112
rect 272024 340060 272076 340112
rect 274876 340060 274928 340112
rect 320600 340060 320652 340112
rect 327868 340060 327920 340112
rect 374144 340060 374196 340112
rect 429436 340060 429488 340112
rect 80204 339992 80256 340044
rect 87288 339992 87340 340044
rect 137520 339992 137572 340044
rect 139636 339992 139688 340044
rect 230532 339992 230584 340044
rect 233476 339992 233528 340044
rect 267884 339992 267936 340044
rect 275152 339992 275204 340044
rect 267148 339312 267200 339364
rect 320416 338768 320468 338820
rect 326580 338768 326632 338820
rect 131816 338700 131868 338752
rect 136140 338700 136192 338752
rect 226484 338700 226536 338752
rect 231912 338700 231964 338752
rect 85080 338632 85132 338684
rect 87472 338632 87524 338684
rect 131908 338632 131960 338684
rect 139636 338632 139688 338684
rect 173492 338632 173544 338684
rect 181588 338632 181640 338684
rect 226392 338632 226444 338684
rect 234120 338632 234172 338684
rect 267792 338632 267844 338684
rect 274876 338632 274928 338684
rect 320508 338632 320560 338684
rect 327224 338632 327276 338684
rect 80204 338564 80256 338616
rect 87564 338564 87616 338616
rect 135404 338564 135456 338616
rect 139728 338564 139780 338616
rect 232004 338564 232056 338616
rect 233476 338564 233528 338616
rect 267516 338564 267568 338616
rect 274968 338564 275020 338616
rect 80112 338496 80164 338548
rect 87196 338496 87248 338548
rect 135312 338496 135364 338548
rect 139820 338496 139872 338548
rect 231820 338496 231872 338548
rect 233660 338496 233712 338548
rect 267884 338496 267936 338548
rect 275244 338496 275296 338548
rect 226392 337612 226444 337664
rect 231544 337612 231596 337664
rect 85172 337272 85224 337324
rect 87196 337272 87248 337324
rect 131816 337272 131868 337324
rect 136232 337272 136284 337324
rect 173676 337272 173728 337324
rect 181772 337272 181824 337324
rect 270828 337272 270880 337324
rect 274876 337272 274928 337324
rect 320416 337272 320468 337324
rect 326764 337272 326816 337324
rect 79836 337204 79888 337256
rect 87380 337204 87432 337256
rect 267332 337204 267384 337256
rect 272024 337204 272076 337256
rect 320416 336048 320468 336100
rect 327316 336048 327368 336100
rect 131908 335980 131960 336032
rect 137612 335980 137664 336032
rect 172848 335980 172900 336032
rect 181588 335980 181640 336032
rect 270736 335980 270788 336032
rect 274968 335980 275020 336032
rect 85816 335912 85868 335964
rect 87196 335912 87248 335964
rect 131816 335912 131868 335964
rect 139820 335912 139872 335964
rect 172940 335912 172992 335964
rect 181772 335912 181824 335964
rect 226392 335912 226444 335964
rect 230716 335912 230768 335964
rect 266780 335912 266832 335964
rect 274876 335912 274928 335964
rect 80204 335844 80256 335896
rect 87288 335844 87340 335896
rect 231912 335844 231964 335896
rect 233476 335844 233528 335896
rect 267884 335844 267936 335896
rect 275060 335844 275112 335896
rect 75972 334756 76024 334808
rect 75880 334688 75932 334740
rect 76064 334688 76116 334740
rect 75972 334527 76024 334536
rect 75972 334493 75981 334527
rect 75981 334493 76015 334527
rect 76015 334493 76024 334527
rect 75972 334484 76024 334493
rect 76064 334484 76116 334536
rect 108264 334416 108316 334468
rect 131632 334416 131684 334468
rect 136140 334416 136192 334468
rect 139636 334416 139688 334468
rect 202472 334416 202524 334468
rect 225380 334416 225432 334468
rect 267332 334416 267384 334468
rect 270828 334416 270880 334468
rect 306248 334416 306300 334468
rect 319128 334416 319180 334468
rect 319680 334416 319732 334468
rect 75880 334348 75932 334400
rect 104860 334348 104912 334400
rect 131724 334348 131776 334400
rect 174044 334348 174096 334400
rect 180300 334348 180352 334400
rect 212316 334348 212368 334400
rect 225196 334348 225248 334400
rect 75972 334280 76024 334332
rect 76984 334280 77036 334332
rect 98236 334280 98288 334332
rect 111392 334280 111444 334332
rect 131540 334280 131592 334332
rect 114796 334212 114848 334264
rect 131448 334212 131500 334264
rect 136232 334212 136284 334264
rect 139636 334212 139688 334264
rect 118200 334144 118252 334196
rect 131356 334144 131408 334196
rect 131724 334144 131776 334196
rect 136876 334144 136928 334196
rect 131540 334076 131592 334128
rect 137060 334076 137112 334128
rect 231544 334076 231596 334128
rect 234304 334076 234356 334128
rect 80204 334008 80256 334060
rect 85172 334008 85224 334060
rect 116084 334008 116136 334060
rect 127860 334008 127912 334060
rect 131632 334008 131684 334060
rect 137336 334008 137388 334060
rect 103664 333940 103716 333992
rect 124548 333940 124600 333992
rect 131448 333940 131500 333992
rect 137520 333940 137572 333992
rect 211304 333940 211356 333992
rect 221884 333940 221936 333992
rect 305144 333940 305196 333992
rect 316184 333940 316236 333992
rect 80112 333872 80164 333924
rect 85080 333872 85132 333924
rect 91244 333872 91296 333924
rect 121236 333872 121288 333924
rect 131356 333872 131408 333924
rect 137704 333872 137756 333924
rect 197504 333872 197556 333924
rect 218572 333872 218624 333924
rect 292724 333872 292776 333924
rect 312872 333872 312924 333924
rect 98236 333804 98288 333856
rect 137796 333804 137848 333856
rect 185084 333804 185136 333856
rect 215628 333804 215680 333856
rect 280304 333804 280356 333856
rect 309560 333804 309612 333856
rect 91888 333736 91940 333788
rect 134852 333736 134904 333788
rect 185912 333736 185964 333788
rect 228692 333736 228744 333788
rect 279568 333736 279620 333788
rect 323820 333736 323872 333788
rect 225196 333532 225248 333584
rect 230992 333532 231044 333584
rect 231820 333532 231872 333584
rect 225380 333124 225432 333176
rect 231360 333124 231412 333176
rect 319680 333124 319732 333176
rect 325384 333124 325436 333176
rect 80204 333056 80256 333108
rect 87564 333056 87616 333108
rect 137612 333056 137664 333108
rect 139636 333056 139688 333108
rect 230716 333056 230768 333108
rect 233936 333056 233988 333108
rect 267148 333056 267200 333108
rect 270736 333056 270788 333108
rect 198792 332920 198844 332972
rect 228784 332920 228836 332972
rect 231452 332920 231504 332972
rect 319864 331764 319916 331816
rect 325200 331764 325252 331816
rect 76892 331696 76944 331748
rect 118200 331696 118252 331748
rect 226576 331696 226628 331748
rect 233476 331696 233528 331748
rect 114796 331628 114848 331680
rect 111392 331560 111444 331612
rect 319128 331696 319180 331748
rect 320508 331696 320560 331748
rect 328512 331696 328564 331748
rect 299532 331492 299584 331544
rect 80204 330744 80256 330796
rect 85816 330744 85868 330796
rect 225288 330608 225340 330660
rect 231728 330608 231780 330660
rect 319680 330472 319732 330524
rect 325752 330472 325804 330524
rect 319128 330404 319180 330456
rect 325292 330404 325344 330456
rect 75512 330175 75564 330184
rect 75512 330141 75521 330175
rect 75521 330141 75555 330175
rect 75555 330141 75564 330175
rect 75512 330132 75564 330141
rect 75420 330107 75472 330116
rect 75420 330073 75429 330107
rect 75429 330073 75463 330107
rect 75463 330073 75472 330107
rect 75420 330064 75472 330073
rect 82320 328976 82372 329028
rect 128504 329180 128556 329232
rect 140556 329180 140608 329232
rect 222528 329180 222580 329232
rect 233476 329180 233528 329232
rect 267884 329112 267936 329164
rect 319588 329180 319640 329232
rect 173400 329044 173452 329096
rect 137704 328976 137756 329028
rect 137888 328976 137940 329028
rect 161716 328976 161768 329028
rect 231360 328976 231412 329028
rect 231728 328976 231780 329028
rect 253716 328976 253768 329028
rect 299532 328976 299584 329028
rect 316552 329044 316604 329096
rect 209280 328908 209332 328960
rect 227220 328908 227272 328960
rect 231452 328908 231504 328960
rect 285916 328908 285968 328960
rect 303120 328908 303172 328960
rect 319036 328908 319088 328960
rect 324740 328908 324792 328960
rect 285916 328228 285968 328280
rect 325660 328228 325712 328280
rect 345256 327616 345308 327668
rect 346084 327616 346136 327668
rect 76064 327548 76116 327600
rect 100996 327548 101048 327600
rect 102284 327548 102336 327600
rect 137336 327548 137388 327600
rect 137520 327548 137572 327600
rect 137704 327548 137756 327600
rect 160980 327548 161032 327600
rect 209280 327548 209332 327600
rect 231452 327548 231504 327600
rect 254360 327548 254412 327600
rect 303120 327548 303172 327600
rect 337160 327548 337212 327600
rect 352800 327548 352852 327600
rect 158404 327480 158456 327532
rect 239548 327480 239600 327532
rect 248840 327480 248892 327532
rect 249576 327480 249628 327532
rect 250496 327480 250548 327532
rect 288676 327480 288728 327532
rect 341300 327480 341352 327532
rect 357584 327480 357636 327532
rect 137796 327412 137848 327464
rect 155920 327412 155972 327464
rect 192076 327412 192128 327464
rect 232004 327412 232056 327464
rect 249116 327412 249168 327464
rect 281776 327412 281828 327464
rect 341024 327412 341076 327464
rect 356020 327412 356072 327464
rect 58308 327344 58360 327396
rect 59228 327344 59280 327396
rect 62356 327344 62408 327396
rect 63368 327344 63420 327396
rect 65208 327344 65260 327396
rect 68520 327344 68572 327396
rect 154816 327344 154868 327396
rect 187936 327344 187988 327396
rect 189224 327344 189276 327396
rect 241756 327344 241808 327396
rect 242768 327344 242820 327396
rect 248932 327344 248984 327396
rect 256292 327344 256344 327396
rect 339644 327344 339696 327396
rect 353628 327344 353680 327396
rect 150860 327276 150912 327328
rect 165212 327276 165264 327328
rect 342404 327276 342456 327328
rect 355560 327276 355612 327328
rect 149388 327208 149440 327260
rect 163280 327208 163332 327260
rect 250496 327208 250548 327260
rect 258408 327208 258460 327260
rect 345624 327208 345676 327260
rect 359700 327208 359752 327260
rect 152240 327140 152292 327192
rect 166132 327140 166184 327192
rect 238628 327140 238680 327192
rect 244424 327140 244476 327192
rect 247184 327140 247236 327192
rect 258960 327140 259012 327192
rect 344796 327140 344848 327192
rect 358320 327140 358372 327192
rect 154080 327072 154132 327124
rect 168064 327072 168116 327124
rect 194836 327072 194888 327124
rect 232096 327072 232148 327124
rect 244240 327072 244292 327124
rect 257304 327072 257356 327124
rect 288676 327072 288728 327124
rect 325108 327072 325160 327124
rect 341208 327072 341260 327124
rect 358412 327072 358464 327124
rect 150768 327004 150820 327056
rect 164568 327004 164620 327056
rect 192076 327004 192128 327056
rect 233476 327004 233528 327056
rect 249576 327004 249628 327056
rect 250036 327004 250088 327056
rect 264112 327004 264164 327056
rect 281776 327004 281828 327056
rect 282880 327004 282932 327056
rect 325568 327004 325620 327056
rect 339920 327004 339972 327056
rect 356756 327004 356808 327056
rect 137612 326936 137664 326988
rect 154816 326936 154868 326988
rect 156288 326936 156340 326988
rect 169996 326936 170048 326988
rect 189224 326936 189276 326988
rect 230716 326936 230768 326988
rect 232004 326936 232056 326988
rect 248288 326936 248340 326988
rect 365220 326936 365272 326988
rect 102284 326868 102336 326920
rect 136968 326868 137020 326920
rect 154264 326868 154316 326920
rect 326580 326868 326632 326920
rect 335688 326868 335740 326920
rect 336792 326868 336844 326920
rect 338540 326868 338592 326920
rect 355192 326868 355244 326920
rect 154908 326800 154960 326852
rect 169076 326800 169128 326852
rect 238996 326800 239048 326852
rect 239916 326800 239968 326852
rect 245896 326800 245948 326852
rect 260156 326800 260208 326852
rect 334216 326800 334268 326852
rect 335228 326800 335280 326852
rect 339368 326800 339420 326852
rect 354364 326800 354416 326852
rect 153528 326732 153580 326784
rect 167328 326732 167380 326784
rect 247276 326732 247328 326784
rect 261168 326732 261220 326784
rect 343232 326732 343284 326784
rect 355652 326732 355704 326784
rect 144604 326664 144656 326716
rect 156196 326664 156248 326716
rect 248656 326664 248708 326716
rect 263100 326664 263152 326716
rect 340840 326664 340892 326716
rect 352800 326664 352852 326716
rect 65116 326596 65168 326648
rect 69624 326596 69676 326648
rect 147456 326596 147508 326648
rect 159048 326596 159100 326648
rect 241480 326596 241532 326648
rect 252888 326596 252940 326648
rect 259696 326596 259748 326648
rect 262088 326596 262140 326648
rect 341576 326596 341628 326648
rect 354180 326596 354232 326648
rect 148468 326528 148520 326580
rect 160244 326528 160296 326580
rect 246356 326528 246408 326580
rect 258316 326528 258368 326580
rect 332928 326528 332980 326580
rect 333664 326528 333716 326580
rect 343968 326528 344020 326580
rect 356940 326528 356992 326580
rect 136968 326460 137020 326512
rect 150400 326460 150452 326512
rect 158956 326460 159008 326512
rect 242492 326460 242544 326512
rect 254084 326460 254136 326512
rect 337068 326460 337120 326512
rect 351972 326460 352024 326512
rect 152148 326392 152200 326444
rect 163004 326392 163056 326444
rect 244332 326392 244384 326444
rect 253532 326392 253584 326444
rect 74040 326324 74092 326376
rect 76064 326324 76116 326376
rect 145524 326324 145576 326376
rect 152332 326324 152384 326376
rect 156840 326324 156892 326376
rect 244516 326324 244568 326376
rect 75788 326256 75840 326308
rect 76984 326256 77036 326308
rect 145340 326256 145392 326308
rect 145892 326256 145944 326308
rect 147916 326256 147968 326308
rect 148744 326256 148796 326308
rect 151320 326256 151372 326308
rect 154816 326256 154868 326308
rect 155644 326256 155696 326308
rect 162268 326256 162320 326308
rect 194836 326256 194888 326308
rect 243228 326256 243280 326308
rect 244240 326256 244292 326308
rect 245344 326256 245396 326308
rect 248748 326256 248800 326308
rect 254544 326256 254596 326308
rect 259236 326256 259288 326308
rect 70636 325236 70688 325288
rect 71372 325236 71424 325288
rect 348016 325168 348068 325220
rect 348476 325168 348528 325220
rect 54076 324828 54128 324880
rect 54812 324828 54864 324880
rect 325108 324828 325160 324880
rect 343968 324828 344020 324880
rect 347188 324828 347240 324880
rect 279108 324760 279160 324812
rect 280304 324760 280356 324812
rect 291528 324760 291580 324812
rect 292724 324760 292776 324812
rect 210016 324148 210068 324200
rect 211304 324148 211356 324200
rect 344796 324080 344848 324132
rect 348108 324080 348160 324132
rect 304040 324012 304092 324064
rect 305144 324012 305196 324064
rect 325752 323468 325804 323520
rect 344796 323468 344848 323520
rect 343876 322788 343928 322840
rect 345164 322788 345216 322840
rect 348016 322788 348068 322840
rect 324556 322720 324608 322772
rect 325384 322720 325436 322772
rect 325200 322176 325252 322228
rect 343876 322176 343928 322228
rect 13964 322108 14016 322160
rect 16356 322108 16408 322160
rect 325384 322108 325436 322160
rect 347004 322108 347056 322160
rect 351236 322108 351288 322160
rect 342496 322040 342548 322092
rect 345256 322040 345308 322092
rect 325660 320748 325712 320800
rect 342496 320748 342548 320800
rect 342956 320748 343008 320800
rect 324740 320680 324792 320732
rect 346452 320680 346504 320732
rect 349488 320680 349540 320732
rect 62448 320612 62500 320664
rect 67692 320612 67744 320664
rect 150860 320612 150912 320664
rect 151964 320612 152016 320664
rect 156196 320612 156248 320664
rect 156932 320612 156984 320664
rect 158956 320612 159008 320664
rect 162636 320612 162688 320664
rect 243228 320612 243280 320664
rect 243780 320612 243832 320664
rect 245896 320612 245948 320664
rect 246448 320612 246500 320664
rect 63736 320544 63788 320596
rect 69440 320544 69492 320596
rect 154816 320544 154868 320596
rect 163464 320544 163516 320596
rect 244424 320544 244476 320596
rect 250956 320612 251008 320664
rect 337160 320612 337212 320664
rect 337528 320612 337580 320664
rect 339920 320612 339972 320664
rect 340564 320612 340616 320664
rect 58216 320476 58268 320528
rect 64104 320476 64156 320528
rect 57940 320408 57992 320460
rect 65116 320476 65168 320528
rect 243596 320476 243648 320528
rect 248932 320544 248984 320596
rect 332928 320544 332980 320596
rect 348568 320544 348620 320596
rect 352800 320544 352852 320596
rect 248656 320476 248708 320528
rect 249116 320476 249168 320528
rect 331456 320476 331508 320528
rect 340472 320476 340524 320528
rect 341024 320476 341076 320528
rect 65208 320408 65260 320460
rect 338448 320408 338500 320460
rect 352248 320476 352300 320528
rect 352892 320476 352944 320528
rect 59688 320340 59740 320392
rect 70636 320340 70688 320392
rect 336976 320340 337028 320392
rect 351604 320408 351656 320460
rect 56100 320272 56152 320324
rect 66588 320272 66640 320324
rect 248748 320272 248800 320324
rect 257120 320272 257172 320324
rect 335596 320272 335648 320324
rect 350408 320340 350460 320392
rect 350960 320272 351012 320324
rect 60608 320204 60660 320256
rect 71924 320204 71976 320256
rect 332836 320204 332888 320256
rect 348016 320204 348068 320256
rect 55272 320136 55324 320188
rect 62356 320136 62408 320188
rect 74776 320136 74828 320188
rect 246264 320136 246316 320188
rect 254544 320136 254596 320188
rect 325568 320136 325620 320188
rect 325844 320136 325896 320188
rect 347280 320136 347332 320188
rect 59596 320068 59648 320120
rect 65944 320068 65996 320120
rect 149296 320068 149348 320120
rect 155644 320068 155696 320120
rect 248932 320068 248984 320120
rect 259696 320068 259748 320120
rect 334308 320068 334360 320120
rect 349396 320068 349448 320120
rect 61436 320000 61488 320052
rect 73396 320000 73448 320052
rect 147916 320000 147968 320052
rect 161716 320000 161768 320052
rect 241756 320000 241808 320052
rect 255556 320000 255608 320052
rect 325108 320000 325160 320052
rect 325568 320000 325620 320052
rect 334216 320000 334268 320052
rect 349764 320000 349816 320052
rect 58768 319932 58820 319984
rect 70728 319932 70780 319984
rect 145340 319932 145392 319984
rect 159048 319932 159100 319984
rect 163004 319932 163056 319984
rect 164384 319932 164436 319984
rect 238996 319932 239048 319984
rect 252796 319932 252848 319984
rect 335688 319932 335740 319984
rect 349488 319932 349540 319984
rect 429436 319932 429488 319984
rect 66496 319864 66548 319916
rect 60976 319796 61028 319848
rect 66772 319796 66824 319848
rect 62448 319728 62500 319780
rect 68612 319728 68664 319780
rect 338540 319728 338592 319780
rect 339460 319728 339512 319780
rect 56836 319660 56888 319712
rect 63276 319660 63328 319712
rect 248840 319660 248892 319712
rect 251784 319660 251836 319712
rect 57020 319592 57072 319644
rect 338724 319592 338776 319644
rect 339644 319592 339696 319644
rect 58308 319524 58360 319576
rect 65024 319524 65076 319576
rect 253532 319524 253584 319576
rect 256292 319524 256344 319576
rect 152332 319456 152384 319508
rect 158128 319456 158180 319508
rect 341208 319456 341260 319508
rect 341760 319456 341812 319508
rect 65300 319388 65352 319440
rect 70360 319388 70412 319440
rect 325476 319388 325528 319440
rect 325844 319388 325896 319440
rect 342496 319388 342548 319440
rect 325292 319320 325344 319372
rect 345716 319320 345768 319372
rect 349488 319320 349540 319372
rect 325844 319252 325896 319304
rect 352892 316575 352944 316584
rect 352892 316541 352901 316575
rect 352901 316541 352935 316575
rect 352935 316541 352944 316575
rect 352892 316532 352944 316541
rect 38804 315852 38856 315904
rect 52696 315852 52748 315904
rect 357676 315852 357728 315904
rect 358320 315852 358372 315904
rect 405976 315852 406028 315904
rect 325292 314424 325344 314476
rect 430172 314424 430224 314476
rect 38436 313744 38488 313796
rect 51224 313744 51276 313796
rect 356204 313744 356256 313796
rect 405976 313744 406028 313796
rect 76984 313540 77036 313592
rect 81676 313540 81728 313592
rect 165120 313064 165172 313116
rect 175516 313064 175568 313116
rect 258960 313064 259012 313116
rect 270276 313064 270328 313116
rect 76156 312452 76208 312504
rect 76984 312452 77036 312504
rect 38804 310276 38856 310328
rect 54076 310276 54128 310328
rect 356940 310276 356992 310328
rect 405976 310276 406028 310328
rect 13964 309664 14016 309716
rect 16540 309664 16592 309716
rect 137704 309664 137756 309716
rect 145524 309664 145576 309716
rect 231452 309664 231504 309716
rect 240652 309664 240704 309716
rect 325384 309664 325436 309716
rect 334216 309664 334268 309716
rect 356296 309664 356348 309716
rect 356940 309664 356992 309716
rect 38804 308236 38856 308288
rect 51224 308236 51276 308288
rect 356204 308236 356256 308288
rect 405976 308236 406028 308288
rect 352892 306987 352944 306996
rect 352892 306953 352901 306987
rect 352901 306953 352935 306987
rect 352935 306953 352944 306987
rect 352892 306944 352944 306953
rect 38804 306196 38856 306248
rect 54444 306196 54496 306248
rect 354916 306196 354968 306248
rect 355652 306196 355704 306248
rect 406068 306196 406120 306248
rect 232096 304156 232148 304208
rect 232740 304156 232792 304208
rect 38620 304088 38672 304140
rect 51408 304088 51460 304140
rect 356204 304088 356256 304140
rect 405976 304088 406028 304140
rect 232004 301368 232056 301420
rect 233476 301368 233528 301420
rect 234120 301368 234172 301420
rect 352892 301436 352944 301488
rect 352800 301300 352852 301352
rect 38804 300620 38856 300672
rect 50304 300620 50356 300672
rect 355560 300620 355612 300672
rect 405976 300620 406028 300672
rect 355008 300008 355060 300060
rect 355560 300008 355612 300060
rect 38252 298580 38304 298632
rect 51408 298580 51460 298632
rect 356204 298580 356256 298632
rect 405976 298580 406028 298632
rect 74224 297152 74276 297204
rect 81676 297152 81728 297204
rect 167880 297152 167932 297204
rect 175516 297152 175568 297204
rect 261720 297152 261772 297204
rect 270368 297152 270420 297204
rect 13688 296132 13740 296184
rect 16724 296132 16776 296184
rect 137796 295860 137848 295912
rect 145432 295860 145484 295912
rect 231544 295860 231596 295912
rect 240928 295860 240980 295912
rect 325476 295860 325528 295912
rect 334216 295860 334268 295912
rect 353536 295792 353588 295844
rect 354180 295792 354232 295844
rect 38804 295112 38856 295164
rect 51316 295112 51368 295164
rect 353536 295112 353588 295164
rect 405976 295112 406028 295164
rect 38436 293752 38488 293804
rect 51316 293752 51368 293804
rect 356204 293752 356256 293804
rect 405976 293752 406028 293804
rect 14700 293140 14752 293192
rect 17460 293140 17512 293192
rect 38620 291644 38672 291696
rect 50028 291644 50080 291696
rect 50028 291236 50080 291288
rect 51684 291236 51736 291288
rect 353996 290964 354048 291016
rect 405976 290964 406028 291016
rect 427688 290352 427740 290404
rect 429436 290352 429488 290404
rect 427228 288992 427280 289044
rect 430264 288992 430316 289044
rect 38804 288924 38856 288976
rect 51316 288924 51368 288976
rect 356204 288924 356256 288976
rect 406068 288924 406120 288976
rect 51408 288720 51460 288772
rect 51684 288720 51736 288772
rect 261260 286272 261312 286324
rect 269264 286272 269316 286324
rect 168064 286204 168116 286256
rect 175424 286204 175476 286256
rect 38804 285456 38856 285508
rect 49936 285456 49988 285508
rect 354272 285456 354324 285508
rect 405976 285456 406028 285508
rect 38068 283416 38120 283468
rect 51500 283484 51552 283536
rect 137888 283484 137940 283536
rect 145156 283484 145208 283536
rect 231820 283484 231872 283536
rect 240376 283484 240428 283536
rect 325568 283484 325620 283536
rect 334216 283484 334268 283536
rect 356204 283416 356256 283468
rect 405976 283416 406028 283468
rect 12676 283348 12728 283400
rect 14700 283348 14752 283400
rect 142396 283348 142448 283400
rect 143040 283348 143092 283400
rect 236236 283008 236288 283060
rect 236880 283008 236932 283060
rect 325844 282804 325896 282856
rect 330076 282804 330128 282856
rect 231636 282736 231688 282788
rect 236236 282736 236288 282788
rect 138164 282328 138216 282380
rect 143040 282328 143092 282380
rect 16356 280628 16408 280680
rect 16724 280628 16776 280680
rect 74132 280628 74184 280680
rect 81676 280628 81728 280680
rect 427872 280628 427924 280680
rect 430172 280628 430224 280680
rect 38068 279948 38120 280000
rect 48556 279948 48608 280000
rect 352984 279379 353036 279388
rect 352984 279345 352993 279379
rect 352993 279345 353027 279379
rect 353027 279345 353036 279379
rect 352984 279336 353036 279345
rect 38620 279268 38672 279320
rect 51500 279268 51552 279320
rect 356204 279268 356256 279320
rect 405976 279268 406028 279320
rect 64196 276548 64248 276600
rect 64748 276548 64800 276600
rect 137520 275120 137572 275172
rect 155920 275120 155972 275172
rect 348752 275120 348804 275172
rect 138440 275052 138492 275104
rect 155276 275052 155328 275104
rect 234120 275052 234172 275104
rect 249116 275052 249168 275104
rect 347004 275052 347056 275104
rect 149204 274984 149256 275036
rect 158220 274984 158272 275036
rect 338264 274984 338316 275036
rect 349580 274984 349632 275036
rect 149756 274916 149808 274968
rect 160520 274916 160572 274968
rect 339644 274916 339696 274968
rect 351236 274916 351288 274968
rect 150584 274848 150636 274900
rect 162728 274848 162780 274900
rect 243504 274848 243556 274900
rect 252980 274848 253032 274900
rect 341024 274848 341076 274900
rect 352156 274848 352208 274900
rect 59688 274780 59740 274832
rect 60792 274780 60844 274832
rect 151872 274780 151924 274832
rect 163280 274780 163332 274832
rect 244056 274780 244108 274832
rect 254452 274780 254504 274832
rect 336884 274780 336936 274832
rect 34572 274712 34624 274764
rect 46992 274712 47044 274764
rect 149204 274712 149256 274764
rect 162084 274712 162136 274764
rect 243044 274712 243096 274764
rect 255740 274712 255792 274764
rect 334124 274712 334176 274764
rect 346176 274780 346228 274832
rect 343508 274712 343560 274764
rect 348200 274712 348252 274764
rect 31904 274644 31956 274696
rect 46624 274644 46676 274696
rect 147824 274644 147876 274696
rect 161440 274644 161492 274696
rect 241664 274644 241716 274696
rect 255096 274644 255148 274696
rect 335412 274644 335464 274696
rect 342404 274644 342456 274696
rect 345900 274644 345952 274696
rect 29236 274576 29288 274628
rect 46532 274576 46584 274628
rect 145064 274576 145116 274628
rect 160244 274576 160296 274628
rect 240284 274576 240336 274628
rect 254544 274576 254596 274628
rect 332744 274576 332796 274628
rect 26568 274508 26620 274560
rect 47084 274508 47136 274560
rect 146444 274508 146496 274560
rect 160888 274508 160940 274560
rect 238904 274508 238956 274560
rect 254176 274508 254228 274560
rect 335504 274508 335556 274560
rect 23900 274440 23952 274492
rect 46440 274440 46492 274492
rect 57020 274440 57072 274492
rect 68060 274440 68112 274492
rect 143684 274440 143736 274492
rect 159600 274440 159652 274492
rect 237524 274440 237576 274492
rect 253256 274440 253308 274492
rect 246540 274236 246592 274288
rect 247184 274236 247236 274288
rect 344336 274576 344388 274628
rect 349580 274576 349632 274628
rect 341760 274508 341812 274560
rect 345992 274508 346044 274560
rect 345164 274440 345216 274492
rect 367980 274440 368032 274492
rect 369912 274440 369964 274492
rect 410208 274440 410260 274492
rect 345348 274372 345400 274424
rect 348016 274236 348068 274288
rect 338172 274032 338224 274084
rect 342588 274032 342640 274084
rect 62356 273964 62408 274016
rect 63644 273964 63696 274016
rect 247276 273964 247328 274016
rect 247828 273964 247880 274016
rect 249576 273964 249628 274016
rect 339276 273964 339328 274016
rect 341944 273964 341996 274016
rect 254820 273896 254872 273948
rect 257580 273896 257632 273948
rect 337620 273896 337672 273948
rect 341116 273896 341168 273948
rect 61620 273828 61672 273880
rect 63276 273828 63328 273880
rect 64380 273828 64432 273880
rect 65944 273828 65996 273880
rect 151044 273828 151096 273880
rect 151964 273828 152016 273880
rect 234120 273828 234172 273880
rect 234764 273828 234816 273880
rect 256200 273828 256252 273880
rect 258316 273828 258368 273880
rect 340104 273828 340156 273880
rect 341852 273828 341904 273880
rect 21232 273760 21284 273812
rect 22244 273760 22296 273812
rect 61436 273760 61488 273812
rect 62264 273760 62316 273812
rect 63000 273760 63052 273812
rect 64104 273760 64156 273812
rect 65760 273760 65812 273812
rect 66772 273760 66824 273812
rect 68520 273760 68572 273812
rect 69440 273760 69492 273812
rect 152240 273760 152292 273812
rect 153252 273760 153304 273812
rect 153436 273760 153488 273812
rect 162360 273760 162412 273812
rect 163924 273760 163976 273812
rect 245344 273760 245396 273812
rect 245804 273760 245856 273812
rect 247736 273760 247788 273812
rect 248472 273760 248524 273812
rect 249024 273760 249076 273812
rect 249944 273760 249996 273812
rect 256292 273760 256344 273812
rect 256936 273760 256988 273812
rect 340932 273760 340984 273812
rect 341760 273760 341812 273812
rect 154724 273692 154776 273744
rect 352800 272400 352852 272452
rect 352984 272400 353036 272452
rect 349488 271720 349540 271772
rect 350408 271720 350460 271772
rect 12860 270020 12912 270072
rect 16448 270020 16500 270072
rect 88392 269612 88444 269664
rect 182416 269612 182468 269664
rect 182968 269612 183020 269664
rect 276440 269612 276492 269664
rect 290700 269612 290752 269664
rect 430080 269612 430132 269664
rect 13320 269544 13372 269596
rect 95476 269544 95528 269596
rect 96764 269544 96816 269596
rect 102652 269544 102704 269596
rect 196676 269544 196728 269596
rect 189408 269476 189460 269528
rect 283524 269476 283576 269528
rect 127768 269340 127820 269392
rect 131172 269340 131224 269392
rect 303764 269340 303816 269392
rect 304960 269340 305012 269392
rect 310756 269340 310808 269392
rect 312044 269340 312096 269392
rect 95568 269000 95620 269052
rect 109736 269000 109788 269052
rect 189316 269000 189368 269052
rect 203760 269000 203812 269052
rect 284536 269000 284588 269052
rect 297784 269000 297836 269052
rect 96764 268932 96816 268984
rect 170640 268932 170692 268984
rect 189408 268932 189460 268984
rect 196676 268932 196728 268984
rect 268620 268932 268672 268984
rect 290700 268932 290752 268984
rect 210016 268864 210068 268916
rect 210936 268864 210988 268916
rect 114796 268524 114848 268576
rect 116912 268524 116964 268576
rect 354916 267844 354968 267896
rect 355836 267844 355888 267896
rect 64840 266824 64892 266876
rect 68520 266824 68572 266876
rect 158220 266824 158272 266876
rect 158956 266824 159008 266876
rect 247644 266824 247696 266876
rect 254820 266824 254872 266876
rect 153160 266756 153212 266808
rect 162360 266756 162412 266808
rect 246264 266756 246316 266808
rect 256292 266756 256344 266808
rect 59688 266688 59740 266740
rect 63828 266688 63880 266740
rect 154724 266688 154776 266740
rect 164476 266688 164528 266740
rect 244884 266688 244936 266740
rect 255648 266688 255700 266740
rect 63644 266620 63696 266672
rect 75236 266620 75288 266672
rect 151964 266620 152016 266672
rect 62264 266552 62316 266604
rect 74224 266552 74276 266604
rect 150492 266552 150544 266604
rect 161716 266620 161768 266672
rect 245804 266620 245856 266672
rect 256936 266620 256988 266672
rect 244424 266552 244476 266604
rect 255556 266552 255608 266604
rect 60884 266484 60936 266536
rect 73120 266484 73172 266536
rect 143040 266484 143092 266536
rect 155736 266484 155788 266536
rect 247184 266484 247236 266536
rect 259696 266484 259748 266536
rect 341760 266484 341812 266536
rect 345808 266484 345860 266536
rect 59504 266416 59556 266468
rect 71096 266416 71148 266468
rect 153252 266416 153304 266468
rect 165948 266416 166000 266468
rect 245712 266416 245764 266468
rect 258408 266416 258460 266468
rect 58124 266348 58176 266400
rect 70084 266348 70136 266400
rect 151780 266348 151832 266400
rect 164568 266348 164620 266400
rect 236880 266348 236932 266400
rect 250036 266348 250088 266400
rect 56744 266280 56796 266332
rect 67968 266280 68020 266332
rect 154632 266280 154684 266332
rect 168708 266280 168760 266332
rect 248472 266280 248524 266332
rect 262456 266280 262508 266332
rect 55364 266212 55416 266264
rect 66956 266212 67008 266264
rect 153344 266212 153396 266264
rect 167328 266212 167380 266264
rect 247092 266212 247144 266264
rect 261076 266212 261128 266264
rect 60792 266144 60844 266196
rect 72108 266144 72160 266196
rect 154540 266144 154592 266196
rect 170088 266144 170140 266196
rect 248564 266144 248616 266196
rect 263836 266144 263888 266196
rect 338540 266144 338592 266196
rect 349488 266144 349540 266196
rect 163096 266076 163148 266128
rect 63828 266008 63880 266060
rect 67876 266008 67928 266060
rect 60700 265804 60752 265856
rect 64380 265804 64432 265856
rect 62816 265736 62868 265788
rect 66496 265736 66548 265788
rect 61804 265668 61856 265720
rect 65760 265668 65812 265720
rect 157852 265668 157904 265720
rect 165120 265668 165172 265720
rect 251876 265668 251928 265720
rect 258960 265668 259012 265720
rect 58676 265600 58728 265652
rect 63000 265600 63052 265652
rect 341852 265600 341904 265652
rect 344796 265600 344848 265652
rect 345900 265600 345952 265652
rect 347924 265600 347976 265652
rect 57664 265532 57716 265584
rect 61620 265532 61672 265584
rect 65944 265532 65996 265584
rect 69256 265532 69308 265584
rect 249024 265532 249076 265584
rect 256200 265532 256252 265584
rect 333388 265532 333440 265584
rect 334124 265532 334176 265584
rect 334400 265532 334452 265584
rect 335412 265532 335464 265584
rect 341944 265532 341996 265584
rect 343784 265532 343836 265584
rect 345992 265532 346044 265584
rect 346820 265532 346872 265584
rect 427596 265464 427648 265516
rect 429436 265464 429488 265516
rect 51316 265056 51368 265108
rect 52052 265056 52104 265108
rect 74040 264419 74092 264428
rect 74040 264385 74049 264419
rect 74049 264385 74083 264419
rect 74083 264385 74092 264419
rect 74040 264376 74092 264385
rect 78916 264036 78968 264088
rect 123260 264036 123312 264088
rect 124364 264036 124416 264088
rect 310756 264036 310808 264088
rect 328420 264036 328472 264088
rect 267240 263492 267292 263544
rect 310756 263492 310808 263544
rect 73948 263467 74000 263476
rect 73948 263433 73957 263467
rect 73957 263433 73991 263467
rect 73991 263433 74000 263467
rect 73948 263424 74000 263433
rect 124364 263424 124416 263476
rect 140280 263424 140332 263476
rect 249944 263424 249996 263476
rect 358412 263424 358464 263476
rect 369544 263356 369596 263408
rect 225840 262880 225892 262932
rect 233476 262880 233528 262932
rect 132000 262744 132052 262796
rect 139820 262744 139872 262796
rect 325200 262744 325252 262796
rect 325844 262744 325896 262796
rect 360712 262744 360764 262796
rect 46992 262676 47044 262728
rect 49200 262676 49252 262728
rect 228692 262608 228744 262660
rect 369728 262608 369780 262660
rect 13412 262540 13464 262592
rect 385276 262540 385328 262592
rect 360436 261996 360488 262048
rect 360804 261996 360856 262048
rect 422536 261996 422588 262048
rect 78916 261384 78968 261436
rect 87196 261384 87248 261436
rect 132092 261384 132144 261436
rect 140372 261384 140424 261436
rect 225748 261384 225800 261436
rect 233476 261384 233528 261436
rect 324648 261384 324700 261436
rect 327684 261384 327736 261436
rect 95568 261316 95620 261368
rect 96212 261316 96264 261368
rect 203852 261248 203904 261300
rect 209924 261248 209976 261300
rect 297876 261248 297928 261300
rect 303764 261248 303816 261300
rect 217192 260636 217244 260688
rect 225196 260636 225248 260688
rect 311216 260636 311268 260688
rect 319220 260636 319272 260688
rect 123536 260568 123588 260620
rect 127768 260568 127820 260620
rect 110196 260432 110248 260484
rect 114796 260432 114848 260484
rect 78916 260024 78968 260076
rect 85080 260024 85132 260076
rect 132460 260024 132512 260076
rect 140372 260024 140424 260076
rect 189316 260024 189368 260076
rect 190512 260024 190564 260076
rect 226208 260024 226260 260076
rect 233476 260024 233528 260076
rect 360620 259276 360672 259328
rect 419776 259276 419828 259328
rect 78916 258664 78968 258716
rect 84436 258664 84488 258716
rect 132184 258596 132236 258648
rect 140556 258596 140608 258648
rect 226300 258596 226352 258648
rect 233476 258596 233528 258648
rect 321060 258528 321112 258580
rect 324648 258528 324700 258580
rect 78916 257304 78968 257356
rect 81676 257304 81728 257356
rect 132276 257304 132328 257356
rect 140556 257304 140608 257356
rect 226484 257304 226536 257356
rect 232832 257304 232884 257356
rect 131356 257236 131408 257288
rect 140648 257236 140700 257288
rect 173124 257236 173176 257288
rect 181036 257236 181088 257288
rect 226116 257236 226168 257288
rect 233476 257236 233528 257288
rect 321060 257168 321112 257220
rect 327960 257168 328012 257220
rect 85080 256828 85132 256880
rect 87196 256828 87248 256880
rect 12860 256556 12912 256608
rect 16264 256556 16316 256608
rect 361172 256488 361224 256540
rect 417016 256488 417068 256540
rect 78916 255876 78968 255928
rect 81768 255876 81820 255928
rect 132368 255876 132420 255928
rect 139728 255876 139780 255928
rect 173308 255876 173360 255928
rect 176160 255876 176212 255928
rect 178276 255876 178328 255928
rect 181036 255876 181088 255928
rect 228692 255876 228744 255928
rect 233476 255876 233528 255928
rect 266596 255876 266648 255928
rect 271380 255876 271432 255928
rect 81676 255808 81728 255860
rect 87196 255808 87248 255860
rect 320600 255808 320652 255860
rect 327132 255808 327184 255860
rect 84436 255740 84488 255792
rect 87288 255740 87340 255792
rect 321612 255740 321664 255792
rect 327224 255740 327276 255792
rect 173584 255536 173636 255588
rect 222712 255536 222764 255588
rect 225840 255128 225892 255180
rect 225932 255128 225984 255180
rect 234580 255128 234632 255180
rect 225840 254924 225892 254976
rect 131356 254584 131408 254636
rect 136140 254584 136192 254636
rect 132000 254516 132052 254568
rect 136232 254516 136284 254568
rect 176344 254516 176396 254568
rect 181036 254516 181088 254568
rect 266596 254516 266648 254568
rect 272760 254516 272812 254568
rect 78916 254448 78968 254500
rect 82688 254448 82740 254500
rect 132552 254448 132604 254500
rect 140556 254448 140608 254500
rect 173308 254448 173360 254500
rect 176252 254448 176304 254500
rect 179196 254448 179248 254500
rect 181588 254448 181640 254500
rect 267884 254448 267936 254500
rect 274876 254448 274928 254500
rect 320508 254448 320560 254500
rect 328420 254448 328472 254500
rect 81768 254380 81820 254432
rect 87196 254380 87248 254432
rect 321612 253904 321664 253956
rect 328512 253904 328564 253956
rect 179012 253428 179064 253480
rect 181036 253428 181088 253480
rect 225748 253360 225800 253412
rect 234212 253360 234264 253412
rect 131356 253156 131408 253208
rect 137704 253156 137756 253208
rect 230072 253156 230124 253208
rect 233476 253156 233528 253208
rect 78916 253088 78968 253140
rect 137520 253088 137572 253140
rect 139820 253088 139872 253140
rect 266596 253088 266648 253140
rect 272852 253088 272904 253140
rect 361172 253020 361224 253072
rect 414256 253020 414308 253072
rect 427504 253020 427556 253072
rect 429436 253020 429488 253072
rect 87288 252952 87340 253004
rect 82688 252884 82740 252936
rect 87196 252884 87248 252936
rect 132276 252408 132328 252460
rect 267332 252340 267384 252392
rect 267792 252340 267844 252392
rect 132276 252204 132328 252256
rect 174044 251864 174096 251916
rect 178920 251864 178972 251916
rect 131356 251796 131408 251848
rect 138992 251796 139044 251848
rect 78916 251728 78968 251780
rect 132644 251728 132696 251780
rect 140556 251728 140608 251780
rect 174044 251728 174096 251780
rect 181588 251728 181640 251780
rect 230164 251728 230216 251780
rect 233568 251728 233620 251780
rect 266596 251728 266648 251780
rect 275980 251864 276032 251916
rect 321612 251864 321664 251916
rect 327132 251864 327184 251916
rect 271472 251728 271524 251780
rect 274876 251728 274928 251780
rect 87196 251592 87248 251644
rect 222804 250980 222856 251032
rect 233476 250980 233528 251032
rect 321612 250980 321664 251032
rect 327224 250980 327276 251032
rect 79744 250300 79796 250352
rect 87196 250300 87248 250352
rect 173584 250300 173636 250352
rect 182324 250300 182376 250352
rect 173492 250232 173544 250284
rect 181496 250232 181548 250284
rect 266596 250232 266648 250284
rect 276164 250232 276216 250284
rect 267424 250164 267476 250216
rect 274876 250164 274928 250216
rect 78916 249552 78968 249604
rect 87196 249552 87248 249604
rect 360712 249552 360764 249604
rect 412876 249552 412928 249604
rect 321060 249484 321112 249536
rect 327224 249484 327276 249536
rect 321612 249076 321664 249128
rect 328420 249076 328472 249128
rect 132000 248940 132052 248992
rect 138900 248940 138952 248992
rect 225840 248940 225892 248992
rect 234120 248940 234172 248992
rect 173400 248872 173452 248924
rect 181956 248872 182008 248924
rect 226576 248872 226628 248924
rect 233476 248872 233528 248924
rect 266596 248872 266648 248924
rect 274968 248872 275020 248924
rect 173768 248804 173820 248856
rect 181864 248804 181916 248856
rect 267516 248804 267568 248856
rect 274876 248804 274928 248856
rect 267608 248736 267660 248788
rect 274968 248736 275020 248788
rect 173492 248668 173544 248720
rect 178276 248668 178328 248720
rect 78916 248192 78968 248244
rect 87196 248192 87248 248244
rect 321612 247648 321664 247700
rect 328420 247648 328472 247700
rect 78916 247512 78968 247564
rect 88484 247512 88536 247564
rect 173860 247512 173912 247564
rect 182324 247512 182376 247564
rect 267792 247512 267844 247564
rect 274876 247512 274928 247564
rect 321796 247512 321848 247564
rect 328420 247512 328472 247564
rect 136232 247240 136284 247292
rect 140648 247240 140700 247292
rect 173308 246492 173360 246544
rect 179196 246492 179248 246544
rect 321428 246220 321480 246272
rect 78916 246152 78968 246204
rect 87196 246152 87248 246204
rect 131356 246152 131408 246204
rect 136140 246152 136192 246204
rect 140372 246152 140424 246204
rect 172756 246152 172808 246204
rect 176344 246152 176396 246204
rect 182324 246152 182376 246204
rect 226392 246152 226444 246204
rect 233476 246152 233528 246204
rect 267700 246152 267752 246204
rect 274876 246152 274928 246204
rect 327868 246152 327920 246204
rect 140556 246084 140608 246136
rect 176160 246084 176212 246136
rect 181588 246084 181640 246136
rect 266596 246084 266648 246136
rect 275796 246084 275848 246136
rect 173676 246016 173728 246068
rect 271380 246016 271432 246068
rect 274968 246016 275020 246068
rect 225564 245200 225616 245252
rect 228692 245200 228744 245252
rect 321704 244860 321756 244912
rect 323176 244860 323228 244912
rect 321612 244792 321664 244844
rect 78916 244724 78968 244776
rect 87196 244724 87248 244776
rect 137704 244724 137756 244776
rect 140096 244724 140148 244776
rect 176252 244724 176304 244776
rect 182324 244724 182376 244776
rect 225564 244724 225616 244776
rect 232740 244724 232792 244776
rect 266596 244724 266648 244776
rect 272760 244724 272812 244776
rect 274876 244724 274928 244776
rect 327868 244724 327920 244776
rect 275888 244588 275940 244640
rect 173124 243976 173176 244028
rect 179012 243976 179064 244028
rect 321612 243432 321664 243484
rect 327224 243432 327276 243484
rect 13136 243364 13188 243416
rect 16172 243364 16224 243416
rect 173952 243364 174004 243416
rect 181036 243364 181088 243416
rect 272852 243364 272904 243416
rect 275428 243364 275480 243416
rect 323176 243364 323228 243416
rect 327868 243364 327920 243416
rect 226484 243228 226536 243280
rect 233476 243228 233528 243280
rect 132552 243160 132604 243212
rect 137520 243160 137572 243212
rect 226484 243092 226536 243144
rect 230072 243092 230124 243144
rect 78916 243024 78968 243076
rect 87104 243024 87156 243076
rect 178920 242956 178972 243008
rect 181220 242956 181272 243008
rect 225748 242888 225800 242940
rect 230164 242888 230216 242940
rect 321612 242208 321664 242260
rect 328052 242208 328104 242260
rect 79100 242140 79152 242192
rect 87196 242140 87248 242192
rect 267884 242140 267936 242192
rect 271472 242140 271524 242192
rect 79008 242072 79060 242124
rect 87288 242072 87340 242124
rect 320508 242072 320560 242124
rect 327868 242072 327920 242124
rect 123076 241596 123128 241648
rect 124318 241596 124370 241648
rect 133380 240576 133432 240628
rect 140556 240576 140608 240628
rect 173584 240576 173636 240628
rect 181588 240576 181640 240628
rect 227220 240576 227272 240628
rect 233476 240576 233528 240628
rect 267884 240576 267936 240628
rect 275612 240576 275664 240628
rect 427412 240576 427464 240628
rect 429528 240576 429580 240628
rect 358596 239964 358648 240016
rect 389876 239964 389928 240016
rect 358504 239896 358556 239948
rect 393832 239896 393884 239948
rect 314896 239828 314948 239880
rect 316092 239828 316144 239880
rect 78916 239624 78968 239676
rect 87012 239624 87064 239676
rect 364484 239352 364536 239404
rect 377824 239352 377876 239404
rect 185636 239284 185688 239336
rect 186464 239284 186516 239336
rect 279660 239284 279712 239336
rect 280304 239284 280356 239336
rect 381872 239284 381924 239336
rect 132184 239216 132236 239268
rect 140556 239216 140608 239268
rect 173400 239216 173452 239268
rect 181956 239216 182008 239268
rect 226024 239216 226076 239268
rect 233476 239216 233528 239268
rect 267608 239216 267660 239268
rect 275704 239216 275756 239268
rect 266780 239148 266832 239200
rect 275520 239148 275572 239200
rect 200172 238536 200224 238588
rect 230900 238536 230952 238588
rect 290056 238536 290108 238588
rect 290516 238536 290568 238588
rect 325200 238536 325252 238588
rect 221056 237788 221108 237840
rect 222160 237788 222212 237840
rect 128136 237176 128188 237228
rect 140372 237176 140424 237228
rect 172940 237176 172992 237228
rect 219768 237176 219820 237228
rect 233476 237176 233528 237228
rect 267332 237176 267384 237228
rect 316276 237176 316328 237228
rect 78916 236564 78968 236616
rect 128136 236564 128188 236616
rect 316276 236564 316328 236616
rect 328420 236564 328472 236616
rect 296956 236292 297008 236344
rect 298244 236292 298296 236344
rect 262640 236156 262692 236208
rect 298244 235884 298296 235936
rect 324832 235884 324884 235936
rect 203116 235816 203168 235868
rect 230992 235816 231044 235868
rect 286928 235816 286980 235868
rect 325384 235816 325436 235868
rect 145340 235612 145392 235664
rect 146214 235612 146266 235664
rect 136876 235272 136928 235324
rect 137244 235272 137296 235324
rect 145156 235272 145208 235324
rect 152608 235272 152660 235324
rect 137060 235204 137112 235256
rect 150400 235204 150452 235256
rect 167696 235204 167748 235256
rect 149112 235136 149164 235188
rect 167972 235136 168024 235188
rect 230992 235136 231044 235188
rect 244976 235136 245028 235188
rect 262548 235136 262600 235188
rect 76064 235068 76116 235120
rect 113508 235068 113560 235120
rect 113876 235068 113928 235120
rect 359700 235068 359752 235120
rect 368716 235068 368768 235120
rect 113876 234388 113928 234440
rect 137336 234388 137388 234440
rect 301096 234388 301148 234440
rect 324924 234388 324976 234440
rect 346544 234388 346596 234440
rect 360620 234388 360672 234440
rect 324924 233776 324976 233828
rect 345256 233776 345308 233828
rect 346544 233776 346596 233828
rect 63644 233708 63696 233760
rect 61804 233572 61856 233624
rect 65760 233572 65812 233624
rect 62816 233504 62868 233556
rect 65852 233504 65904 233556
rect 138164 233708 138216 233760
rect 146812 233708 146864 233760
rect 149296 233708 149348 233760
rect 162268 233708 162320 233760
rect 234764 233708 234816 233760
rect 241480 233708 241532 233760
rect 246264 233708 246316 233760
rect 259236 233708 259288 233760
rect 323820 233708 323872 233760
rect 368716 233708 368768 233760
rect 154724 233640 154776 233692
rect 168064 233640 168116 233692
rect 248932 233640 248984 233692
rect 262088 233640 262140 233692
rect 243596 233572 243648 233624
rect 256292 233572 256344 233624
rect 362460 233572 362512 233624
rect 368808 233572 368860 233624
rect 75236 233504 75288 233556
rect 153344 233504 153396 233556
rect 166132 233504 166184 233556
rect 248012 233504 248064 233556
rect 261168 233504 261220 233556
rect 340932 233504 340984 233556
rect 347924 233504 347976 233556
rect 64840 233436 64892 233488
rect 67140 233436 67192 233488
rect 249944 233436 249996 233488
rect 263100 233436 263152 233488
rect 63828 233368 63880 233420
rect 67232 233368 67284 233420
rect 151964 233368 152016 233420
rect 165212 233368 165264 233420
rect 340840 233368 340892 233420
rect 346820 233368 346872 233420
rect 365220 233368 365272 233420
rect 368716 233368 368768 233420
rect 58124 233300 58176 233352
rect 70084 233300 70136 233352
rect 231452 233300 231504 233352
rect 234764 233300 234816 233352
rect 250680 233300 250732 233352
rect 264020 233300 264072 233352
rect 56744 233232 56796 233284
rect 67968 233232 68020 233284
rect 153712 233232 153764 233284
rect 167328 233232 167380 233284
rect 231728 233232 231780 233284
rect 243044 233232 243096 233284
rect 245344 233232 245396 233284
rect 258408 233232 258460 233284
rect 62264 233164 62316 233216
rect 74224 233164 74276 233216
rect 55364 233096 55416 233148
rect 66956 233096 67008 233148
rect 74132 233096 74184 233148
rect 60792 233028 60844 233080
rect 73120 233028 73172 233080
rect 137152 233096 137204 233148
rect 150676 233164 150728 233216
rect 151044 233164 151096 233216
rect 164568 233164 164620 233216
rect 231636 233164 231688 233216
rect 242124 233164 242176 233216
rect 244332 233164 244384 233216
rect 257304 233164 257356 233216
rect 144604 233096 144656 233148
rect 165120 233096 165172 233148
rect 238628 233096 238680 233148
rect 145248 233028 145300 233080
rect 156380 232960 156432 233012
rect 169996 232960 170048 233012
rect 59504 232892 59556 232944
rect 71096 232892 71148 232944
rect 155460 232892 155512 232944
rect 169076 232892 169128 232944
rect 60884 232824 60936 232876
rect 72108 232824 72160 232876
rect 150584 232824 150636 232876
rect 163280 232824 163332 232876
rect 109276 232756 109328 232808
rect 352892 233028 352944 233080
rect 247092 232892 247144 232944
rect 260156 232892 260208 232944
rect 258960 232824 259012 232876
rect 158864 232688 158916 232740
rect 161808 232688 161860 232740
rect 58676 232620 58728 232672
rect 63092 232620 63144 232672
rect 156104 232620 156156 232672
rect 158036 232620 158088 232672
rect 158128 232620 158180 232672
rect 160336 232620 160388 232672
rect 256016 232620 256068 232672
rect 258316 232620 258368 232672
rect 59688 232552 59740 232604
rect 63184 232552 63236 232604
rect 155184 232552 155236 232604
rect 157576 232552 157628 232604
rect 252704 232552 252756 232604
rect 255556 232552 255608 232604
rect 57664 232484 57716 232536
rect 61620 232484 61672 232536
rect 65944 232484 65996 232536
rect 68520 232484 68572 232536
rect 157116 232484 157168 232536
rect 159140 232484 159192 232536
rect 160060 232484 160112 232536
rect 162268 232484 162320 232536
rect 254084 232484 254136 232536
rect 255648 232484 255700 232536
rect 60700 232416 60752 232468
rect 63000 232416 63052 232468
rect 67324 232416 67376 232468
rect 68980 232416 69032 232468
rect 154264 232416 154316 232468
rect 156748 232416 156800 232468
rect 160980 232416 161032 232468
rect 163188 232416 163240 232468
rect 248288 232416 248340 232468
rect 250772 232416 250824 232468
rect 252152 232416 252204 232468
rect 254176 232416 254228 232468
rect 255004 232416 255056 232468
rect 256936 232416 256988 232468
rect 333388 232416 333440 232468
rect 334124 232416 334176 232468
rect 334400 232416 334452 232468
rect 335412 232416 335464 232468
rect 338540 232416 338592 232468
rect 339644 232416 339696 232468
rect 342680 232416 342732 232468
rect 344796 232416 344848 232468
rect 348108 232416 348160 232468
rect 349948 232416 350000 232468
rect 134852 232348 134904 232400
rect 368900 232348 368952 232400
rect 229980 232280 230032 232332
rect 368716 232280 368768 232332
rect 326580 232212 326632 232264
rect 368808 232212 368860 232264
rect 345716 231668 345768 231720
rect 360528 231668 360580 231720
rect 222620 230988 222672 231040
rect 222804 230988 222856 231040
rect 324832 230988 324884 231040
rect 325752 230988 325804 231040
rect 345440 230988 345492 231040
rect 345716 230988 345768 231040
rect 358320 231031 358372 231040
rect 358320 230997 358329 231031
rect 358329 230997 358363 231031
rect 358363 230997 358372 231031
rect 358320 230988 358372 230997
rect 47084 230920 47136 230972
rect 368900 230920 368952 230972
rect 76800 230852 76852 230904
rect 368716 230852 368768 230904
rect 134760 230784 134812 230836
rect 368808 230784 368860 230836
rect 115992 230376 116044 230428
rect 127216 230376 127268 230428
rect 210016 230376 210068 230428
rect 221056 230376 221108 230428
rect 304040 230376 304092 230428
rect 314896 230376 314948 230428
rect 103480 230308 103532 230360
rect 123076 230308 123128 230360
rect 197504 230308 197556 230360
rect 218296 230308 218348 230360
rect 291528 230308 291580 230360
rect 312136 230308 312188 230360
rect 91060 230240 91112 230292
rect 120316 230240 120368 230292
rect 185084 230240 185136 230292
rect 214156 230240 214208 230292
rect 279108 230240 279160 230292
rect 307996 230240 308048 230292
rect 343784 230240 343836 230292
rect 360896 230240 360948 230292
rect 324648 229628 324700 229680
rect 325476 229628 325528 229680
rect 343232 229628 343284 229680
rect 343784 229628 343836 229680
rect 13044 229560 13096 229612
rect 16080 229560 16132 229612
rect 22244 229560 22296 229612
rect 368716 229560 368768 229612
rect 370004 229016 370056 229068
rect 345256 228880 345308 228932
rect 346084 228880 346136 228932
rect 354916 228880 354968 228932
rect 355836 228880 355888 228932
rect 369820 228880 369872 228932
rect 370004 228880 370056 228932
rect 74040 228404 74092 228456
rect 368716 228404 368768 228456
rect 47084 228336 47136 228388
rect 368808 228336 368860 228388
rect 34020 228268 34072 228320
rect 368716 228268 368768 228320
rect 305144 227656 305196 227708
rect 322992 227656 323044 227708
rect 345164 227656 345216 227708
rect 360804 227656 360856 227708
rect 222436 227588 222488 227640
rect 222620 227588 222672 227640
rect 280304 227588 280356 227640
rect 353076 227588 353128 227640
rect 186464 227520 186516 227572
rect 369268 227520 369320 227572
rect 325384 226976 325436 227028
rect 325660 226976 325712 227028
rect 343876 226976 343928 227028
rect 345164 226976 345216 227028
rect 76800 226908 76852 226960
rect 368808 226908 368860 226960
rect 34572 226840 34624 226892
rect 368716 226840 368768 226892
rect 324740 226296 324792 226348
rect 347188 226296 347240 226348
rect 239548 226228 239600 226280
rect 353168 226228 353220 226280
rect 231360 226160 231412 226212
rect 353260 226160 353312 226212
rect 137612 226092 137664 226144
rect 353352 226092 353404 226144
rect 347188 225684 347240 225736
rect 359700 225820 359752 225872
rect 360436 225956 360488 226008
rect 172020 225616 172072 225668
rect 368808 225616 368860 225668
rect 137520 225548 137572 225600
rect 368716 225548 368768 225600
rect 134760 225480 134812 225532
rect 368900 225480 368952 225532
rect 158036 225412 158088 225464
rect 159048 225412 159100 225464
rect 161992 225412 162044 225464
rect 164384 225412 164436 225464
rect 251324 225412 251376 225464
rect 253992 225412 254044 225464
rect 338356 225412 338408 225464
rect 343508 225412 343560 225464
rect 350960 225412 351012 225464
rect 63000 225344 63052 225396
rect 65944 225344 65996 225396
rect 67140 225344 67192 225396
rect 69440 225344 69492 225396
rect 228692 225344 228744 225396
rect 368716 225344 368768 225396
rect 56100 225276 56152 225328
rect 56744 225276 56796 225328
rect 59688 225276 59740 225328
rect 60884 225276 60936 225328
rect 61436 225276 61488 225328
rect 62264 225276 62316 225328
rect 62356 225276 62408 225328
rect 63644 225276 63696 225328
rect 65760 225276 65812 225328
rect 66772 225276 66824 225328
rect 68520 225276 68572 225328
rect 70360 225276 70412 225328
rect 137612 225276 137664 225328
rect 368992 225276 369044 225328
rect 249208 225208 249260 225260
rect 252152 225208 252204 225260
rect 337160 225208 337212 225260
rect 341116 225208 341168 225260
rect 341208 225208 341260 225260
rect 352248 225208 352300 225260
rect 65852 225140 65904 225192
rect 67692 225140 67744 225192
rect 249760 225140 249812 225192
rect 253072 225140 253124 225192
rect 339000 225140 339052 225192
rect 342036 225140 342088 225192
rect 348108 225140 348160 225192
rect 63092 225072 63144 225124
rect 64104 225072 64156 225124
rect 337712 225072 337764 225124
rect 342496 225072 342548 225124
rect 58768 225004 58820 225056
rect 59504 225004 59556 225056
rect 335412 225004 335464 225056
rect 348568 225004 348620 225056
rect 332744 224936 332796 224988
rect 347280 224936 347332 224988
rect 360712 224936 360764 224988
rect 361172 224936 361224 224988
rect 334124 224868 334176 224920
rect 347924 224868 347976 224920
rect 335504 224800 335556 224852
rect 349396 224800 349448 224852
rect 57020 224732 57072 224784
rect 67324 224732 67376 224784
rect 339644 224732 339696 224784
rect 358044 224800 358096 224852
rect 358228 224800 358280 224852
rect 360988 224732 361040 224784
rect 339552 224664 339604 224716
rect 342680 224664 342732 224716
rect 345348 224596 345400 224648
rect 336884 224528 336936 224580
rect 349764 224528 349816 224580
rect 341392 224460 341444 224512
rect 348016 224460 348068 224512
rect 338264 224392 338316 224444
rect 350684 224392 350736 224444
rect 339460 224324 339512 224376
rect 351604 224324 351656 224376
rect 63184 224256 63236 224308
rect 65024 224256 65076 224308
rect 67232 224256 67284 224308
rect 68612 224256 68664 224308
rect 325844 224256 325896 224308
rect 345164 224256 345216 224308
rect 61620 224188 61672 224240
rect 63276 224188 63328 224240
rect 324924 224188 324976 224240
rect 325200 224188 325252 224240
rect 344520 224188 344572 224240
rect 361172 224188 361224 224240
rect 322532 224120 322584 224172
rect 368808 224120 368860 224172
rect 369176 224163 369228 224172
rect 369176 224129 369185 224163
rect 369185 224129 369219 224163
rect 369219 224129 369228 224163
rect 369176 224120 369228 224129
rect 369084 223984 369136 224036
rect 369360 223984 369412 224036
rect 342726 223032 342778 223084
rect 325568 222896 325620 222948
rect 342726 222896 342778 222948
rect 362460 222896 362512 222948
rect 369084 222896 369136 222948
rect 323820 222828 323872 222880
rect 368716 222828 368768 222880
rect 322624 222760 322676 222812
rect 368808 222760 368860 222812
rect 38528 222012 38580 222064
rect 50580 222012 50632 222064
rect 34572 221740 34624 221792
rect 34940 221740 34992 221792
rect 34020 221672 34072 221724
rect 34756 221672 34808 221724
rect 361080 221468 361132 221520
rect 369084 221468 369136 221520
rect 325200 221400 325252 221452
rect 368808 221400 368860 221452
rect 322808 221332 322860 221384
rect 368716 221332 368768 221384
rect 369912 221375 369964 221384
rect 369912 221341 369921 221375
rect 369921 221341 369955 221375
rect 369955 221341 369964 221375
rect 369912 221332 369964 221341
rect 325292 220584 325344 220636
rect 353444 220584 353496 220636
rect 34664 220516 34716 220568
rect 34940 220516 34992 220568
rect 325384 220516 325436 220568
rect 368808 220516 368860 220568
rect 34756 220448 34808 220500
rect 322716 220448 322768 220500
rect 368716 220448 368768 220500
rect 359792 220040 359844 220092
rect 368992 220040 369044 220092
rect 38068 219904 38120 219956
rect 52052 219904 52104 219956
rect 76156 219496 76208 219548
rect 81676 219496 81728 219548
rect 165120 219224 165172 219276
rect 178920 219224 178972 219276
rect 258960 219224 259012 219276
rect 272944 219224 272996 219276
rect 365220 218680 365272 218732
rect 368808 218680 368860 218732
rect 352800 218612 352852 218664
rect 368716 218612 368768 218664
rect 394844 218612 394896 218664
rect 405976 218612 406028 218664
rect 352892 218544 352944 218596
rect 368808 218544 368860 218596
rect 352984 217184 353036 217236
rect 368716 217184 368768 217236
rect 38528 217116 38580 217168
rect 53248 217116 53300 217168
rect 353352 217048 353404 217100
rect 368716 217048 368768 217100
rect 368992 216436 369044 216488
rect 137704 215824 137756 215876
rect 145156 215824 145208 215876
rect 231360 215824 231412 215876
rect 240928 215824 240980 215876
rect 325292 215824 325344 215876
rect 334216 215824 334268 215876
rect 353168 215756 353220 215808
rect 368716 215756 368768 215808
rect 427320 215756 427372 215808
rect 429712 215756 429764 215808
rect 353260 215688 353312 215740
rect 368808 215688 368860 215740
rect 358412 215620 358464 215672
rect 368716 215620 368768 215672
rect 358228 215484 358280 215536
rect 358412 215484 358464 215536
rect 368992 214464 369044 214516
rect 369176 214464 369228 214516
rect 38528 214396 38580 214448
rect 51408 214396 51460 214448
rect 353076 214260 353128 214312
rect 368716 214260 368768 214312
rect 361264 214192 361316 214244
rect 368900 214192 368952 214244
rect 356204 214056 356256 214108
rect 405976 214056 406028 214108
rect 357676 213988 357728 214040
rect 406620 213988 406672 214040
rect 355100 213920 355152 213972
rect 394844 213920 394896 213972
rect 34848 213895 34900 213904
rect 34848 213861 34857 213895
rect 34857 213861 34891 213895
rect 34891 213861 34900 213895
rect 34848 213852 34900 213861
rect 353444 213036 353496 213088
rect 368716 213036 368768 213088
rect 369912 211608 369964 211660
rect 370740 211608 370792 211660
rect 38712 210928 38764 210980
rect 54076 210928 54128 210980
rect 354916 210928 354968 210980
rect 405976 210928 406028 210980
rect 383896 210860 383948 210912
rect 385184 210860 385236 210912
rect 369544 209636 369596 209688
rect 369912 209636 369964 209688
rect 38528 209568 38580 209620
rect 51408 209568 51460 209620
rect 356204 209568 356256 209620
rect 405976 209568 406028 209620
rect 34848 206891 34900 206900
rect 34848 206857 34857 206891
rect 34857 206857 34891 206891
rect 34891 206857 34900 206891
rect 34848 206848 34900 206857
rect 38528 206780 38580 206832
rect 51408 206780 51460 206832
rect 355008 206780 355060 206832
rect 405976 206780 406028 206832
rect 38528 204740 38580 204792
rect 51408 204740 51460 204792
rect 136876 204740 136928 204792
rect 145340 204740 145392 204792
rect 356204 204740 356256 204792
rect 406068 204740 406120 204792
rect 34848 204715 34900 204724
rect 34848 204681 34857 204715
rect 34857 204681 34891 204715
rect 34891 204681 34900 204715
rect 34848 204672 34900 204681
rect 368992 204672 369044 204724
rect 369176 204672 369228 204724
rect 231636 204060 231688 204112
rect 237524 204060 237576 204112
rect 74224 203312 74276 203364
rect 81676 203312 81728 203364
rect 167880 203312 167932 203364
rect 178920 203312 178972 203364
rect 261720 203312 261772 203364
rect 272944 203312 272996 203364
rect 13964 202020 14016 202072
rect 16448 202020 16500 202072
rect 137796 202020 137848 202072
rect 145156 202020 145208 202072
rect 231452 202020 231504 202072
rect 240376 202020 240428 202072
rect 325476 202020 325528 202072
rect 334216 202020 334268 202072
rect 358412 202020 358464 202072
rect 358596 202020 358648 202072
rect 38528 201272 38580 201324
rect 51500 201272 51552 201324
rect 353536 201272 353588 201324
rect 405976 201272 406028 201324
rect 369544 199912 369596 199964
rect 369912 199912 369964 199964
rect 427136 199708 427188 199760
rect 428792 199708 428844 199760
rect 13412 199300 13464 199352
rect 17644 199300 17696 199352
rect 38528 199232 38580 199284
rect 51224 199232 51276 199284
rect 356204 199232 356256 199284
rect 405976 199232 406028 199284
rect 38528 195764 38580 195816
rect 51316 195764 51368 195816
rect 352708 195764 352760 195816
rect 405976 195764 406028 195816
rect 368808 195220 368860 195272
rect 38804 195084 38856 195136
rect 51316 195152 51368 195204
rect 369084 195152 369136 195204
rect 369360 195152 369412 195204
rect 356204 195084 356256 195136
rect 406068 195084 406120 195136
rect 167972 192568 168024 192620
rect 173400 192568 173452 192620
rect 262364 192364 262416 192416
rect 273128 192364 273180 192416
rect 368716 192407 368768 192416
rect 368716 192373 368725 192407
rect 368725 192373 368759 192407
rect 368759 192373 368768 192407
rect 368716 192364 368768 192373
rect 38804 191616 38856 191668
rect 49936 191616 49988 191668
rect 173400 191616 173452 191668
rect 178920 191616 178972 191668
rect 352800 191616 352852 191668
rect 405976 191616 406028 191668
rect 368992 190256 369044 190308
rect 369360 190256 369412 190308
rect 369544 190256 369596 190308
rect 369912 190256 369964 190308
rect 13320 189576 13372 189628
rect 13504 189576 13556 189628
rect 38068 189576 38120 189628
rect 51224 189576 51276 189628
rect 137336 189576 137388 189628
rect 137704 189576 137756 189628
rect 356204 189576 356256 189628
rect 405976 189576 406028 189628
rect 13320 189372 13372 189424
rect 17460 189372 17512 189424
rect 324556 188896 324608 188948
rect 330076 188896 330128 188948
rect 232004 188760 232056 188812
rect 236236 188760 236288 188812
rect 236880 188760 236932 188812
rect 137796 188284 137848 188336
rect 142396 188284 142448 188336
rect 143040 188284 143092 188336
rect 232740 188284 232792 188336
rect 240376 188284 240428 188336
rect 138900 188216 138952 188268
rect 145616 188216 145668 188268
rect 326580 188216 326632 188268
rect 334216 188216 334268 188268
rect 75420 186788 75472 186840
rect 81676 186788 81728 186840
rect 38068 186108 38120 186160
rect 48556 186108 48608 186160
rect 352800 186108 352852 186160
rect 405976 186108 406028 186160
rect 368716 185496 368768 185548
rect 13504 185428 13556 185480
rect 17460 185428 17512 185480
rect 427228 185428 427280 185480
rect 430080 185428 430132 185480
rect 368808 185360 368860 185412
rect 38804 184000 38856 184052
rect 51408 184000 51460 184052
rect 356204 184000 356256 184052
rect 405976 184000 406028 184052
rect 34388 183184 34440 183236
rect 34940 183184 34992 183236
rect 34572 182640 34624 182692
rect 34756 182640 34808 182692
rect 352156 181688 352208 181740
rect 21600 181280 21652 181332
rect 34388 181280 34440 181332
rect 59688 181280 59740 181332
rect 60884 181280 60936 181332
rect 61436 181280 61488 181332
rect 62264 181280 62316 181332
rect 63000 181280 63052 181332
rect 64104 181280 64156 181332
rect 65760 181280 65812 181332
rect 66772 181280 66824 181332
rect 151044 181280 151096 181332
rect 151872 181280 151924 181332
rect 152240 181280 152292 181332
rect 153252 181280 153304 181332
rect 153436 181280 153488 181332
rect 154724 181280 154776 181332
rect 245344 181280 245396 181332
rect 245804 181280 245856 181332
rect 252060 181280 252112 181332
rect 257580 181280 257632 181332
rect 337620 181280 337672 181332
rect 341116 181280 341168 181332
rect 345164 181280 345216 181332
rect 359792 181280 359844 181332
rect 361172 181280 361224 181332
rect 412876 181280 412928 181332
rect 149204 181144 149256 181196
rect 158220 181144 158272 181196
rect 149756 181076 149808 181128
rect 160336 181076 160388 181128
rect 150584 181008 150636 181060
rect 162728 181008 162780 181060
rect 243504 181008 243556 181060
rect 252796 181008 252848 181060
rect 151964 180940 152016 180992
rect 163280 180940 163332 180992
rect 244056 180940 244108 180992
rect 254176 180940 254228 180992
rect 334124 180940 334176 180992
rect 346176 181212 346228 181264
rect 370740 181212 370792 181264
rect 410208 181212 410260 181264
rect 338264 181144 338316 181196
rect 341852 181144 341904 181196
rect 340104 181076 340156 181128
rect 343876 181076 343928 181128
rect 336884 181008 336936 181060
rect 348752 181008 348804 181060
rect 339644 180940 339696 180992
rect 351236 180940 351288 180992
rect 34664 180872 34716 180924
rect 46992 180872 47044 180924
rect 149204 180872 149256 180924
rect 162084 180872 162136 180924
rect 243044 180872 243096 180924
rect 255740 180872 255792 180924
rect 31812 180804 31864 180856
rect 45796 180804 45848 180856
rect 147824 180804 147876 180856
rect 161440 180804 161492 180856
rect 240284 180804 240336 180856
rect 254544 180804 254596 180856
rect 341024 180804 341076 180856
rect 29512 180736 29564 180788
rect 46624 180736 46676 180788
rect 145064 180736 145116 180788
rect 160244 180736 160296 180788
rect 241664 180736 241716 180788
rect 255096 180736 255148 180788
rect 335412 180736 335464 180788
rect 347004 180736 347056 180788
rect 26936 180668 26988 180720
rect 46532 180668 46584 180720
rect 238904 180668 238956 180720
rect 254268 180668 254320 180720
rect 332744 180668 332796 180720
rect 345348 180668 345400 180720
rect 24176 180600 24228 180652
rect 46440 180600 46492 180652
rect 57020 180600 57072 180652
rect 68060 180600 68112 180652
rect 146444 180600 146496 180652
rect 160888 180600 160940 180652
rect 237524 180600 237576 180652
rect 253440 180600 253492 180652
rect 335504 180600 335556 180652
rect 348016 180600 348068 180652
rect 143684 180532 143736 180584
rect 159600 180532 159652 180584
rect 338264 180532 338316 180584
rect 349580 180532 349632 180584
rect 62356 180464 62408 180516
rect 63644 180464 63696 180516
rect 68520 180464 68572 180516
rect 69440 180464 69492 180516
rect 247736 180464 247788 180516
rect 248564 180464 248616 180516
rect 339276 180464 339328 180516
rect 341760 180464 341812 180516
rect 340932 180396 340984 180448
rect 344612 180396 344664 180448
rect 246540 180328 246592 180380
rect 247184 180328 247236 180380
rect 343508 180124 343560 180176
rect 348016 180124 348068 180176
rect 341668 180056 341720 180108
rect 344704 180056 344756 180108
rect 344336 179988 344388 180040
rect 347280 179988 347332 180040
rect 254820 179920 254872 179972
rect 258408 179920 258460 179972
rect 342404 179920 342456 179972
rect 344520 179920 344572 179972
rect 368992 179920 369044 179972
rect 369360 179920 369412 179972
rect 369544 179920 369596 179972
rect 369912 179920 369964 179972
rect 324556 179852 324608 179904
rect 326580 179852 326632 179904
rect 230992 179716 231044 179768
rect 232740 179716 232792 179768
rect 427596 178492 427648 178544
rect 429896 178492 429948 178544
rect 368532 177880 368584 177932
rect 368716 177880 368768 177932
rect 358320 175908 358372 175960
rect 88392 175772 88444 175824
rect 178276 175772 178328 175824
rect 182416 175772 182468 175824
rect 182876 175772 182928 175824
rect 276440 175772 276492 175824
rect 358320 175772 358372 175824
rect 95476 175704 95528 175756
rect 170640 175704 170692 175756
rect 189500 175704 189552 175756
rect 283524 175704 283576 175756
rect 196676 175636 196728 175688
rect 268620 175636 268672 175688
rect 290700 175636 290752 175688
rect 96764 175160 96816 175212
rect 109736 175160 109788 175212
rect 190604 175160 190656 175212
rect 203760 175160 203812 175212
rect 102652 175092 102704 175144
rect 176160 175092 176212 175144
rect 196676 175092 196728 175144
rect 285824 175092 285876 175144
rect 297784 175092 297836 175144
rect 124364 174412 124416 174464
rect 131172 174412 131224 174464
rect 60700 172984 60752 173036
rect 65944 172984 65996 173036
rect 153160 172984 153212 173036
rect 153344 172984 153396 173036
rect 158220 172984 158272 173036
rect 158956 172984 159008 173036
rect 249024 172984 249076 173036
rect 254820 172984 254872 173036
rect 333388 172984 333440 173036
rect 334124 172984 334176 173036
rect 341852 172984 341904 173036
rect 342680 172984 342732 173036
rect 347280 172984 347332 173036
rect 349948 172984 350000 173036
rect 64840 172916 64892 172968
rect 68520 172916 68572 172968
rect 154540 172916 154592 172968
rect 164660 172916 164712 172968
rect 246264 172916 246316 172968
rect 257304 172916 257356 172968
rect 341760 172916 341812 172968
rect 343784 172916 343836 172968
rect 59688 172848 59740 172900
rect 65024 172848 65076 172900
rect 153344 172848 153396 172900
rect 163924 172848 163976 172900
rect 244884 172848 244936 172900
rect 256752 172848 256804 172900
rect 63644 172780 63696 172832
rect 75236 172780 75288 172832
rect 150308 172780 150360 172832
rect 161716 172780 161768 172832
rect 245804 172780 245856 172832
rect 256936 172780 256988 172832
rect 60884 172712 60936 172764
rect 72108 172712 72160 172764
rect 151872 172712 151924 172764
rect 163096 172712 163148 172764
rect 244424 172712 244476 172764
rect 255556 172712 255608 172764
rect 62264 172644 62316 172696
rect 74224 172644 74276 172696
rect 143040 172644 143092 172696
rect 155736 172644 155788 172696
rect 157852 172644 157904 172696
rect 165120 172644 165172 172696
rect 247184 172644 247236 172696
rect 259696 172644 259748 172696
rect 59504 172576 59556 172628
rect 71096 172576 71148 172628
rect 153252 172576 153304 172628
rect 165856 172576 165908 172628
rect 246816 172576 246868 172628
rect 258316 172576 258368 172628
rect 354916 172576 354968 172628
rect 355836 172576 355888 172628
rect 58032 172508 58084 172560
rect 70084 172508 70136 172560
rect 151688 172508 151740 172560
rect 164476 172508 164528 172560
rect 236880 172508 236932 172560
rect 250036 172508 250088 172560
rect 55364 172440 55416 172492
rect 66956 172440 67008 172492
rect 154724 172440 154776 172492
rect 168616 172440 168668 172492
rect 247644 172440 247696 172492
rect 252060 172440 252112 172492
rect 56744 172372 56796 172424
rect 67968 172372 68020 172424
rect 153160 172372 153212 172424
rect 167236 172372 167288 172424
rect 248564 172372 248616 172424
rect 262456 172440 262508 172492
rect 261168 172372 261220 172424
rect 60608 172304 60660 172356
rect 73120 172304 73172 172356
rect 154632 172304 154684 172356
rect 169996 172304 170048 172356
rect 248012 172304 248064 172356
rect 263836 172304 263888 172356
rect 338540 172304 338592 172356
rect 350684 172304 350736 172356
rect 63828 172236 63880 172288
rect 68612 172236 68664 172288
rect 245528 172236 245580 172288
rect 58676 172032 58728 172084
rect 63000 172032 63052 172084
rect 65944 172032 65996 172084
rect 70452 172032 70504 172084
rect 334400 172032 334452 172084
rect 335412 172032 335464 172084
rect 57664 171896 57716 171948
rect 63276 171896 63328 171948
rect 62816 171828 62868 171880
rect 67692 171828 67744 171880
rect 344520 171828 344572 171880
rect 347924 171828 347976 171880
rect 344704 171760 344756 171812
rect 346820 171760 346872 171812
rect 61804 171692 61856 171744
rect 65760 171692 65812 171744
rect 251876 171692 251928 171744
rect 258960 171692 259012 171744
rect 344612 171692 344664 171744
rect 345808 171692 345860 171744
rect 358412 171556 358464 171608
rect 358596 171556 358648 171608
rect 79744 170196 79796 170248
rect 123996 170196 124048 170248
rect 312044 170196 312096 170248
rect 328420 170196 328472 170248
rect 123996 169516 124048 169568
rect 140280 169516 140332 169568
rect 267240 169516 267292 169568
rect 312044 169516 312096 169568
rect 71648 169423 71700 169432
rect 71648 169389 71657 169423
rect 71657 169389 71691 169423
rect 71691 169389 71700 169423
rect 71648 169380 71700 169389
rect 132184 168904 132236 168956
rect 140556 168904 140608 168956
rect 225840 168904 225892 168956
rect 233476 168904 233528 168956
rect 46992 168836 47044 168888
rect 49200 168836 49252 168888
rect 359700 168836 359752 168888
rect 423640 168836 423692 168888
rect 222160 168564 222212 168616
rect 369268 168564 369320 168616
rect 128136 168496 128188 168548
rect 368992 168496 369044 168548
rect 368716 168156 368768 168208
rect 368992 168156 369044 168208
rect 77260 167544 77312 167596
rect 87196 167544 87248 167596
rect 132276 167544 132328 167596
rect 140556 167544 140608 167596
rect 226024 167544 226076 167596
rect 233476 167544 233528 167596
rect 203852 166932 203904 166984
rect 210936 166932 210988 166984
rect 110196 166796 110248 166848
rect 116912 166796 116964 166848
rect 217192 166796 217244 166848
rect 225196 166796 225248 166848
rect 297876 166796 297928 166848
rect 304960 166796 305012 166848
rect 311216 166796 311268 166848
rect 319220 166796 319272 166848
rect 123536 166320 123588 166372
rect 124364 166320 124416 166372
rect 284536 166252 284588 166304
rect 285824 166252 285876 166304
rect 77260 166184 77312 166236
rect 85724 166184 85776 166236
rect 132092 166184 132144 166236
rect 140556 166184 140608 166236
rect 225932 166184 225984 166236
rect 233476 166184 233528 166236
rect 324556 166184 324608 166236
rect 328420 166184 328472 166236
rect 361264 165436 361316 165488
rect 420880 165436 420932 165488
rect 79744 164824 79796 164876
rect 85632 164824 85684 164876
rect 132552 164756 132604 164808
rect 139636 164756 139688 164808
rect 225748 164756 225800 164808
rect 233476 164756 233528 164808
rect 321796 164756 321848 164808
rect 328512 164756 328564 164808
rect 132644 163464 132696 163516
rect 139636 163464 139688 163516
rect 226300 163464 226352 163516
rect 232832 163464 232884 163516
rect 321612 163464 321664 163516
rect 327224 163464 327276 163516
rect 131356 163396 131408 163448
rect 140556 163396 140608 163448
rect 179012 163396 179064 163448
rect 182324 163396 182376 163448
rect 226116 163396 226168 163448
rect 233476 163396 233528 163448
rect 85724 163328 85776 163380
rect 87196 163328 87248 163380
rect 320968 163328 321020 163380
rect 324556 163328 324608 163380
rect 358596 163371 358648 163380
rect 358596 163337 358605 163371
rect 358605 163337 358639 163371
rect 358639 163337 358648 163371
rect 358596 163328 358648 163337
rect 12860 163192 12912 163244
rect 16356 163192 16408 163244
rect 360528 162648 360580 162700
rect 418212 162648 418264 162700
rect 226300 162376 226352 162428
rect 230992 162376 231044 162428
rect 132000 162104 132052 162156
rect 138164 162104 138216 162156
rect 131908 162036 131960 162088
rect 139636 162036 139688 162088
rect 178828 162036 178880 162088
rect 181772 162036 181824 162088
rect 226300 162036 226352 162088
rect 233476 162036 233528 162088
rect 266872 162036 266924 162088
rect 274876 162036 274928 162088
rect 321704 162036 321756 162088
rect 328420 162036 328472 162088
rect 77260 161968 77312 162020
rect 87196 161968 87248 162020
rect 132000 161968 132052 162020
rect 132276 161968 132328 162020
rect 85632 161900 85684 161952
rect 87288 161900 87340 161952
rect 222436 161560 222488 161612
rect 172848 161492 172900 161544
rect 320784 161288 320836 161340
rect 327224 161288 327276 161340
rect 131356 160676 131408 160728
rect 140464 160676 140516 160728
rect 131724 160608 131776 160660
rect 139636 160608 139688 160660
rect 173952 160608 174004 160660
rect 177540 160608 177592 160660
rect 179104 160608 179156 160660
rect 182324 160608 182376 160660
rect 226392 160608 226444 160660
rect 232924 160744 232976 160796
rect 266964 160744 267016 160796
rect 267332 160744 267384 160796
rect 274876 160744 274928 160796
rect 266596 160676 266648 160728
rect 274324 160676 274376 160728
rect 231360 160608 231412 160660
rect 233476 160608 233528 160660
rect 267332 160608 267384 160660
rect 271380 160608 271432 160660
rect 274876 160608 274928 160660
rect 77168 160540 77220 160592
rect 87196 160540 87248 160592
rect 225564 159928 225616 159980
rect 226300 159928 226352 159980
rect 173952 159316 174004 159368
rect 180392 159316 180444 159368
rect 226300 159316 226352 159368
rect 232740 159316 232792 159368
rect 79284 159248 79336 159300
rect 137612 159248 137664 159300
rect 139636 159248 139688 159300
rect 178920 159248 178972 159300
rect 182324 159248 182376 159300
rect 227220 159248 227272 159300
rect 233476 159248 233528 159300
rect 266596 159248 266648 159300
rect 274232 159248 274284 159300
rect 87288 159112 87340 159164
rect 81676 159044 81728 159096
rect 87196 159044 87248 159096
rect 361264 158500 361316 158552
rect 415544 158500 415596 158552
rect 321612 158160 321664 158212
rect 327224 158160 327276 158212
rect 321060 158024 321112 158076
rect 327316 158024 327368 158076
rect 131356 157956 131408 158008
rect 138900 157956 138952 158008
rect 173860 157956 173912 158008
rect 79744 157888 79796 157940
rect 87196 157888 87248 157940
rect 131632 157888 131684 157940
rect 139636 157888 139688 157940
rect 173768 157888 173820 157940
rect 176252 157888 176304 157940
rect 226392 157956 226444 158008
rect 228784 157956 228836 158008
rect 266596 157956 266648 158008
rect 274416 157956 274468 158008
rect 182324 157888 182376 157940
rect 227312 157888 227364 157940
rect 233476 157888 233528 157940
rect 321612 157208 321664 157260
rect 327224 157208 327276 157260
rect 222804 157140 222856 157192
rect 233476 157140 233528 157192
rect 77260 156460 77312 156512
rect 173768 156460 173820 156512
rect 181772 156460 181824 156512
rect 87196 156392 87248 156444
rect 173584 156392 173636 156444
rect 182324 156392 182376 156444
rect 267424 156392 267476 156444
rect 274876 156392 274928 156444
rect 358596 156435 358648 156444
rect 358596 156401 358605 156435
rect 358605 156401 358639 156435
rect 358639 156401 358648 156435
rect 358596 156392 358648 156401
rect 321612 155916 321664 155968
rect 327224 155916 327276 155968
rect 173952 155100 174004 155152
rect 182232 155100 182284 155152
rect 267792 155100 267844 155152
rect 274968 155100 275020 155152
rect 321612 155100 321664 155152
rect 79744 155032 79796 155084
rect 87196 155032 87248 155084
rect 138164 155032 138216 155084
rect 139728 155032 139780 155084
rect 174044 155032 174096 155084
rect 179012 155032 179064 155084
rect 173400 154964 173452 155016
rect 181128 155032 181180 155084
rect 230992 155032 231044 155084
rect 234028 155032 234080 155084
rect 267700 155032 267752 155084
rect 274876 155032 274928 155084
rect 328420 155032 328472 155084
rect 266596 154964 266648 155016
rect 274508 154964 274560 155016
rect 267056 154896 267108 154948
rect 267700 154896 267752 154948
rect 79744 154352 79796 154404
rect 87196 154352 87248 154404
rect 172940 153876 172992 153928
rect 178828 153876 178880 153928
rect 368532 153808 368584 153860
rect 368992 153808 369044 153860
rect 320876 153740 320928 153792
rect 328420 153740 328472 153792
rect 131540 153672 131592 153724
rect 139636 153672 139688 153724
rect 173308 153672 173360 153724
rect 181404 153672 181456 153724
rect 267148 153672 267200 153724
rect 274968 153672 275020 153724
rect 427504 153672 427556 153724
rect 429436 153672 429488 153724
rect 173492 153604 173544 153656
rect 181956 153604 182008 153656
rect 267516 153604 267568 153656
rect 274876 153604 274928 153656
rect 173216 153128 173268 153180
rect 179104 153128 179156 153180
rect 79744 152992 79796 153044
rect 87196 152992 87248 153044
rect 320508 152448 320560 152500
rect 323176 152448 323228 152500
rect 85816 152380 85868 152432
rect 87196 152380 87248 152432
rect 321612 152380 321664 152432
rect 328420 152380 328472 152432
rect 174044 152312 174096 152364
rect 182324 152312 182376 152364
rect 267884 152312 267936 152364
rect 274876 152312 274928 152364
rect 368532 152312 368584 152364
rect 368716 152312 368768 152364
rect 85908 151360 85960 151412
rect 87472 151360 87524 151412
rect 320784 151360 320836 151412
rect 323268 151360 323320 151412
rect 225564 150952 225616 151004
rect 226208 150952 226260 151004
rect 173676 150884 173728 150936
rect 182324 150884 182376 150936
rect 225656 150884 225708 150936
rect 233476 150884 233528 150936
rect 267700 150884 267752 150936
rect 274876 150884 274928 150936
rect 323176 150884 323228 150936
rect 328420 150884 328472 150936
rect 177540 150816 177592 150868
rect 182232 150816 182284 150868
rect 225564 150816 225616 150868
rect 231360 150816 231412 150868
rect 266596 150816 266648 150868
rect 271380 150816 271432 150868
rect 174044 150748 174096 150800
rect 181036 150748 181088 150800
rect 181036 150612 181088 150664
rect 181680 150612 181732 150664
rect 77260 149796 77312 149848
rect 85816 149796 85868 149848
rect 321612 149728 321664 149780
rect 327224 149728 327276 149780
rect 80112 149592 80164 149644
rect 87196 149592 87248 149644
rect 321060 149592 321112 149644
rect 323176 149592 323228 149644
rect 131816 149524 131868 149576
rect 139636 149524 139688 149576
rect 176252 149524 176304 149576
rect 182324 149524 182376 149576
rect 323268 149524 323320 149576
rect 328420 149524 328472 149576
rect 131356 149456 131408 149508
rect 137612 149456 137664 149508
rect 174044 149456 174096 149508
rect 178920 149456 178972 149508
rect 225288 149388 225340 149440
rect 227220 149388 227272 149440
rect 266596 149388 266648 149440
rect 275704 149388 275756 149440
rect 12860 149320 12912 149372
rect 16264 149320 16316 149372
rect 225196 148640 225248 148692
rect 227312 148640 227364 148692
rect 78916 148436 78968 148488
rect 85908 148436 85960 148488
rect 321612 148368 321664 148420
rect 327868 148368 327920 148420
rect 174044 148164 174096 148216
rect 180300 148164 180352 148216
rect 228784 148164 228836 148216
rect 233476 148164 233528 148216
rect 266596 148164 266648 148216
rect 274140 148164 274192 148216
rect 323176 148164 323228 148216
rect 328420 148164 328472 148216
rect 78916 147688 78968 147740
rect 87012 147688 87064 147740
rect 132276 146736 132328 146788
rect 140556 146736 140608 146788
rect 226300 146736 226352 146788
rect 233476 146736 233528 146788
rect 267884 146736 267936 146788
rect 275520 146736 275572 146788
rect 79376 145376 79428 145428
rect 87196 145376 87248 145428
rect 91704 145376 91756 145428
rect 128136 145376 128188 145428
rect 132460 145376 132512 145428
rect 140556 145376 140608 145428
rect 185636 145376 185688 145428
rect 222160 145376 222212 145428
rect 226392 145376 226444 145428
rect 233476 145376 233528 145428
rect 266780 145376 266832 145428
rect 275612 145376 275664 145428
rect 279660 145376 279712 145428
rect 322808 145376 322860 145428
rect 116084 144832 116136 144884
rect 128044 144832 128096 144884
rect 292724 144832 292776 144884
rect 312320 144832 312372 144884
rect 103664 144764 103716 144816
rect 124272 144764 124324 144816
rect 171284 144764 171336 144816
rect 189224 144764 189276 144816
rect 197504 144764 197556 144816
rect 218296 144764 218348 144816
rect 280304 144764 280356 144816
rect 308732 144764 308784 144816
rect 91244 144696 91296 144748
rect 120684 144696 120736 144748
rect 185084 144696 185136 144748
rect 214708 144696 214760 144748
rect 218940 144696 218992 144748
rect 221976 144696 222028 144748
rect 290516 144696 290568 144748
rect 326580 144696 326632 144748
rect 312780 144084 312832 144136
rect 316000 144084 316052 144136
rect 132368 144016 132420 144068
rect 140556 144016 140608 144068
rect 226484 144016 226536 144068
rect 233476 144016 233528 144068
rect 321796 144016 321848 144068
rect 327316 144016 327368 144068
rect 95292 143880 95344 143932
rect 211028 143404 211080 143456
rect 231360 143404 231412 143456
rect 76892 143336 76944 143388
rect 88576 143336 88628 143388
rect 203760 143336 203812 143388
rect 231176 143336 231228 143388
rect 294288 143336 294340 143388
rect 325292 143336 325344 143388
rect 78916 143200 78968 143252
rect 87104 143200 87156 143252
rect 200172 142248 200224 142300
rect 167972 142180 168024 142232
rect 168524 142180 168576 142232
rect 196860 142180 196912 142232
rect 236880 142180 236932 142232
rect 238996 142180 239048 142232
rect 239916 142180 239968 142232
rect 261904 142180 261956 142232
rect 76064 142087 76116 142096
rect 76064 142053 76073 142087
rect 76073 142053 76107 142087
rect 76107 142053 76116 142087
rect 76064 142044 76116 142053
rect 305052 142044 305104 142096
rect 324556 142044 324608 142096
rect 127584 141976 127636 142028
rect 140372 141976 140424 142028
rect 173584 141976 173636 142028
rect 219676 141976 219728 142028
rect 233476 141976 233528 142028
rect 267332 141976 267384 142028
rect 316276 141976 316328 142028
rect 136876 141364 136928 141416
rect 150400 141364 150452 141416
rect 167972 141364 168024 141416
rect 78916 141296 78968 141348
rect 127216 141296 127268 141348
rect 127584 141296 127636 141348
rect 147456 141296 147508 141348
rect 171284 141296 171336 141348
rect 231360 141296 231412 141348
rect 246908 141296 246960 141348
rect 261904 141296 261956 141348
rect 316276 141296 316328 141348
rect 327316 141296 327368 141348
rect 74132 141228 74184 141280
rect 75420 141228 75472 141280
rect 113416 141228 113468 141280
rect 113876 141228 113928 141280
rect 231176 141228 231228 141280
rect 231452 141228 231504 141280
rect 427320 140752 427372 140804
rect 429528 140752 429580 140804
rect 113876 140616 113928 140668
rect 137244 140616 137296 140668
rect 73948 140548 74000 140600
rect 102376 140548 102428 140600
rect 137336 140548 137388 140600
rect 207256 140548 207308 140600
rect 231084 140548 231136 140600
rect 301096 140548 301148 140600
rect 325108 140548 325160 140600
rect 76064 140183 76116 140192
rect 76064 140149 76073 140183
rect 76073 140149 76107 140183
rect 76107 140149 76116 140183
rect 76064 140140 76116 140149
rect 164568 139868 164620 139920
rect 251140 139868 251192 139920
rect 253992 139868 254044 139920
rect 150584 139800 150636 139852
rect 162268 139800 162320 139852
rect 239548 139800 239600 139852
rect 322716 139800 322768 139852
rect 64840 139732 64892 139784
rect 70452 139732 70504 139784
rect 156104 139732 156156 139784
rect 157576 139732 157628 139784
rect 63644 139664 63696 139716
rect 75236 139664 75288 139716
rect 151780 139664 151832 139716
rect 157484 139664 157536 139716
rect 169996 139732 170048 139784
rect 241756 139732 241808 139784
rect 244976 139732 245028 139784
rect 247092 139732 247144 139784
rect 259236 139732 259288 139784
rect 160060 139664 160112 139716
rect 162636 139664 162688 139716
rect 169076 139664 169128 139716
rect 244332 139664 244384 139716
rect 256292 139664 256344 139716
rect 62264 139596 62316 139648
rect 74224 139596 74276 139648
rect 156104 139596 156156 139648
rect 249208 139596 249260 139648
rect 252060 139596 252112 139648
rect 60884 139528 60936 139580
rect 73120 139528 73172 139580
rect 154264 139528 154316 139580
rect 157300 139528 157352 139580
rect 158864 139528 158916 139580
rect 160980 139528 161032 139580
rect 161992 139528 162044 139580
rect 163004 139528 163056 139580
rect 241480 139528 241532 139580
rect 249668 139528 249720 139580
rect 249852 139528 249904 139580
rect 253072 139528 253124 139580
rect 59504 139460 59556 139512
rect 71096 139460 71148 139512
rect 56744 139392 56796 139444
rect 67968 139392 68020 139444
rect 116176 139460 116228 139512
rect 154724 139460 154776 139512
rect 167328 139460 167380 139512
rect 151872 139392 151924 139444
rect 158128 139392 158180 139444
rect 160796 139392 160848 139444
rect 160888 139392 160940 139444
rect 163464 139392 163516 139444
rect 251324 139392 251376 139444
rect 264112 139596 264164 139648
rect 58124 139324 58176 139376
rect 70084 139324 70136 139376
rect 75144 139324 75196 139376
rect 55364 139256 55416 139308
rect 66956 139256 67008 139308
rect 150492 139324 150544 139376
rect 163280 139324 163332 139376
rect 249944 139324 249996 139376
rect 263100 139528 263152 139580
rect 261260 139460 261312 139512
rect 260156 139392 260208 139444
rect 258316 139324 258368 139376
rect 154632 139256 154684 139308
rect 168064 139256 168116 139308
rect 244424 139256 244476 139308
rect 257304 139256 257356 139308
rect 60792 139188 60844 139240
rect 72108 139188 72160 139240
rect 144604 139188 144656 139240
rect 170732 139188 170784 139240
rect 238628 139188 238680 139240
rect 264480 139188 264532 139240
rect 333388 139188 333440 139240
rect 334124 139188 334176 139240
rect 152700 139120 152752 139172
rect 153344 139120 153396 139172
rect 63828 139052 63880 139104
rect 68612 139052 68664 139104
rect 136876 138984 136928 139036
rect 165212 139120 165264 139172
rect 249852 139120 249904 139172
rect 262088 139120 262140 139172
rect 248564 139052 248616 139104
rect 166132 138984 166184 139036
rect 247184 138984 247236 139036
rect 58676 138916 58728 138968
rect 63000 138916 63052 138968
rect 64380 138916 64432 138968
rect 68980 138916 69032 138968
rect 157576 138916 157628 138968
rect 158220 138916 158272 138968
rect 245804 138916 245856 138968
rect 62816 138848 62868 138900
rect 67692 138848 67744 138900
rect 157116 138848 157168 138900
rect 159968 138848 160020 138900
rect 244976 138848 245028 138900
rect 252244 138848 252296 138900
rect 341760 138848 341812 138900
rect 59688 138780 59740 138832
rect 63092 138780 63144 138832
rect 242492 138780 242544 138832
rect 249116 138780 249168 138832
rect 253900 138780 253952 138832
rect 256660 138780 256712 138832
rect 338264 138780 338316 138832
rect 342680 138780 342732 138832
rect 345808 138780 345860 138832
rect 61804 138712 61856 138764
rect 65760 138712 65812 138764
rect 145248 138712 145300 138764
rect 365220 138712 365272 138764
rect 60700 138644 60752 138696
rect 63184 138644 63236 138696
rect 252152 138644 252204 138696
rect 254176 138644 254228 138696
rect 256016 138644 256068 138696
rect 258684 138644 258736 138696
rect 338172 138644 338224 138696
rect 341668 138644 341720 138696
rect 341944 138644 341996 138696
rect 344796 138644 344848 138696
rect 57664 138576 57716 138628
rect 61620 138576 61672 138628
rect 65944 138576 65996 138628
rect 70544 138576 70596 138628
rect 155184 138576 155236 138628
rect 158036 138576 158088 138628
rect 252704 138576 252756 138628
rect 254820 138576 254872 138628
rect 255004 138576 255056 138628
rect 257488 138576 257540 138628
rect 334400 138576 334452 138628
rect 335504 138576 335556 138628
rect 338540 138576 338592 138628
rect 339644 138576 339696 138628
rect 341852 138576 341904 138628
rect 343784 138576 343836 138628
rect 348660 138576 348712 138628
rect 349948 138576 350000 138628
rect 284444 137828 284496 137880
rect 324832 137828 324884 137880
rect 12860 137080 12912 137132
rect 16080 137080 16132 137132
rect 137152 137080 137204 137132
rect 137428 137080 137480 137132
rect 210016 136672 210068 136724
rect 218940 136672 218992 136724
rect 346636 136468 346688 136520
rect 347556 136468 347608 136520
rect 304040 136400 304092 136452
rect 312780 136400 312832 136452
rect 291528 136264 291580 136316
rect 292724 136264 292776 136316
rect 279108 136128 279160 136180
rect 280304 136128 280356 136180
rect 324556 135788 324608 135840
rect 347004 135788 347056 135840
rect 359056 135720 359108 135772
rect 286744 135040 286796 135092
rect 324648 135040 324700 135092
rect 343876 135040 343928 135092
rect 360804 135040 360856 135092
rect 324648 134428 324700 134480
rect 343876 134428 343928 134480
rect 51500 134360 51552 134412
rect 51592 134360 51644 134412
rect 343968 133680 344020 133732
rect 360712 133680 360764 133732
rect 326580 133000 326632 133052
rect 343968 133000 344020 133052
rect 344244 133000 344296 133052
rect 346084 132456 346136 132508
rect 360436 132456 360488 132508
rect 354916 132388 354968 132440
rect 355836 132388 355888 132440
rect 136876 132320 136928 132372
rect 137336 132320 137388 132372
rect 343324 132320 343376 132372
rect 360988 132320 361040 132372
rect 258960 132252 259012 132304
rect 368900 132252 368952 132304
rect 324556 132184 324608 132236
rect 324740 132184 324792 132236
rect 324832 131708 324884 131760
rect 325476 131708 325528 131760
rect 343324 131708 343376 131760
rect 325108 131640 325160 131692
rect 346084 131640 346136 131692
rect 56100 131572 56152 131624
rect 56744 131572 56796 131624
rect 59688 131572 59740 131624
rect 60792 131572 60844 131624
rect 155460 131572 155512 131624
rect 156104 131572 156156 131624
rect 245344 131572 245396 131624
rect 245804 131572 245856 131624
rect 248012 131572 248064 131624
rect 248564 131572 248616 131624
rect 341668 131572 341720 131624
rect 348016 131572 348068 131624
rect 339644 131504 339696 131556
rect 350960 131504 351012 131556
rect 160980 131436 161032 131488
rect 161716 131436 161768 131488
rect 341024 131436 341076 131488
rect 352248 131436 352300 131488
rect 339552 131368 339604 131420
rect 351604 131368 351656 131420
rect 338080 131300 338132 131352
rect 350408 131300 350460 131352
rect 231360 131232 231412 131284
rect 322624 131232 322676 131284
rect 335504 131232 335556 131284
rect 348568 131232 348620 131284
rect 248472 131164 248524 131216
rect 250956 131164 251008 131216
rect 336884 131164 336936 131216
rect 349764 131164 349816 131216
rect 332744 131096 332796 131148
rect 341024 131096 341076 131148
rect 346636 131096 346688 131148
rect 334124 131028 334176 131080
rect 348016 131028 348068 131080
rect 335412 130960 335464 131012
rect 349396 130960 349448 131012
rect 340564 130892 340616 130944
rect 346728 130892 346780 130944
rect 63184 130688 63236 130740
rect 65944 130688 65996 130740
rect 243596 130688 243648 130740
rect 244332 130688 244384 130740
rect 250680 130688 250732 130740
rect 251324 130688 251376 130740
rect 57020 130552 57072 130604
rect 64380 130552 64432 130604
rect 63092 130484 63144 130536
rect 65024 130484 65076 130536
rect 61620 130416 61672 130468
rect 63276 130416 63328 130468
rect 246264 130416 246316 130468
rect 247092 130416 247144 130468
rect 248932 130416 248984 130468
rect 249852 130416 249904 130468
rect 325384 130416 325436 130468
rect 342496 130824 342548 130876
rect 342404 130756 342456 130808
rect 348660 130756 348712 130808
rect 347280 130688 347332 130740
rect 62356 130348 62408 130400
rect 63644 130348 63696 130400
rect 324740 130348 324792 130400
rect 325292 130348 325344 130400
rect 338724 130552 338776 130604
rect 341852 130552 341904 130604
rect 339368 130484 339420 130536
rect 341944 130484 341996 130536
rect 345164 130484 345216 130536
rect 360896 130892 360948 130944
rect 360344 130416 360396 130468
rect 360528 130416 360580 130468
rect 337528 130348 337580 130400
rect 338172 130348 338224 130400
rect 339552 130348 339604 130400
rect 341760 130348 341812 130400
rect 61436 130280 61488 130332
rect 62264 130280 62316 130332
rect 63000 130280 63052 130332
rect 64104 130280 64156 130332
rect 65760 130280 65812 130332
rect 66772 130280 66824 130332
rect 149296 130280 149348 130332
rect 150584 130280 150636 130332
rect 151044 130280 151096 130332
rect 151780 130280 151832 130332
rect 153712 130280 153764 130332
rect 154724 130280 154776 130332
rect 156380 130280 156432 130332
rect 157484 130280 157536 130332
rect 158220 130280 158272 130332
rect 159048 130280 159100 130332
rect 163004 130280 163056 130332
rect 164384 130280 164436 130332
rect 254820 130280 254872 130332
rect 255556 130280 255608 130332
rect 324648 130280 324700 130332
rect 345716 130280 345768 130332
rect 361080 130280 361132 130332
rect 231084 130212 231136 130264
rect 246448 130212 246500 130264
rect 137060 127492 137112 127544
rect 137428 127492 137480 127544
rect 84712 127424 84764 127476
rect 85816 127424 85868 127476
rect 38804 126744 38856 126796
rect 48464 126744 48516 126796
rect 357676 126744 357728 126796
rect 405976 126744 406028 126796
rect 38252 126064 38304 126116
rect 52604 126064 52656 126116
rect 356204 126064 356256 126116
rect 405976 126064 406028 126116
rect 76892 125452 76944 125504
rect 82688 125452 82740 125504
rect 169996 125384 170048 125436
rect 170732 125384 170784 125436
rect 175516 125384 175568 125436
rect 263836 125248 263888 125300
rect 264480 125248 264532 125300
rect 270368 125248 270420 125300
rect 76156 125044 76208 125096
rect 76892 125044 76944 125096
rect 12676 123276 12728 123328
rect 16172 123276 16224 123328
rect 38804 122596 38856 122648
rect 54076 122596 54128 122648
rect 356296 122596 356348 122648
rect 405976 122596 406028 122648
rect 137612 121984 137664 122036
rect 144236 121984 144288 122036
rect 231452 121984 231504 122036
rect 240376 121984 240428 122036
rect 325292 121984 325344 122036
rect 334216 121984 334268 122036
rect 38804 120556 38856 120608
rect 52604 120556 52656 120608
rect 356204 120556 356256 120608
rect 405976 120556 406028 120608
rect 324556 119876 324608 119928
rect 326580 119876 326632 119928
rect 262364 117904 262416 117956
rect 270000 117904 270052 117956
rect 167880 117836 167932 117888
rect 176252 117836 176304 117888
rect 38252 117088 38304 117140
rect 54076 117088 54128 117140
rect 354916 117088 354968 117140
rect 405976 117088 406028 117140
rect 427412 116408 427464 116460
rect 429436 116408 429488 116460
rect 51684 115116 51736 115168
rect 38804 115048 38856 115100
rect 52144 115048 52196 115100
rect 356204 115048 356256 115100
rect 405976 115048 406028 115100
rect 51592 113731 51644 113740
rect 51592 113697 51601 113731
rect 51601 113697 51635 113731
rect 51635 113697 51644 113731
rect 51592 113688 51644 113697
rect 38804 112940 38856 112992
rect 51868 112940 51920 112992
rect 136876 112940 136928 112992
rect 146628 112940 146680 112992
rect 355008 112940 355060 112992
rect 405976 112940 406028 112992
rect 38252 110900 38304 110952
rect 52604 110968 52656 111020
rect 427596 110968 427648 111020
rect 428792 110968 428844 111020
rect 136876 110900 136928 110952
rect 145340 110900 145392 110952
rect 356204 110900 356256 110952
rect 406068 110900 406120 110952
rect 84712 109744 84764 109796
rect 85816 109744 85868 109796
rect 232004 109540 232056 109592
rect 238996 109540 239048 109592
rect 240100 109540 240152 109592
rect 74316 109472 74368 109524
rect 82596 109472 82648 109524
rect 51592 108248 51644 108300
rect 137704 108180 137756 108232
rect 143960 108180 144012 108232
rect 231544 108180 231596 108232
rect 240836 108180 240888 108232
rect 325384 108180 325436 108232
rect 334216 108180 334268 108232
rect 358320 108180 358372 108232
rect 358320 108044 358372 108096
rect 38804 107432 38856 107484
rect 353536 107432 353588 107484
rect 405976 107432 406028 107484
rect 13320 105460 13372 105512
rect 18104 105460 18156 105512
rect 427596 105460 427648 105512
rect 430080 105460 430132 105512
rect 38804 105392 38856 105444
rect 52604 105392 52656 105444
rect 356204 105392 356256 105444
rect 405976 105392 406028 105444
rect 358320 105367 358372 105376
rect 358320 105333 358329 105367
rect 358329 105333 358363 105367
rect 358363 105333 358372 105367
rect 358320 105324 358372 105333
rect 51684 104075 51736 104084
rect 51684 104041 51693 104075
rect 51693 104041 51727 104075
rect 51727 104041 51736 104075
rect 51684 104032 51736 104041
rect 427596 102672 427648 102724
rect 429436 102672 429488 102724
rect 352708 101924 352760 101976
rect 405976 101924 406028 101976
rect 50028 101516 50080 101568
rect 51316 101516 51368 101568
rect 38620 101312 38672 101364
rect 50028 101312 50080 101364
rect 38804 100564 38856 100616
rect 52604 100564 52656 100616
rect 356204 100564 356256 100616
rect 405976 100564 406028 100616
rect 13504 99884 13556 99936
rect 17460 99884 17512 99936
rect 167880 98524 167932 98576
rect 173400 98524 173452 98576
rect 261168 98524 261220 98576
rect 267240 98524 267292 98576
rect 38804 97776 38856 97828
rect 49936 97776 49988 97828
rect 352800 97776 352852 97828
rect 405976 97776 406028 97828
rect 13136 95804 13188 95856
rect 18104 95804 18156 95856
rect 38068 95736 38120 95788
rect 52604 95804 52656 95856
rect 358320 95847 358372 95856
rect 358320 95813 358329 95847
rect 358329 95813 358363 95847
rect 358363 95813 358372 95847
rect 358320 95804 358372 95813
rect 427228 95804 427280 95856
rect 430172 95804 430224 95856
rect 356204 95736 356256 95788
rect 405976 95736 406028 95788
rect 324556 95056 324608 95108
rect 330076 95056 330128 95108
rect 232004 94988 232056 95040
rect 236236 94988 236288 95040
rect 138164 94376 138216 94428
rect 142396 94376 142448 94428
rect 235500 94376 235552 94428
rect 240376 94376 240428 94428
rect 329340 94376 329392 94428
rect 334216 94376 334268 94428
rect 73396 93696 73448 93748
rect 73672 93696 73724 93748
rect 84804 93424 84856 93476
rect 85816 93424 85868 93476
rect 267240 92948 267292 93000
rect 270368 92948 270420 93000
rect 75420 92676 75472 92728
rect 82688 92676 82740 92728
rect 173400 92540 173452 92592
rect 175516 92540 175568 92592
rect 37608 92268 37660 92320
rect 48556 92268 48608 92320
rect 352800 92268 352852 92320
rect 405976 92268 406028 92320
rect 13412 91588 13464 91640
rect 18104 91588 18156 91640
rect 73396 91452 73448 91504
rect 76800 91452 76852 91504
rect 38804 90160 38856 90212
rect 52604 90160 52656 90212
rect 356204 90160 356256 90212
rect 405976 90160 406028 90212
rect 51684 89004 51736 89056
rect 358320 88868 358372 88920
rect 358412 88664 358464 88716
rect 23900 87440 23952 87492
rect 72016 87440 72068 87492
rect 150400 87440 150452 87492
rect 154080 87440 154132 87492
rect 154724 87440 154776 87492
rect 172020 87440 172072 87492
rect 361080 87440 361132 87492
rect 418212 87440 418264 87492
rect 36044 87372 36096 87424
rect 73856 87372 73908 87424
rect 160980 87372 161032 87424
rect 163924 87372 163976 87424
rect 249024 87372 249076 87424
rect 258960 87372 259012 87424
rect 359700 87372 359752 87424
rect 360344 87372 360396 87424
rect 415544 87372 415596 87424
rect 29236 87304 29288 87356
rect 73580 87304 73632 87356
rect 149756 87304 149808 87356
rect 154172 87304 154224 87356
rect 343508 87304 343560 87356
rect 348200 87304 348252 87356
rect 370004 87304 370056 87356
rect 410208 87304 410260 87356
rect 31904 87236 31956 87288
rect 73488 87236 73540 87288
rect 151044 87236 151096 87288
rect 155460 87236 155512 87288
rect 244424 87236 244476 87288
rect 254176 87236 254228 87288
rect 340932 87236 340984 87288
rect 345256 87236 345308 87288
rect 34572 87168 34624 87220
rect 73672 87168 73724 87220
rect 336884 87168 336936 87220
rect 348752 87168 348804 87220
rect 21232 87100 21284 87152
rect 34664 87100 34716 87152
rect 64380 87100 64432 87152
rect 65944 87100 65996 87152
rect 149204 87100 149256 87152
rect 157576 87100 157628 87152
rect 243044 87100 243096 87152
rect 255096 87100 255148 87152
rect 338080 87100 338132 87152
rect 349580 87100 349632 87152
rect 26568 87032 26620 87084
rect 36044 87032 36096 87084
rect 150584 87032 150636 87084
rect 162084 87032 162136 87084
rect 339644 87032 339696 87084
rect 351236 87032 351288 87084
rect 59688 86964 59740 87016
rect 67140 86964 67192 87016
rect 149204 86964 149256 87016
rect 161440 86964 161492 87016
rect 241664 86964 241716 87016
rect 254544 86964 254596 87016
rect 334124 86964 334176 87016
rect 146444 86896 146496 86948
rect 160244 86896 160296 86948
rect 244056 86896 244108 86948
rect 252980 86896 253032 86948
rect 335412 86896 335464 86948
rect 341024 86964 341076 87016
rect 352156 86964 352208 87016
rect 346176 86896 346228 86948
rect 57020 86828 57072 86880
rect 67876 86828 67928 86880
rect 147824 86828 147876 86880
rect 160888 86828 160940 86880
rect 240284 86828 240336 86880
rect 254268 86828 254320 86880
rect 335504 86828 335556 86880
rect 348016 86828 348068 86880
rect 56100 86760 56152 86812
rect 66680 86760 66732 86812
rect 145064 86760 145116 86812
rect 159600 86760 159652 86812
rect 238904 86760 238956 86812
rect 253440 86760 253492 86812
rect 332744 86760 332796 86812
rect 345348 86760 345400 86812
rect 347004 86692 347056 86744
rect 344336 86624 344388 86676
rect 347280 86624 347332 86676
rect 257580 86488 257632 86540
rect 258408 86488 258460 86540
rect 345072 86488 345124 86540
rect 362460 86488 362512 86540
rect 252152 86216 252204 86268
rect 255740 86216 255792 86268
rect 61620 86148 61672 86200
rect 63276 86148 63328 86200
rect 67232 86148 67284 86200
rect 68612 86148 68664 86200
rect 162360 86148 162412 86200
rect 164568 86148 164620 86200
rect 245344 86148 245396 86200
rect 252060 86148 252112 86200
rect 51500 86123 51552 86132
rect 51500 86089 51509 86123
rect 51509 86089 51543 86123
rect 51543 86089 51552 86123
rect 51500 86080 51552 86089
rect 61436 86080 61488 86132
rect 62264 86080 62316 86132
rect 62356 86080 62408 86132
rect 63644 86080 63696 86132
rect 63736 86080 63788 86132
rect 64748 86080 64800 86132
rect 65760 86080 65812 86132
rect 66772 86080 66824 86132
rect 68520 86080 68572 86132
rect 69440 86080 69492 86132
rect 152240 86080 152292 86132
rect 153252 86080 153304 86132
rect 153436 86080 153488 86132
rect 154724 86080 154776 86132
rect 162452 86080 162504 86132
rect 163280 86080 163332 86132
rect 243504 86080 243556 86132
rect 245160 86080 245212 86132
rect 246540 86080 246592 86132
rect 247092 86080 247144 86132
rect 247736 86080 247788 86132
rect 248564 86080 248616 86132
rect 257672 86148 257724 86200
rect 337620 86148 337672 86200
rect 339092 86148 339144 86200
rect 341668 86148 341720 86200
rect 344612 86148 344664 86200
rect 256292 86080 256344 86132
rect 256936 86080 256988 86132
rect 338264 86080 338316 86132
rect 339000 86080 339052 86132
rect 340104 86080 340156 86132
rect 341760 86080 341812 86132
rect 342404 86080 342456 86132
rect 344520 86080 344572 86132
rect 345900 86080 345952 86132
rect 350408 86080 350460 86132
rect 66588 86012 66640 86064
rect 67324 86012 67376 86064
rect 137888 86012 137940 86064
rect 145800 86012 145852 86064
rect 256200 86012 256252 86064
rect 324556 86012 324608 86064
rect 329340 86012 329392 86064
rect 358412 86055 358464 86064
rect 358412 86021 358421 86055
rect 358421 86021 358455 86055
rect 358455 86021 358464 86055
rect 358412 86012 358464 86021
rect 231084 85740 231136 85792
rect 235500 85740 235552 85792
rect 354916 84040 354968 84092
rect 355836 84040 355888 84092
rect 88484 81932 88536 81984
rect 178736 81932 178788 81984
rect 182416 81932 182468 81984
rect 276348 81932 276400 81984
rect 95752 81864 95804 81916
rect 170640 81864 170692 81916
rect 189500 81864 189552 81916
rect 283156 81864 283208 81916
rect 102928 81796 102980 81848
rect 176160 81796 176212 81848
rect 196676 81796 196728 81848
rect 290332 81796 290384 81848
rect 285824 81320 285876 81372
rect 297508 81320 297560 81372
rect 96764 81252 96816 81304
rect 109828 81252 109880 81304
rect 190604 81252 190656 81304
rect 203760 81252 203812 81304
rect 276348 81252 276400 81304
rect 428056 81252 428108 81304
rect 224460 80572 224512 80624
rect 225196 80572 225248 80624
rect 318300 80572 318352 80624
rect 319128 80572 319180 80624
rect 236236 79348 236288 79400
rect 237248 79348 237300 79400
rect 60240 79144 60292 79196
rect 64380 79144 64432 79196
rect 66588 79144 66640 79196
rect 75788 79144 75840 79196
rect 76892 79144 76944 79196
rect 155460 79144 155512 79196
rect 161716 79144 161768 79196
rect 245160 79144 245212 79196
rect 251416 79144 251468 79196
rect 252060 79144 252112 79196
rect 255556 79144 255608 79196
rect 333388 79144 333440 79196
rect 334124 79144 334176 79196
rect 334400 79144 334452 79196
rect 335412 79144 335464 79196
rect 339552 79144 339604 79196
rect 343784 79144 343836 79196
rect 344520 79144 344572 79196
rect 65484 79076 65536 79128
rect 69348 79076 69400 79128
rect 154172 79076 154224 79128
rect 158956 79076 159008 79128
rect 249024 79076 249076 79128
rect 256200 79076 256252 79128
rect 339000 79076 339052 79128
rect 342680 79076 342732 79128
rect 344612 79076 344664 79128
rect 346820 79076 346872 79128
rect 347280 79144 347332 79196
rect 349948 79144 350000 79196
rect 347924 79076 347976 79128
rect 57204 79008 57256 79060
rect 61620 79008 61672 79060
rect 154724 79008 154776 79060
rect 160980 79008 161032 79060
rect 337528 79008 337580 79060
rect 338264 79008 338316 79060
rect 341760 79008 341812 79060
rect 344796 79008 344848 79060
rect 62356 78940 62408 78992
rect 58124 78872 58176 78924
rect 64380 78872 64432 78924
rect 68520 78872 68572 78924
rect 63644 78804 63696 78856
rect 74776 78804 74828 78856
rect 62264 78736 62316 78788
rect 67140 78736 67192 78788
rect 71648 78736 71700 78788
rect 151964 78940 152016 78992
rect 154080 78940 154132 78992
rect 160336 78940 160388 78992
rect 244884 78940 244936 78992
rect 252152 78940 252204 78992
rect 153344 78872 153396 78924
rect 162452 78872 162504 78924
rect 247644 78872 247696 78924
rect 256292 78872 256344 78924
rect 151964 78804 152016 78856
rect 161808 78804 161860 78856
rect 246264 78804 246316 78856
rect 255648 78804 255700 78856
rect 163096 78736 163148 78788
rect 245804 78736 245856 78788
rect 256936 78736 256988 78788
rect 60884 78668 60936 78720
rect 72660 78668 72712 78720
rect 153252 78668 153304 78720
rect 164568 78668 164620 78720
rect 247092 78668 247144 78720
rect 258408 78668 258460 78720
rect 339092 78668 339144 78720
rect 341668 78668 341720 78720
rect 59228 78600 59280 78652
rect 63736 78600 63788 78652
rect 59504 78532 59556 78584
rect 70636 78600 70688 78652
rect 153436 78600 153488 78652
rect 165948 78600 166000 78652
rect 248564 78600 248616 78652
rect 261076 78600 261128 78652
rect 338540 78600 338592 78652
rect 345900 78600 345952 78652
rect 69624 78532 69676 78584
rect 154632 78532 154684 78584
rect 167328 78532 167380 78584
rect 247184 78532 247236 78584
rect 259696 78532 259748 78584
rect 55364 78464 55416 78516
rect 66496 78464 66548 78516
rect 73764 78464 73816 78516
rect 154448 78464 154500 78516
rect 168708 78464 168760 78516
rect 248472 78464 248524 78516
rect 262456 78464 262508 78516
rect 63368 78396 63420 78448
rect 67232 78396 67284 78448
rect 58216 78328 58268 78380
rect 63828 78328 63880 78380
rect 156104 78328 156156 78380
rect 162360 78328 162412 78380
rect 250404 78328 250456 78380
rect 257580 78328 257632 78380
rect 61344 78056 61396 78108
rect 65760 78056 65812 78108
rect 427412 77784 427464 77836
rect 429528 77784 429580 77836
rect 88024 76424 88076 76476
rect 88208 76424 88260 76476
rect 358504 76424 358556 76476
rect 79468 76356 79520 76408
rect 123996 76356 124048 76408
rect 139636 76356 139688 76408
rect 173860 76356 173912 76408
rect 218020 76356 218072 76408
rect 233476 76356 233528 76408
rect 266596 76356 266648 76408
rect 312044 76356 312096 76408
rect 328420 76356 328472 76408
rect 80204 73704 80256 73756
rect 87932 73704 87984 73756
rect 174044 73704 174096 73756
rect 181036 73704 181088 73756
rect 226576 73704 226628 73756
rect 233476 73704 233528 73756
rect 266596 73704 266648 73756
rect 274876 73704 274928 73756
rect 304868 73704 304920 73756
rect 305052 73704 305104 73756
rect 321796 73704 321848 73756
rect 328328 73704 328380 73756
rect 110196 73432 110248 73484
rect 116820 73432 116872 73484
rect 204128 72956 204180 73008
rect 210936 72956 210988 73008
rect 217560 72956 217612 73008
rect 224460 72956 224512 73008
rect 311216 72616 311268 72668
rect 318300 72616 318352 72668
rect 79836 72344 79888 72396
rect 85724 72344 85776 72396
rect 123536 72344 123588 72396
rect 130988 72344 131040 72396
rect 172940 72344 172992 72396
rect 180944 72344 180996 72396
rect 230164 72344 230216 72396
rect 233476 72344 233528 72396
rect 266596 72344 266648 72396
rect 274692 72344 274744 72396
rect 284536 72344 284588 72396
rect 285824 72344 285876 72396
rect 297876 72344 297928 72396
rect 304868 72344 304920 72396
rect 78916 70984 78968 71036
rect 85632 70984 85684 71036
rect 174044 70984 174096 71036
rect 178460 70984 178512 71036
rect 266596 70984 266648 71036
rect 272024 70984 272076 71036
rect 132552 70916 132604 70968
rect 139636 70916 139688 70968
rect 173308 70916 173360 70968
rect 178276 70916 178328 70968
rect 230624 70916 230676 70968
rect 233568 70916 233620 70968
rect 266688 70916 266740 70968
rect 274784 70916 274836 70968
rect 321244 70916 321296 70968
rect 328512 70916 328564 70968
rect 174044 69896 174096 69948
rect 178368 69896 178420 69948
rect 80204 69556 80256 69608
rect 87288 69556 87340 69608
rect 266596 69556 266648 69608
rect 274968 69556 275020 69608
rect 358504 69624 358556 69676
rect 131356 69488 131408 69540
rect 139728 69488 139780 69540
rect 225932 69488 225984 69540
rect 230164 69488 230216 69540
rect 358412 69488 358464 69540
rect 131816 69420 131868 69472
rect 139544 69420 139596 69472
rect 321612 69080 321664 69132
rect 327224 69080 327276 69132
rect 85724 68944 85776 68996
rect 87656 68944 87708 68996
rect 79284 68196 79336 68248
rect 85080 68196 85132 68248
rect 136784 68196 136836 68248
rect 139636 68196 139688 68248
rect 172940 68196 172992 68248
rect 180944 68196 180996 68248
rect 266596 68196 266648 68248
rect 274692 68196 274744 68248
rect 85632 68128 85684 68180
rect 87840 68128 87892 68180
rect 132368 68128 132420 68180
rect 139912 68128 139964 68180
rect 178276 68128 178328 68180
rect 181404 68128 181456 68180
rect 226300 68128 226352 68180
rect 233476 68128 233528 68180
rect 79560 67516 79612 67568
rect 129424 67516 129476 67568
rect 173400 67516 173452 67568
rect 223448 67516 223500 67568
rect 267240 67516 267292 67568
rect 317564 67516 317616 67568
rect 80204 67176 80256 67228
rect 82780 67176 82832 67228
rect 321612 67040 321664 67092
rect 327040 67040 327092 67092
rect 174044 66904 174096 66956
rect 179104 66904 179156 66956
rect 135956 66836 136008 66888
rect 139728 66836 139780 66888
rect 266688 66836 266740 66888
rect 272668 66836 272720 66888
rect 80204 66768 80256 66820
rect 87380 66768 87432 66820
rect 136140 66768 136192 66820
rect 139636 66768 139688 66820
rect 173860 66768 173912 66820
rect 181772 66768 181824 66820
rect 266596 66768 266648 66820
rect 274232 66768 274284 66820
rect 80296 66700 80348 66752
rect 87196 66700 87248 66752
rect 88208 66743 88260 66752
rect 88208 66709 88217 66743
rect 88217 66709 88251 66743
rect 88251 66709 88260 66743
rect 88208 66700 88260 66709
rect 132368 66700 132420 66752
rect 139820 66700 139872 66752
rect 226392 66700 226444 66752
rect 233568 66700 233620 66752
rect 272024 66700 272076 66752
rect 274876 66700 274928 66752
rect 317380 66700 317432 66752
rect 226300 66632 226352 66684
rect 230624 66632 230676 66684
rect 178368 66428 178420 66480
rect 182140 66428 182192 66480
rect 178460 66156 178512 66208
rect 181956 66156 182008 66208
rect 321612 65952 321664 66004
rect 327132 65952 327184 66004
rect 173860 65680 173912 65732
rect 178828 65680 178880 65732
rect 80204 65408 80256 65460
rect 87288 65408 87340 65460
rect 266596 65408 266648 65460
rect 274784 65408 274836 65460
rect 82780 65340 82832 65392
rect 87196 65340 87248 65392
rect 131356 65340 131408 65392
rect 136784 65340 136836 65392
rect 225932 65340 225984 65392
rect 233476 65340 233528 65392
rect 272668 65340 272720 65392
rect 274876 65340 274928 65392
rect 85080 65272 85132 65324
rect 87472 65272 87524 65324
rect 132184 65272 132236 65324
rect 135956 65272 136008 65324
rect 226208 65272 226260 65324
rect 233660 65272 233712 65324
rect 173492 64864 173544 64916
rect 175884 64864 175936 64916
rect 321612 64592 321664 64644
rect 327224 64592 327276 64644
rect 79468 64456 79520 64508
rect 82412 64456 82464 64508
rect 229428 64320 229480 64372
rect 233476 64320 233528 64372
rect 321612 64116 321664 64168
rect 328236 64116 328288 64168
rect 266596 64048 266648 64100
rect 273404 64048 273456 64100
rect 132368 63980 132420 64032
rect 136140 63980 136192 64032
rect 179104 63980 179156 64032
rect 182324 63980 182376 64032
rect 225748 63980 225800 64032
rect 234212 63980 234264 64032
rect 320508 63640 320560 63692
rect 326948 63640 327000 63692
rect 80204 62960 80256 63012
rect 82596 62960 82648 63012
rect 80204 62688 80256 62740
rect 85724 62688 85776 62740
rect 174044 62688 174096 62740
rect 178276 62688 178328 62740
rect 266596 62688 266648 62740
rect 272852 62688 272904 62740
rect 173492 62620 173544 62672
rect 175608 62620 175660 62672
rect 230440 62620 230492 62672
rect 233476 62620 233528 62672
rect 266688 62620 266740 62672
rect 274876 62620 274928 62672
rect 82412 62552 82464 62604
rect 87196 62552 87248 62604
rect 131724 62552 131776 62604
rect 139636 62552 139688 62604
rect 175884 62552 175936 62604
rect 181588 62552 181640 62604
rect 226300 62552 226352 62604
rect 234396 62552 234448 62604
rect 273404 62552 273456 62604
rect 274968 62552 275020 62604
rect 321060 62552 321112 62604
rect 327132 62552 327184 62604
rect 131356 62484 131408 62536
rect 139912 62484 139964 62536
rect 178828 62484 178880 62536
rect 182324 62484 182376 62536
rect 173124 61600 173176 61652
rect 175516 61600 175568 61652
rect 320692 61532 320744 61584
rect 327316 61532 327368 61584
rect 226300 61396 226352 61448
rect 229428 61396 229480 61448
rect 80204 61328 80256 61380
rect 81676 61328 81728 61380
rect 230532 61260 230584 61312
rect 233476 61260 233528 61312
rect 266596 61260 266648 61312
rect 272760 61260 272812 61312
rect 82596 61192 82648 61244
rect 87196 61192 87248 61244
rect 131356 61192 131408 61244
rect 139728 61192 139780 61244
rect 175608 61192 175660 61244
rect 181220 61192 181272 61244
rect 225748 61192 225800 61244
rect 230440 61192 230492 61244
rect 173124 60512 173176 60564
rect 175792 60512 175844 60564
rect 321060 60240 321112 60292
rect 328420 60240 328472 60292
rect 80204 60104 80256 60156
rect 81768 60104 81820 60156
rect 230624 59900 230676 59952
rect 233476 59900 233528 59952
rect 266596 59900 266648 59952
rect 272668 59900 272720 59952
rect 131356 59832 131408 59884
rect 139820 59832 139872 59884
rect 175516 59832 175568 59884
rect 181128 59832 181180 59884
rect 226300 59832 226352 59884
rect 233568 59832 233620 59884
rect 272760 59832 272812 59884
rect 275428 59832 275480 59884
rect 358412 59832 358464 59884
rect 358596 59832 358648 59884
rect 131448 59764 131500 59816
rect 139636 59764 139688 59816
rect 272852 59764 272904 59816
rect 275704 59764 275756 59816
rect 85724 59696 85776 59748
rect 87840 59696 87892 59748
rect 178276 59696 178328 59748
rect 181036 59696 181088 59748
rect 81676 59492 81728 59544
rect 87196 59492 87248 59544
rect 225748 59424 225800 59476
rect 230532 59424 230584 59476
rect 173032 58744 173084 58796
rect 175700 58744 175752 58796
rect 320508 58676 320560 58728
rect 327224 58676 327276 58728
rect 79652 58608 79704 58660
rect 82964 58608 83016 58660
rect 173584 58608 173636 58660
rect 175608 58608 175660 58660
rect 267884 58608 267936 58660
rect 272116 58608 272168 58660
rect 80204 58540 80256 58592
rect 82412 58540 82464 58592
rect 267332 58540 267384 58592
rect 272300 58540 272352 58592
rect 320416 58540 320468 58592
rect 328328 58540 328380 58592
rect 81768 58472 81820 58524
rect 87196 58472 87248 58524
rect 131356 58472 131408 58524
rect 139728 58472 139780 58524
rect 175792 58472 175844 58524
rect 181036 58472 181088 58524
rect 225564 58472 225616 58524
rect 230624 58472 230676 58524
rect 272668 58472 272720 58524
rect 275704 58472 275756 58524
rect 320416 57792 320468 57844
rect 328420 57792 328472 57844
rect 267700 57384 267752 57436
rect 272208 57384 272260 57436
rect 80204 57112 80256 57164
rect 81860 57112 81912 57164
rect 88300 57112 88352 57164
rect 173308 57112 173360 57164
rect 175516 57112 175568 57164
rect 317564 57155 317616 57164
rect 317564 57121 317573 57155
rect 317573 57121 317607 57155
rect 317607 57121 317616 57155
rect 317564 57112 317616 57121
rect 82964 57044 83016 57096
rect 87196 57044 87248 57096
rect 132184 57044 132236 57096
rect 140372 57044 140424 57096
rect 226300 57044 226352 57096
rect 233660 57044 233712 57096
rect 272300 57044 272352 57096
rect 275704 57044 275756 57096
rect 82412 56976 82464 57028
rect 87288 56976 87340 57028
rect 131356 56976 131408 57028
rect 140464 56976 140516 57028
rect 225656 56976 225708 57028
rect 233476 56976 233528 57028
rect 272116 56976 272168 57028
rect 275244 56976 275296 57028
rect 175608 56568 175660 56620
rect 181128 56568 181180 56620
rect 175700 56500 175752 56552
rect 181036 56500 181088 56552
rect 320416 56500 320468 56552
rect 327500 56500 327552 56552
rect 320508 56296 320560 56348
rect 328604 56296 328656 56348
rect 173492 56024 173544 56076
rect 175608 56024 175660 56076
rect 78916 55752 78968 55804
rect 82964 55752 83016 55804
rect 136508 55752 136560 55804
rect 140464 55752 140516 55804
rect 226484 55752 226536 55804
rect 233476 55752 233528 55804
rect 267332 55752 267384 55804
rect 272116 55752 272168 55804
rect 13136 55684 13188 55736
rect 16356 55684 16408 55736
rect 81860 55684 81912 55736
rect 87196 55684 87248 55736
rect 131356 55684 131408 55736
rect 140280 55684 140332 55736
rect 175516 55684 175568 55736
rect 181036 55684 181088 55736
rect 226392 55684 226444 55736
rect 233568 55684 233620 55736
rect 272208 55684 272260 55736
rect 275428 55684 275480 55736
rect 320416 55616 320468 55668
rect 328420 55616 328472 55668
rect 129424 55004 129476 55056
rect 140648 55004 140700 55056
rect 223448 55004 223500 55056
rect 233476 55004 233528 55056
rect 317564 55004 317616 55056
rect 328512 55004 328564 55056
rect 80204 54392 80256 54444
rect 82964 54256 83016 54308
rect 87196 54256 87248 54308
rect 134116 54392 134168 54444
rect 140372 54392 140424 54444
rect 173584 54392 173636 54444
rect 131356 54324 131408 54376
rect 136508 54324 136560 54376
rect 134116 54256 134168 54308
rect 233476 54392 233528 54444
rect 267884 54392 267936 54444
rect 272116 54324 272168 54376
rect 275704 54324 275756 54376
rect 328420 54392 328472 54444
rect 175608 54188 175660 54240
rect 181036 54188 181088 54240
rect 369176 54256 369228 54308
rect 369544 54256 369596 54308
rect 320416 54188 320468 54240
rect 327500 54188 327552 54240
rect 123536 54120 123588 54172
rect 217560 54120 217612 54172
rect 311584 54120 311636 54172
rect 80204 53644 80256 53696
rect 118660 53644 118712 53696
rect 140556 53644 140608 53696
rect 173584 53644 173636 53696
rect 212500 53644 212552 53696
rect 233476 53644 233528 53696
rect 267884 53644 267936 53696
rect 306616 53644 306668 53696
rect 328420 53644 328472 53696
rect 207900 53236 207952 53288
rect 80204 52964 80256 53016
rect 113968 52964 114020 53016
rect 140004 52964 140056 53016
rect 171836 52964 171888 53016
rect 267884 52964 267936 53016
rect 301648 52964 301700 53016
rect 233476 52896 233528 52948
rect 328512 52896 328564 52948
rect 91244 51536 91296 51588
rect 134760 51536 134812 51588
rect 187292 51536 187344 51588
rect 232096 51536 232148 51588
rect 279016 51536 279068 51588
rect 323820 51536 323872 51588
rect 88300 51468 88352 51520
rect 93636 51468 93688 51520
rect 184992 51468 185044 51520
rect 228692 51468 228744 51520
rect 312780 51468 312832 51520
rect 314252 51468 314304 51520
rect 314804 51468 314856 51520
rect 316644 51468 316696 51520
rect 220964 51400 221016 51452
rect 222620 51400 222672 51452
rect 125100 51264 125152 51316
rect 125928 51264 125980 51316
rect 111944 51128 111996 51180
rect 121236 51128 121288 51180
rect 205784 51128 205836 51180
rect 215536 51128 215588 51180
rect 299624 51128 299676 51180
rect 309560 51128 309612 51180
rect 106424 51060 106476 51112
rect 119120 51060 119172 51112
rect 200264 51060 200316 51112
rect 213236 51060 213288 51112
rect 294104 51060 294156 51112
rect 307260 51060 307312 51112
rect 102284 50992 102336 51044
rect 116544 50992 116596 51044
rect 196124 50992 196176 51044
rect 210844 50992 210896 51044
rect 289964 50992 290016 51044
rect 304868 50992 304920 51044
rect 114152 50924 114204 50976
rect 170456 50924 170508 50976
rect 189684 50924 189736 50976
rect 190604 50924 190656 50976
rect 208452 50924 208504 50976
rect 218940 50924 218992 50976
rect 220228 50924 220280 50976
rect 284444 50924 284496 50976
rect 302476 50924 302528 50976
rect 91244 50856 91296 50908
rect 112036 50856 112088 50908
rect 116084 50856 116136 50908
rect 123628 50856 123680 50908
rect 185084 50856 185136 50908
rect 206152 50856 206204 50908
rect 280304 50856 280356 50908
rect 300176 50856 300228 50908
rect 305144 50856 305196 50908
rect 311952 50856 312004 50908
rect 127124 50380 127176 50432
rect 128688 50380 128740 50432
rect 211304 50380 211356 50432
rect 217928 50380 217980 50432
rect 78916 50312 78968 50364
rect 108632 50312 108684 50364
rect 140648 50312 140700 50364
rect 173308 50312 173360 50364
rect 202564 50312 202616 50364
rect 233568 50312 233620 50364
rect 267516 50312 267568 50364
rect 296588 50312 296640 50364
rect 327684 50312 327736 50364
rect 80204 50244 80256 50296
rect 103572 50244 103624 50296
rect 140372 50244 140424 50296
rect 173584 50244 173636 50296
rect 197504 50244 197556 50296
rect 233476 50244 233528 50296
rect 266780 50244 266832 50296
rect 291528 50244 291580 50296
rect 328420 50244 328472 50296
rect 88392 49496 88444 49548
rect 102376 49496 102428 49548
rect 182140 49496 182192 49548
rect 194376 49496 194428 49548
rect 276164 49496 276216 49548
rect 288400 49496 288452 49548
rect 80204 48884 80256 48936
rect 98604 48884 98656 48936
rect 140556 48884 140608 48936
rect 172940 48884 172992 48936
rect 192536 48884 192588 48936
rect 233476 48884 233528 48936
rect 267884 48884 267936 48936
rect 286560 48884 286612 48936
rect 328420 48884 328472 48936
rect 96764 48519 96816 48528
rect 96764 48485 96773 48519
rect 96773 48485 96807 48519
rect 96807 48485 96816 48519
rect 96764 48476 96816 48485
rect 181864 48136 181916 48188
rect 182232 48136 182284 48188
rect 196676 48136 196728 48188
rect 232096 48136 232148 48188
rect 238628 48136 238680 48188
rect 241112 48136 241164 48188
rect 276072 48136 276124 48188
rect 293092 48136 293144 48188
rect 80204 47660 80256 47712
rect 140004 47660 140056 47712
rect 93728 47524 93780 47576
rect 142856 47524 142908 47576
rect 159508 47524 159560 47576
rect 100260 47456 100312 47508
rect 100444 47456 100496 47508
rect 156840 47456 156892 47508
rect 167696 47456 167748 47508
rect 173308 47456 173360 47508
rect 187568 47456 187620 47508
rect 233476 47456 233528 47508
rect 267884 47456 267936 47508
rect 281592 47456 281644 47508
rect 327868 47456 327920 47508
rect 60700 47388 60752 47440
rect 74224 47388 74276 47440
rect 295484 47388 295536 47440
rect 353628 47388 353680 47440
rect 419776 47388 419828 47440
rect 286008 47320 286060 47372
rect 338356 47320 338408 47372
rect 74684 46776 74736 46828
rect 88116 46776 88168 46828
rect 88024 46708 88076 46760
rect 100260 46708 100312 46760
rect 275980 46708 276032 46760
rect 295484 46708 295536 46760
rect 338356 46640 338408 46692
rect 339644 46640 339696 46692
rect 73120 46164 73172 46216
rect 88208 46164 88260 46216
rect 106608 46164 106660 46216
rect 74224 46096 74276 46148
rect 88024 46096 88076 46148
rect 88116 46096 88168 46148
rect 109460 46096 109512 46148
rect 317472 46139 317524 46148
rect 317472 46105 317481 46139
rect 317481 46105 317515 46139
rect 317515 46105 317524 46139
rect 317472 46096 317524 46105
rect 167236 46028 167288 46080
rect 169720 46028 169772 46080
rect 298244 46071 298296 46080
rect 298244 46037 298253 46071
rect 298253 46037 298287 46071
rect 298287 46037 298296 46071
rect 298244 46028 298296 46037
rect 350132 46028 350184 46080
rect 361080 46028 361132 46080
rect 53708 45960 53760 46012
rect 95476 45960 95528 46012
rect 144696 45960 144748 46012
rect 369728 45960 369780 46012
rect 57204 45892 57256 45944
rect 98052 45892 98104 45944
rect 153436 45892 153488 45944
rect 238628 45892 238680 45944
rect 322532 45892 322584 45944
rect 332652 45892 332704 45944
rect 369820 45892 369872 45944
rect 95476 45824 95528 45876
rect 95752 45824 95804 45876
rect 150584 45824 150636 45876
rect 170180 45824 170232 45876
rect 250956 45824 251008 45876
rect 275520 45824 275572 45876
rect 276164 45824 276216 45876
rect 357124 45824 357176 45876
rect 253992 45756 254044 45808
rect 262548 45756 262600 45808
rect 263100 45756 263152 45808
rect 284352 45756 284404 45808
rect 336148 45756 336200 45808
rect 347924 45756 347976 45808
rect 359700 45756 359752 45808
rect 50212 45688 50264 45740
rect 369176 45688 369228 45740
rect 169536 45348 169588 45400
rect 181956 45348 182008 45400
rect 182048 45348 182100 45400
rect 201460 45348 201512 45400
rect 276072 45348 276124 45400
rect 290700 45348 290752 45400
rect 324556 45348 324608 45400
rect 346636 45348 346688 45400
rect 347924 45348 347976 45400
rect 357124 45348 357176 45400
rect 376996 45348 377048 45400
rect 422536 45348 422588 45400
rect 262824 45280 262876 45332
rect 275888 45280 275940 45332
rect 317472 44804 317524 44856
rect 169720 44736 169772 44788
rect 182048 44736 182100 44788
rect 263100 44736 263152 44788
rect 276072 44736 276124 44788
rect 12860 42560 12912 42612
rect 16264 42560 16316 42612
rect 358412 40631 358464 40640
rect 358412 40597 358421 40631
rect 358421 40597 358455 40631
rect 358455 40597 358464 40631
rect 358412 40588 358464 40597
rect 317104 37843 317156 37852
rect 317104 37809 317113 37843
rect 317113 37809 317147 37843
rect 317147 37809 317156 37843
rect 317104 37800 317156 37809
rect 358412 37843 358464 37852
rect 358412 37809 358421 37843
rect 358421 37809 358455 37843
rect 358455 37809 358464 37843
rect 358412 37800 358464 37809
rect 101364 37732 101416 37784
rect 102284 37732 102336 37784
rect 210016 37732 210068 37784
rect 211304 37732 211356 37784
rect 215076 37732 215128 37784
rect 218940 37732 218992 37784
rect 220044 37732 220096 37784
rect 220964 37732 221016 37784
rect 289044 37732 289096 37784
rect 289964 37732 290016 37784
rect 304040 37732 304092 37784
rect 305144 37732 305196 37784
rect 96396 37460 96448 37512
rect 96764 37460 96816 37512
rect 195020 37392 195072 37444
rect 196124 37392 196176 37444
rect 279108 37324 279160 37376
rect 280304 37324 280356 37376
rect 121420 37120 121472 37172
rect 125100 37120 125152 37172
rect 314068 37120 314120 37172
rect 314804 37120 314856 37172
rect 309100 36712 309152 36764
rect 312780 36712 312832 36764
rect 111392 36644 111444 36696
rect 111944 36644 111996 36696
rect 126388 36576 126440 36628
rect 127124 36576 127176 36628
rect 276164 33040 276216 33092
rect 369636 33040 369688 33092
rect 182324 32972 182376 33024
rect 369452 32972 369504 33024
rect 88484 32904 88536 32956
rect 369176 32904 369228 32956
rect 12676 29436 12728 29488
rect 16172 29436 16224 29488
rect 358228 28119 358280 28128
rect 358228 28085 358237 28119
rect 358237 28085 358271 28119
rect 358271 28085 358280 28119
rect 358228 28076 358280 28085
rect 427504 28076 427556 28128
rect 429804 28076 429856 28128
rect 358320 18488 358372 18540
rect 185176 17060 185228 17112
rect 186372 17060 186424 17112
rect 191340 17060 191392 17112
rect 192076 17060 192128 17112
rect 196124 17060 196176 17112
rect 196308 17060 196360 17112
rect 92624 16788 92676 16840
rect 105136 16788 105188 16840
rect 80756 16720 80808 16772
rect 102376 16720 102428 16772
rect 285364 16720 285416 16772
rect 299716 16720 299768 16772
rect 67876 16652 67928 16704
rect 107068 16652 107120 16704
rect 170916 16652 170968 16704
rect 201368 16652 201420 16704
rect 273956 16652 274008 16704
rect 295392 16652 295444 16704
rect 54996 16584 55048 16636
rect 112036 16584 112088 16636
rect 158036 16584 158088 16636
rect 206336 16584 206388 16636
rect 261076 16584 261128 16636
rect 300360 16584 300412 16636
rect 29236 16516 29288 16568
rect 122064 16516 122116 16568
rect 145156 16516 145208 16568
rect 211304 16516 211356 16568
rect 248196 16516 248248 16568
rect 305328 16516 305380 16568
rect 42116 16448 42168 16500
rect 117004 16448 117056 16500
rect 119396 16448 119448 16500
rect 221332 16448 221384 16500
rect 235316 16448 235368 16500
rect 310388 16448 310440 16500
rect 16356 16380 16408 16432
rect 127216 16380 127268 16432
rect 132276 16380 132328 16432
rect 216364 16380 216416 16432
rect 222436 16380 222488 16432
rect 315356 16380 315408 16432
rect 13044 15564 13096 15616
rect 16080 15564 16132 15616
rect 427320 15428 427372 15480
rect 429436 15428 429488 15480
rect 351236 12912 351288 12964
rect 358320 12912 358372 12964
rect 286836 12436 286888 12488
rect 290056 12436 290108 12488
rect 280396 12368 280448 12420
rect 312596 12368 312648 12420
rect 105136 12300 105188 12352
rect 106516 12300 106568 12352
rect 183796 12300 183848 12352
rect 196124 12300 196176 12352
rect 265860 12300 265912 12352
rect 402756 12300 402808 12352
rect 93636 12232 93688 12284
rect 96856 12232 96908 12284
rect 185176 12232 185228 12284
rect 209556 12232 209608 12284
rect 228600 12232 228652 12284
rect 415636 12232 415688 12284
rect 192076 12096 192128 12148
rect 196676 12096 196728 12148
rect 385184 12096 385236 12148
rect 389876 12096 389928 12148
rect 324556 9376 324608 9428
rect 325476 9376 325528 9428
rect 428056 9376 428108 9428
rect 428516 9376 428568 9428
<< metal2 >>
rect 18746 396344 18802 396824
rect 36410 396344 36466 396824
rect 54166 396344 54222 396824
rect 71830 396344 71886 396824
rect 89586 396344 89642 396824
rect 107250 396344 107306 396824
rect 125006 396344 125062 396824
rect 142670 396344 142726 396824
rect 160426 396344 160482 396824
rect 178090 396344 178146 396824
rect 195846 396344 195902 396824
rect 213510 396344 213566 396824
rect 231266 396344 231322 396824
rect 248930 396344 248986 396824
rect 266686 396344 266742 396824
rect 284350 396344 284406 396824
rect 302106 396344 302162 396824
rect 319770 396344 319826 396824
rect 337526 396344 337582 396824
rect 355190 396344 355246 396824
rect 372946 396344 373002 396824
rect 390610 396344 390666 396824
rect 408366 396344 408422 396824
rect 426030 396344 426086 396824
rect 18760 392818 18788 396344
rect 36424 396234 36452 396344
rect 54180 396234 54208 396344
rect 36148 396206 36452 396234
rect 54088 396206 54208 396234
rect 18196 392812 18248 392818
rect 18196 392754 18248 392760
rect 18748 392812 18800 392818
rect 18748 392754 18800 392760
rect 13318 390128 13374 390137
rect 13318 390063 13374 390072
rect 12676 283400 12728 283406
rect 12676 283342 12728 283348
rect 12688 283105 12716 283342
rect 12674 283096 12730 283105
rect 12674 283031 12730 283040
rect 12860 270072 12912 270078
rect 12860 270014 12912 270020
rect 12872 269777 12900 270014
rect 12858 269768 12914 269777
rect 12858 269703 12914 269712
rect 13332 269602 13360 390063
rect 18208 389010 18236 392754
rect 36148 389146 36176 396206
rect 54088 389282 54116 396206
rect 71844 393702 71872 396344
rect 89600 393838 89628 396344
rect 107264 393838 107292 396344
rect 125020 393838 125048 396344
rect 88576 393832 88628 393838
rect 88576 393774 88628 393780
rect 89588 393832 89640 393838
rect 89588 393774 89640 393780
rect 106516 393832 106568 393838
rect 106516 393774 106568 393780
rect 107252 393832 107304 393838
rect 107252 393774 107304 393780
rect 124456 393832 124508 393838
rect 124456 393774 124508 393780
rect 125008 393832 125060 393838
rect 125008 393774 125060 393780
rect 70636 393696 70688 393702
rect 70636 393638 70688 393644
rect 71832 393696 71884 393702
rect 71832 393638 71884 393644
rect 70648 389350 70676 393638
rect 70636 389344 70688 389350
rect 70636 389286 70688 389292
rect 54076 389276 54128 389282
rect 54076 389218 54128 389224
rect 36136 389140 36188 389146
rect 36136 389082 36188 389088
rect 88588 389078 88616 393774
rect 106332 393220 106384 393226
rect 106332 393162 106384 393168
rect 91336 393152 91388 393158
rect 91336 393094 91388 393100
rect 88576 389072 88628 389078
rect 88576 389014 88628 389020
rect 18196 389004 18248 389010
rect 18196 388946 18248 388952
rect 13412 388528 13464 388534
rect 13412 388470 13464 388476
rect 13424 350017 13452 388470
rect 13504 388460 13556 388466
rect 13504 388402 13556 388408
rect 13516 363345 13544 388402
rect 13596 388392 13648 388398
rect 13596 388334 13648 388340
rect 13608 376809 13636 388334
rect 91348 386700 91376 393094
rect 96304 388596 96356 388602
rect 96304 388538 96356 388544
rect 96316 386700 96344 388538
rect 101272 388528 101324 388534
rect 101272 388470 101324 388476
rect 101284 386700 101312 388470
rect 106344 386700 106372 393162
rect 106528 389214 106556 393774
rect 111300 389344 111352 389350
rect 111300 389286 111352 389292
rect 106516 389208 106568 389214
rect 106516 389150 106568 389156
rect 111312 386700 111340 389286
rect 124468 389282 124496 393774
rect 142684 389282 142712 396344
rect 116268 389276 116320 389282
rect 116268 389218 116320 389224
rect 124456 389276 124508 389282
rect 124456 389218 124508 389224
rect 142672 389276 142724 389282
rect 142672 389218 142724 389224
rect 116280 386700 116308 389218
rect 121328 389140 121380 389146
rect 121328 389082 121380 389088
rect 121340 386700 121368 389082
rect 160440 389010 160468 396344
rect 178104 389146 178132 396344
rect 195860 389282 195888 396344
rect 213524 393838 213552 396344
rect 231280 396234 231308 396344
rect 231004 396206 231308 396234
rect 248944 396234 248972 396344
rect 266700 396234 266728 396344
rect 248944 396206 249064 396234
rect 212776 393832 212828 393838
rect 212776 393774 212828 393780
rect 213512 393832 213564 393838
rect 213512 393774 213564 393780
rect 194836 389276 194888 389282
rect 194836 389218 194888 389224
rect 195848 389276 195900 389282
rect 195848 389218 195900 389224
rect 178092 389140 178144 389146
rect 178092 389082 178144 389088
rect 126296 389004 126348 389010
rect 126296 388946 126348 388952
rect 160428 389004 160480 389010
rect 160428 388946 160480 388952
rect 126308 386700 126336 388946
rect 127860 388596 127912 388602
rect 127860 388538 127912 388544
rect 185360 388596 185412 388602
rect 185360 388538 185412 388544
rect 13594 376800 13650 376809
rect 13594 376735 13650 376744
rect 89864 367720 89916 367726
rect 89864 367662 89916 367668
rect 13502 363336 13558 363345
rect 13502 363271 13558 363280
rect 67692 359900 67744 359906
rect 67692 359842 67744 359848
rect 75972 359900 76024 359906
rect 75972 359842 76024 359848
rect 53708 359832 53760 359838
rect 53708 359774 53760 359780
rect 50212 359764 50264 359770
rect 50212 359706 50264 359712
rect 50224 357732 50252 359706
rect 53720 357732 53748 359774
rect 64196 359696 64248 359702
rect 64196 359638 64248 359644
rect 60700 359628 60752 359634
rect 60700 359570 60752 359576
rect 57204 359560 57256 359566
rect 57204 359502 57256 359508
rect 57216 357732 57244 359502
rect 60712 357732 60740 359570
rect 64208 357732 64236 359638
rect 67704 357732 67732 359842
rect 75696 359696 75748 359702
rect 75696 359638 75748 359644
rect 71188 359424 71240 359430
rect 71188 359366 71240 359372
rect 71200 357732 71228 359366
rect 75708 357594 75736 359638
rect 75788 359628 75840 359634
rect 75788 359570 75840 359576
rect 75696 357588 75748 357594
rect 75696 357530 75748 357536
rect 75800 357526 75828 359570
rect 75880 359424 75932 359430
rect 75880 359366 75932 359372
rect 75788 357520 75840 357526
rect 74710 357458 74816 357474
rect 75788 357462 75840 357468
rect 74710 357452 74828 357458
rect 74710 357446 74776 357452
rect 74776 357394 74828 357400
rect 13410 350008 13466 350017
rect 13410 349943 13466 349952
rect 13410 336680 13466 336689
rect 13410 336615 13466 336624
rect 13320 269596 13372 269602
rect 13320 269538 13372 269544
rect 13424 262598 13452 336615
rect 75892 334746 75920 359366
rect 75984 334814 76012 359842
rect 76984 359832 77036 359838
rect 76984 359774 77036 359780
rect 76800 359764 76852 359770
rect 76800 359706 76852 359712
rect 76064 359560 76116 359566
rect 76064 359502 76116 359508
rect 76076 354058 76104 359502
rect 76432 357588 76484 357594
rect 76432 357530 76484 357536
rect 76156 357520 76208 357526
rect 76156 357462 76208 357468
rect 76064 354052 76116 354058
rect 76064 353994 76116 354000
rect 76062 353952 76118 353961
rect 76062 353887 76118 353896
rect 76076 344130 76104 353887
rect 76168 344130 76196 357462
rect 76444 353961 76472 357530
rect 76430 353952 76486 353961
rect 76248 353916 76300 353922
rect 76430 353887 76486 353896
rect 76248 353858 76300 353864
rect 76064 344124 76116 344130
rect 76064 344066 76116 344072
rect 76156 344124 76208 344130
rect 76156 344066 76208 344072
rect 76260 343874 76288 353858
rect 76076 343846 76288 343874
rect 75972 334808 76024 334814
rect 75972 334750 76024 334756
rect 76076 334746 76104 343846
rect 76156 343784 76208 343790
rect 76156 343726 76208 343732
rect 75880 334740 75932 334746
rect 75880 334682 75932 334688
rect 76064 334740 76116 334746
rect 76064 334682 76116 334688
rect 76168 334626 76196 343726
rect 75892 334598 76196 334626
rect 75892 334406 75920 334598
rect 75972 334536 76024 334542
rect 75972 334478 76024 334484
rect 76064 334536 76116 334542
rect 76064 334478 76116 334484
rect 75880 334400 75932 334406
rect 75880 334342 75932 334348
rect 75512 330184 75564 330190
rect 75512 330126 75564 330132
rect 75420 330116 75472 330122
rect 75420 330058 75472 330064
rect 48568 329838 48950 329866
rect 13962 323216 14018 323225
rect 13962 323151 14018 323160
rect 13976 322166 14004 323151
rect 13964 322160 14016 322166
rect 13964 322102 14016 322108
rect 16356 322160 16408 322166
rect 16356 322102 16408 322108
rect 16078 313832 16134 313841
rect 16078 313767 16134 313776
rect 13962 309888 14018 309897
rect 13962 309823 14018 309832
rect 13976 309722 14004 309823
rect 13964 309716 14016 309722
rect 13964 309658 14016 309664
rect 13686 296424 13742 296433
rect 13686 296359 13742 296368
rect 13700 296190 13728 296359
rect 13688 296184 13740 296190
rect 13688 296126 13740 296132
rect 14700 293192 14752 293198
rect 14700 293134 14752 293140
rect 14712 283406 14740 293134
rect 14700 283400 14752 283406
rect 14700 283342 14752 283348
rect 13412 262592 13464 262598
rect 13412 262534 13464 262540
rect 12860 256608 12912 256614
rect 12860 256550 12912 256556
rect 12872 256313 12900 256550
rect 12858 256304 12914 256313
rect 12858 256239 12914 256248
rect 13136 243416 13188 243422
rect 13136 243358 13188 243364
rect 13148 242985 13176 243358
rect 13134 242976 13190 242985
rect 13134 242911 13190 242920
rect 13042 229648 13098 229657
rect 16092 229618 16120 313767
rect 16170 308392 16226 308401
rect 16170 308327 16226 308336
rect 16184 243422 16212 308327
rect 16262 304176 16318 304185
rect 16262 304111 16318 304120
rect 16276 256614 16304 304111
rect 16368 280686 16396 322102
rect 38804 315904 38856 315910
rect 38804 315846 38856 315852
rect 38816 315609 38844 315846
rect 38802 315600 38858 315609
rect 38802 315535 38858 315544
rect 38436 313796 38488 313802
rect 38436 313738 38488 313744
rect 38448 313161 38476 313738
rect 38434 313152 38490 313161
rect 38434 313087 38490 313096
rect 38802 310432 38858 310441
rect 38802 310367 38858 310376
rect 38816 310334 38844 310367
rect 38804 310328 38856 310334
rect 38804 310270 38856 310276
rect 16540 309716 16592 309722
rect 16540 309658 16592 309664
rect 16446 298736 16502 298745
rect 16446 298671 16502 298680
rect 16356 280680 16408 280686
rect 16356 280622 16408 280628
rect 16460 270078 16488 298671
rect 16552 283513 16580 309658
rect 38804 308288 38856 308294
rect 38804 308230 38856 308236
rect 38816 308129 38844 308230
rect 38802 308120 38858 308129
rect 38802 308055 38858 308064
rect 38804 306248 38856 306254
rect 38804 306190 38856 306196
rect 38816 305681 38844 306190
rect 38802 305672 38858 305681
rect 38802 305607 38858 305616
rect 38620 304140 38672 304146
rect 38620 304082 38672 304088
rect 38632 303097 38660 304082
rect 38618 303088 38674 303097
rect 38618 303023 38674 303032
rect 38804 300672 38856 300678
rect 38802 300640 38804 300649
rect 38856 300640 38858 300649
rect 38802 300575 38858 300584
rect 38252 298632 38304 298638
rect 38252 298574 38304 298580
rect 38264 298201 38292 298574
rect 38250 298192 38306 298201
rect 38250 298127 38306 298136
rect 16724 296184 16776 296190
rect 16724 296126 16776 296132
rect 16736 289089 16764 296126
rect 38802 295472 38858 295481
rect 38802 295407 38858 295416
rect 38816 295170 38844 295407
rect 38804 295164 38856 295170
rect 38804 295106 38856 295112
rect 17458 293840 17514 293849
rect 17458 293775 17514 293784
rect 38436 293804 38488 293810
rect 17472 293198 17500 293775
rect 38436 293746 38488 293752
rect 17460 293192 17512 293198
rect 38448 293169 38476 293746
rect 17460 293134 17512 293140
rect 38434 293160 38490 293169
rect 38434 293095 38490 293104
rect 38620 291696 38672 291702
rect 38620 291638 38672 291644
rect 38632 290585 38660 291638
rect 38618 290576 38674 290585
rect 38618 290511 38674 290520
rect 16722 289080 16778 289089
rect 16722 289015 16778 289024
rect 38804 288976 38856 288982
rect 38804 288918 38856 288924
rect 38816 288137 38844 288918
rect 38802 288128 38858 288137
rect 38802 288063 38858 288072
rect 38802 285544 38858 285553
rect 38802 285479 38804 285488
rect 38856 285479 38858 285488
rect 38804 285450 38856 285456
rect 16538 283504 16594 283513
rect 16538 283439 16594 283448
rect 38068 283468 38120 283474
rect 38068 283410 38120 283416
rect 38080 283105 38108 283410
rect 38066 283096 38122 283105
rect 38066 283031 38122 283040
rect 16724 280680 16776 280686
rect 16724 280622 16776 280628
rect 16736 279433 16764 280622
rect 38066 280376 38122 280385
rect 38066 280311 38122 280320
rect 38080 280006 38108 280311
rect 48568 280006 48596 329838
rect 49948 285514 49976 329852
rect 50040 329838 50974 329866
rect 51328 329838 51986 329866
rect 50040 291702 50068 329838
rect 51222 313832 51278 313841
rect 51222 313767 51224 313776
rect 51276 313767 51278 313776
rect 51224 313738 51276 313744
rect 51222 308664 51278 308673
rect 51222 308599 51278 308608
rect 51236 308294 51264 308599
rect 51224 308288 51276 308294
rect 51224 308230 51276 308236
rect 50304 300672 50356 300678
rect 50302 300640 50304 300649
rect 50356 300640 50358 300649
rect 50302 300575 50358 300584
rect 51328 295170 51356 329838
rect 53076 327441 53104 329852
rect 54088 327441 54116 329852
rect 54824 329838 55114 329866
rect 53062 327432 53118 327441
rect 53062 327367 53118 327376
rect 54074 327432 54130 327441
rect 54074 327367 54130 327376
rect 54824 324886 54852 329838
rect 56112 327441 56140 329852
rect 56848 329838 57230 329866
rect 56098 327432 56154 327441
rect 56098 327367 56154 327376
rect 54076 324880 54128 324886
rect 54076 324822 54128 324828
rect 54812 324880 54864 324886
rect 54812 324822 54864 324828
rect 54088 317921 54116 324822
rect 56100 320324 56152 320330
rect 56100 320266 56152 320272
rect 55272 320188 55324 320194
rect 55272 320130 55324 320136
rect 54074 317912 54130 317921
rect 54074 317847 54130 317856
rect 55284 316796 55312 320130
rect 56112 316796 56140 320266
rect 56848 319718 56876 329838
rect 58228 320534 58256 329852
rect 59240 327402 59268 329852
rect 59608 329838 60266 329866
rect 60988 329838 61370 329866
rect 62382 329838 62488 329866
rect 58308 327396 58360 327402
rect 58308 327338 58360 327344
rect 59228 327396 59280 327402
rect 59228 327338 59280 327344
rect 58216 320528 58268 320534
rect 58216 320470 58268 320476
rect 57940 320460 57992 320466
rect 57940 320402 57992 320408
rect 56836 319712 56888 319718
rect 56836 319654 56888 319660
rect 57020 319644 57072 319650
rect 57020 319586 57072 319592
rect 57032 316796 57060 319586
rect 57952 316796 57980 320402
rect 58320 319582 58348 327338
rect 59608 320126 59636 329838
rect 59688 320392 59740 320398
rect 59688 320334 59740 320340
rect 59596 320120 59648 320126
rect 59596 320062 59648 320068
rect 58768 319984 58820 319990
rect 58768 319926 58820 319932
rect 58308 319576 58360 319582
rect 58308 319518 58360 319524
rect 58780 316796 58808 319926
rect 59700 316796 59728 320334
rect 60608 320256 60660 320262
rect 60608 320198 60660 320204
rect 60620 316796 60648 320198
rect 60988 319854 61016 329838
rect 62356 327396 62408 327402
rect 62356 327338 62408 327344
rect 62368 320516 62396 327338
rect 62460 320670 62488 329838
rect 63380 327402 63408 329852
rect 63748 329838 64406 329866
rect 65312 329838 65510 329866
rect 63368 327396 63420 327402
rect 63368 327338 63420 327344
rect 62448 320664 62500 320670
rect 62448 320606 62500 320612
rect 63748 320602 63776 329838
rect 65208 327396 65260 327402
rect 65208 327338 65260 327344
rect 65116 326648 65168 326654
rect 65116 326590 65168 326596
rect 63736 320596 63788 320602
rect 63736 320538 63788 320544
rect 65128 320534 65156 326590
rect 64104 320528 64156 320534
rect 62368 320488 62488 320516
rect 62356 320188 62408 320194
rect 62356 320130 62408 320136
rect 61436 320052 61488 320058
rect 61436 319994 61488 320000
rect 60976 319848 61028 319854
rect 60976 319790 61028 319796
rect 61448 316796 61476 319994
rect 62368 316796 62396 320130
rect 62460 319786 62488 320488
rect 64104 320470 64156 320476
rect 65116 320528 65168 320534
rect 65116 320470 65168 320476
rect 62448 319780 62500 319786
rect 62448 319722 62500 319728
rect 63276 319712 63328 319718
rect 63276 319654 63328 319660
rect 63288 316796 63316 319654
rect 64116 316796 64144 320470
rect 65220 320466 65248 327338
rect 65208 320460 65260 320466
rect 65208 320402 65260 320408
rect 65024 319576 65076 319582
rect 65024 319518 65076 319524
rect 65036 316796 65064 319518
rect 65312 319446 65340 329838
rect 65944 320120 65996 320126
rect 65944 320062 65996 320068
rect 65300 319440 65352 319446
rect 65300 319382 65352 319388
rect 65956 316796 65984 320062
rect 66508 319922 66536 329852
rect 66600 329838 67534 329866
rect 66600 320330 66628 329838
rect 68532 327402 68560 329852
rect 68520 327396 68572 327402
rect 68520 327338 68572 327344
rect 69636 326654 69664 329852
rect 70662 329838 70768 329866
rect 69624 326648 69676 326654
rect 69624 326590 69676 326596
rect 70636 325288 70688 325294
rect 70636 325230 70688 325236
rect 67692 320664 67744 320670
rect 67692 320606 67744 320612
rect 66588 320324 66640 320330
rect 66588 320266 66640 320272
rect 66496 319916 66548 319922
rect 66496 319858 66548 319864
rect 66772 319848 66824 319854
rect 66772 319790 66824 319796
rect 66784 316796 66812 319790
rect 67704 316796 67732 320606
rect 69440 320596 69492 320602
rect 69440 320538 69492 320544
rect 68612 319780 68664 319786
rect 68612 319722 68664 319728
rect 68624 316796 68652 319722
rect 69452 316796 69480 320538
rect 70648 320398 70676 325230
rect 70636 320392 70688 320398
rect 70636 320334 70688 320340
rect 70740 319990 70768 329838
rect 71384 329838 71674 329866
rect 72028 329838 72686 329866
rect 73408 329838 73790 329866
rect 71384 325294 71412 329838
rect 72028 326330 72056 329838
rect 71936 326302 72056 326330
rect 71372 325288 71424 325294
rect 71372 325230 71424 325236
rect 71936 320262 71964 326302
rect 71924 320256 71976 320262
rect 71924 320198 71976 320204
rect 73408 320058 73436 329838
rect 74040 326376 74092 326382
rect 74040 326318 74092 326324
rect 73396 320052 73448 320058
rect 73396 319994 73448 320000
rect 70728 319984 70780 319990
rect 70728 319926 70780 319932
rect 70360 319440 70412 319446
rect 70360 319382 70412 319388
rect 70372 316796 70400 319382
rect 52696 315904 52748 315910
rect 52694 315872 52696 315881
rect 52748 315872 52750 315881
rect 52694 315807 52750 315816
rect 54074 310432 54130 310441
rect 54074 310367 54130 310376
rect 54088 310334 54116 310367
rect 54076 310328 54128 310334
rect 54076 310270 54128 310276
rect 73394 307168 73450 307177
rect 73394 307103 73450 307112
rect 54444 306248 54496 306254
rect 54442 306216 54444 306225
rect 54496 306216 54498 306225
rect 54442 306151 54498 306160
rect 73408 305681 73436 307103
rect 73394 305672 73450 305681
rect 73394 305607 73450 305616
rect 51406 304176 51462 304185
rect 51406 304111 51408 304120
rect 51460 304111 51462 304120
rect 51408 304082 51460 304088
rect 51406 298872 51462 298881
rect 51406 298807 51462 298816
rect 51420 298638 51448 298807
rect 51408 298632 51460 298638
rect 51408 298574 51460 298580
rect 51316 295164 51368 295170
rect 51316 295106 51368 295112
rect 51328 293962 51356 295106
rect 51236 293934 51356 293962
rect 51236 293690 51264 293934
rect 51314 293840 51370 293849
rect 51314 293775 51316 293784
rect 51368 293775 51370 293784
rect 51316 293746 51368 293752
rect 51236 293662 51356 293690
rect 50028 291696 50080 291702
rect 50028 291638 50080 291644
rect 50040 291294 50068 291638
rect 50028 291288 50080 291294
rect 50028 291230 50080 291236
rect 51328 289202 51356 293662
rect 51684 291288 51736 291294
rect 51684 291230 51736 291236
rect 51236 289174 51356 289202
rect 51236 288794 51264 289174
rect 51314 289080 51370 289089
rect 51314 289015 51370 289024
rect 51328 288982 51356 289015
rect 51316 288976 51368 288982
rect 51316 288918 51368 288924
rect 51236 288766 51356 288794
rect 51696 288778 51724 291230
rect 74052 290177 74080 326318
rect 74788 320194 74816 329852
rect 74776 320188 74828 320194
rect 74776 320130 74828 320136
rect 74222 314512 74278 314521
rect 74222 314447 74278 314456
rect 74130 311112 74186 311121
rect 74130 311047 74186 311056
rect 74038 290168 74094 290177
rect 74038 290103 74094 290112
rect 49936 285508 49988 285514
rect 49936 285450 49988 285456
rect 38068 280000 38120 280006
rect 38068 279942 38120 279948
rect 48556 280000 48608 280006
rect 48556 279942 48608 279948
rect 16722 279424 16778 279433
rect 16722 279359 16778 279368
rect 38620 279320 38672 279326
rect 38620 279262 38672 279268
rect 38632 278209 38660 279262
rect 38618 278200 38674 278209
rect 38618 278135 38674 278144
rect 21244 273818 21272 276948
rect 23912 274498 23940 276948
rect 26580 274566 26608 276948
rect 29248 274634 29276 276948
rect 31916 274702 31944 276948
rect 34584 274770 34612 276948
rect 34572 274764 34624 274770
rect 34572 274706 34624 274712
rect 46992 274764 47044 274770
rect 46992 274706 47044 274712
rect 31904 274696 31956 274702
rect 31904 274638 31956 274644
rect 46624 274696 46676 274702
rect 46624 274638 46676 274644
rect 29236 274628 29288 274634
rect 29236 274570 29288 274576
rect 46532 274628 46584 274634
rect 46532 274570 46584 274576
rect 26568 274560 26620 274566
rect 26568 274502 26620 274508
rect 23900 274492 23952 274498
rect 23900 274434 23952 274440
rect 46440 274492 46492 274498
rect 46440 274434 46492 274440
rect 21232 273812 21284 273818
rect 21232 273754 21284 273760
rect 22244 273812 22296 273818
rect 22244 273754 22296 273760
rect 16448 270072 16500 270078
rect 16448 270014 16500 270020
rect 16264 256608 16316 256614
rect 16264 256550 16316 256556
rect 16172 243416 16224 243422
rect 16172 243358 16224 243364
rect 22256 229618 22284 273754
rect 46452 249785 46480 274434
rect 46544 256041 46572 274570
rect 46636 259169 46664 274638
rect 47004 262734 47032 274706
rect 47084 274560 47136 274566
rect 47084 274502 47136 274508
rect 47096 271681 47124 274502
rect 47082 271672 47138 271681
rect 47082 271607 47138 271616
rect 46992 262728 47044 262734
rect 46992 262670 47044 262676
rect 46622 259160 46678 259169
rect 46622 259095 46678 259104
rect 46530 256032 46586 256041
rect 46530 255967 46586 255976
rect 47096 252913 47124 271607
rect 48568 263906 48596 279942
rect 48568 263878 49148 263906
rect 49120 263770 49148 263878
rect 49948 263770 49976 285450
rect 51328 265114 51356 288766
rect 51408 288772 51460 288778
rect 51408 288714 51460 288720
rect 51684 288772 51736 288778
rect 51684 288714 51736 288720
rect 51316 265108 51368 265114
rect 51316 265050 51368 265056
rect 49120 263742 49410 263770
rect 49948 263742 50422 263770
rect 51420 263756 51448 288714
rect 51498 283776 51554 283785
rect 51498 283711 51554 283720
rect 51512 283542 51540 283711
rect 51500 283536 51552 283542
rect 51500 283478 51552 283484
rect 74144 280686 74172 311047
rect 74236 297210 74264 314447
rect 75432 299969 75460 330058
rect 75524 304049 75552 330126
rect 75800 326314 75828 329852
rect 75788 326308 75840 326314
rect 75788 326250 75840 326256
rect 75510 304040 75566 304049
rect 75510 303975 75566 303984
rect 75418 299960 75474 299969
rect 75418 299895 75474 299904
rect 74224 297204 74276 297210
rect 74224 297146 74276 297152
rect 74222 296968 74278 296977
rect 74222 296903 74278 296912
rect 74132 280680 74184 280686
rect 74132 280622 74184 280628
rect 51498 279424 51554 279433
rect 51498 279359 51554 279368
rect 51512 279326 51540 279359
rect 51500 279320 51552 279326
rect 51500 279262 51552 279268
rect 74038 278200 74094 278209
rect 74038 278135 74094 278144
rect 67152 277070 67718 277098
rect 69636 277070 70386 277098
rect 55298 276934 55404 276962
rect 56126 276934 56784 276962
rect 55376 266270 55404 276934
rect 55546 266640 55602 266649
rect 55546 266575 55602 266584
rect 55364 266264 55416 266270
rect 55364 266206 55416 266212
rect 53522 265552 53578 265561
rect 53522 265487 53578 265496
rect 54534 265552 54590 265561
rect 54534 265487 54590 265496
rect 52052 265108 52104 265114
rect 52052 265050 52104 265056
rect 52064 263770 52092 265050
rect 52064 263742 52446 263770
rect 53536 263756 53564 265487
rect 54548 263756 54576 265487
rect 55560 263756 55588 266575
rect 56756 266338 56784 276934
rect 57032 274498 57060 276948
rect 57966 276934 58164 276962
rect 58794 276934 59544 276962
rect 57020 274492 57072 274498
rect 57020 274434 57072 274440
rect 58136 266406 58164 276934
rect 59516 266474 59544 276934
rect 59700 274838 59728 276948
rect 60634 276934 60924 276962
rect 59688 274832 59740 274838
rect 59688 274774 59740 274780
rect 60792 274832 60844 274838
rect 60792 274774 60844 274780
rect 59688 266740 59740 266746
rect 59688 266682 59740 266688
rect 59504 266468 59556 266474
rect 59504 266410 59556 266416
rect 58124 266400 58176 266406
rect 58124 266342 58176 266348
rect 56744 266332 56796 266338
rect 56744 266274 56796 266280
rect 58676 265652 58728 265658
rect 58676 265594 58728 265600
rect 57664 265584 57716 265590
rect 56558 265552 56614 265561
rect 57664 265526 57716 265532
rect 56558 265487 56614 265496
rect 56572 263756 56600 265487
rect 57676 263756 57704 265526
rect 58688 263756 58716 265594
rect 59700 263756 59728 266682
rect 60804 266202 60832 274774
rect 60896 266542 60924 276934
rect 61448 273818 61476 276948
rect 62368 274022 62396 276948
rect 62356 274016 62408 274022
rect 62356 273958 62408 273964
rect 63288 273886 63316 276948
rect 63644 274016 63696 274022
rect 63644 273958 63696 273964
rect 61620 273880 61672 273886
rect 61620 273822 61672 273828
rect 63276 273880 63328 273886
rect 63276 273822 63328 273828
rect 61436 273812 61488 273818
rect 61436 273754 61488 273760
rect 60884 266536 60936 266542
rect 60884 266478 60936 266484
rect 60792 266196 60844 266202
rect 60792 266138 60844 266144
rect 60700 265856 60752 265862
rect 60700 265798 60752 265804
rect 60712 263756 60740 265798
rect 61632 265590 61660 273822
rect 62264 273812 62316 273818
rect 62264 273754 62316 273760
rect 63000 273812 63052 273818
rect 63000 273754 63052 273760
rect 62276 266610 62304 273754
rect 62264 266604 62316 266610
rect 62264 266546 62316 266552
rect 62816 265788 62868 265794
rect 62816 265730 62868 265736
rect 61804 265720 61856 265726
rect 61804 265662 61856 265668
rect 61620 265584 61672 265590
rect 61620 265526 61672 265532
rect 61816 263756 61844 265662
rect 62828 263756 62856 265730
rect 63012 265658 63040 273754
rect 63656 266678 63684 273958
rect 64116 273818 64144 276948
rect 64760 276934 65050 276962
rect 64760 276606 64788 276934
rect 64196 276600 64248 276606
rect 64196 276542 64248 276548
rect 64748 276600 64800 276606
rect 64748 276542 64800 276548
rect 64104 273812 64156 273818
rect 64104 273754 64156 273760
rect 64208 271794 64236 276542
rect 65956 273886 65984 276948
rect 64380 273880 64432 273886
rect 64380 273822 64432 273828
rect 65944 273880 65996 273886
rect 65944 273822 65996 273828
rect 63840 271766 64236 271794
rect 63840 266746 63868 271766
rect 63828 266740 63880 266746
rect 63828 266682 63880 266688
rect 63644 266672 63696 266678
rect 63644 266614 63696 266620
rect 63828 266060 63880 266066
rect 63828 266002 63880 266008
rect 63000 265652 63052 265658
rect 63000 265594 63052 265600
rect 63840 263756 63868 266002
rect 64392 265862 64420 273822
rect 66784 273818 66812 276948
rect 65760 273812 65812 273818
rect 65760 273754 65812 273760
rect 66772 273812 66824 273818
rect 66772 273754 66824 273760
rect 64840 266876 64892 266882
rect 64840 266818 64892 266824
rect 64380 265856 64432 265862
rect 64380 265798 64432 265804
rect 64852 263756 64880 266818
rect 65772 265726 65800 273754
rect 67152 271794 67180 277070
rect 66508 271766 67180 271794
rect 67980 276934 68638 276962
rect 66508 265794 66536 271766
rect 67980 266490 68008 276934
rect 68060 274492 68112 274498
rect 68060 274434 68112 274440
rect 67888 266462 68008 266490
rect 66956 266264 67008 266270
rect 66956 266206 67008 266212
rect 66496 265788 66548 265794
rect 66496 265730 66548 265736
rect 65760 265720 65812 265726
rect 65760 265662 65812 265668
rect 65944 265584 65996 265590
rect 65944 265526 65996 265532
rect 65956 263756 65984 265526
rect 66968 263756 66996 266206
rect 67888 266066 67916 266462
rect 67968 266332 68020 266338
rect 67968 266274 68020 266280
rect 67876 266060 67928 266066
rect 67876 266002 67928 266008
rect 67980 263756 68008 266274
rect 68072 263634 68100 274434
rect 69452 273818 69480 276948
rect 68520 273812 68572 273818
rect 68520 273754 68572 273760
rect 69440 273812 69492 273818
rect 69440 273754 69492 273760
rect 68532 266882 68560 273754
rect 69636 271794 69664 277070
rect 69268 271766 69664 271794
rect 68520 266876 68572 266882
rect 68520 266818 68572 266824
rect 69268 265590 69296 271766
rect 73120 266536 73172 266542
rect 73120 266478 73172 266484
rect 71096 266468 71148 266474
rect 71096 266410 71148 266416
rect 70084 266400 70136 266406
rect 70084 266342 70136 266348
rect 69256 265584 69308 265590
rect 69256 265526 69308 265532
rect 70096 263756 70124 266342
rect 71108 263756 71136 266410
rect 72108 266196 72160 266202
rect 72108 266138 72160 266144
rect 72120 263756 72148 266138
rect 73132 263756 73160 266478
rect 74052 264434 74080 278135
rect 74236 271681 74264 296903
rect 75892 293033 75920 334342
rect 75984 334338 76012 334478
rect 75972 334332 76024 334338
rect 75972 334274 76024 334280
rect 75984 296977 76012 334274
rect 76076 327606 76104 334478
rect 76064 327600 76116 327606
rect 76064 327542 76116 327548
rect 76076 326382 76104 327542
rect 76064 326376 76116 326382
rect 76064 326318 76116 326324
rect 76156 312504 76208 312510
rect 76156 312446 76208 312452
rect 75970 296968 76026 296977
rect 75970 296903 76026 296912
rect 75878 293024 75934 293033
rect 75878 292959 75934 292968
rect 74222 271672 74278 271681
rect 74222 271607 74278 271616
rect 74236 271137 74264 271607
rect 74222 271128 74278 271137
rect 74222 271063 74278 271072
rect 75236 266672 75288 266678
rect 75236 266614 75288 266620
rect 74224 266604 74276 266610
rect 74224 266546 74276 266552
rect 74040 264428 74092 264434
rect 74040 264370 74092 264376
rect 74236 263756 74264 266546
rect 75248 263756 75276 266614
rect 76168 263770 76196 312446
rect 76168 263742 76274 263770
rect 68072 263606 69006 263634
rect 73946 263512 74002 263521
rect 73946 263447 73948 263456
rect 74000 263447 74002 263456
rect 73948 263418 74000 263424
rect 49200 262728 49252 262734
rect 49198 262696 49200 262705
rect 49252 262696 49254 262705
rect 49198 262631 49254 262640
rect 47082 252904 47138 252913
rect 47082 252839 47138 252848
rect 46438 249776 46494 249785
rect 46438 249711 46494 249720
rect 47082 237400 47138 237409
rect 47082 237335 47138 237344
rect 47096 230978 47124 237335
rect 55744 235998 56586 236026
rect 48568 235862 49410 235890
rect 49948 235862 50422 235890
rect 51328 235862 51434 235890
rect 51512 235862 52446 235890
rect 47084 230972 47136 230978
rect 47084 230914 47136 230920
rect 13042 229583 13044 229592
rect 13096 229583 13098 229592
rect 16080 229612 16132 229618
rect 13044 229554 13096 229560
rect 16080 229554 16132 229560
rect 22244 229612 22296 229618
rect 22244 229554 22296 229560
rect 47084 228388 47136 228394
rect 47084 228330 47136 228336
rect 34020 228320 34072 228326
rect 34020 228262 34072 228268
rect 34032 221730 34060 228262
rect 34572 226892 34624 226898
rect 34572 226834 34624 226840
rect 34584 221798 34612 226834
rect 38528 222064 38580 222070
rect 38528 222006 38580 222012
rect 34572 221792 34624 221798
rect 34572 221734 34624 221740
rect 34940 221792 34992 221798
rect 38540 221769 38568 222006
rect 34940 221734 34992 221740
rect 38526 221760 38582 221769
rect 34020 221724 34072 221730
rect 34020 221666 34072 221672
rect 34756 221724 34808 221730
rect 34756 221666 34808 221672
rect 34664 220568 34716 220574
rect 34664 220510 34716 220516
rect 16170 219992 16226 220001
rect 16170 219927 16226 219936
rect 13318 216184 13374 216193
rect 13318 216119 13374 216128
rect 13332 189634 13360 216119
rect 16078 214552 16134 214561
rect 16078 214487 16134 214496
rect 13962 202856 14018 202865
rect 13962 202791 14018 202800
rect 13976 202078 14004 202791
rect 13964 202072 14016 202078
rect 13964 202014 14016 202020
rect 13412 199352 13464 199358
rect 13412 199294 13464 199300
rect 13320 189628 13372 189634
rect 13320 189570 13372 189576
rect 13320 189424 13372 189430
rect 13318 189392 13320 189401
rect 13372 189392 13374 189401
rect 13318 189327 13374 189336
rect 13424 176073 13452 199294
rect 13504 189628 13556 189634
rect 13504 189570 13556 189576
rect 13516 185486 13544 189570
rect 13504 185480 13556 185486
rect 13504 185422 13556 185428
rect 13410 176064 13466 176073
rect 13410 175999 13466 176008
rect 12860 163244 12912 163250
rect 12860 163186 12912 163192
rect 12872 162745 12900 163186
rect 12858 162736 12914 162745
rect 12858 162671 12914 162680
rect 12860 149372 12912 149378
rect 12860 149314 12912 149320
rect 12872 149281 12900 149314
rect 12858 149272 12914 149281
rect 12858 149207 12914 149216
rect 16092 137138 16120 214487
rect 12860 137132 12912 137138
rect 12860 137074 12912 137080
rect 16080 137132 16132 137138
rect 16080 137074 16132 137080
rect 12872 135953 12900 137074
rect 12858 135944 12914 135953
rect 12858 135879 12914 135888
rect 16078 126152 16134 126161
rect 16078 126087 16134 126096
rect 12676 123328 12728 123334
rect 12676 123270 12728 123276
rect 12688 122625 12716 123270
rect 12674 122616 12730 122625
rect 12674 122551 12730 122560
rect 13410 109152 13466 109161
rect 13410 109087 13466 109096
rect 13320 105512 13372 105518
rect 13320 105454 13372 105460
rect 13136 95856 13188 95862
rect 13134 95824 13136 95833
rect 13188 95824 13190 95833
rect 13134 95759 13190 95768
rect 13332 69041 13360 105454
rect 13424 91646 13452 109087
rect 13504 99936 13556 99942
rect 13504 99878 13556 99884
rect 13412 91640 13464 91646
rect 13412 91582 13464 91588
rect 13516 82369 13544 99878
rect 13502 82360 13558 82369
rect 13502 82295 13558 82304
rect 13318 69032 13374 69041
rect 13318 68967 13374 68976
rect 13136 55736 13188 55742
rect 13134 55704 13136 55713
rect 13188 55704 13190 55713
rect 13134 55639 13190 55648
rect 12860 42612 12912 42618
rect 12860 42554 12912 42560
rect 12872 42249 12900 42554
rect 12858 42240 12914 42249
rect 12858 42175 12914 42184
rect 12676 29488 12728 29494
rect 12676 29430 12728 29436
rect 12688 28921 12716 29430
rect 12674 28912 12730 28921
rect 12674 28847 12730 28856
rect 16092 15622 16120 126087
rect 16184 123334 16212 219927
rect 17550 209656 17606 209665
rect 17550 209591 17606 209600
rect 17564 208985 17592 209591
rect 16262 208976 16318 208985
rect 16262 208911 16318 208920
rect 17550 208976 17606 208985
rect 17550 208911 17606 208920
rect 16276 149378 16304 208911
rect 34676 206922 34704 220510
rect 34768 220506 34796 221666
rect 34952 220574 34980 221734
rect 38526 221695 38582 221704
rect 34940 220568 34992 220574
rect 34940 220510 34992 220516
rect 34756 220500 34808 220506
rect 34756 220442 34808 220448
rect 38068 219956 38120 219962
rect 38068 219898 38120 219904
rect 38080 219457 38108 219898
rect 38066 219448 38122 219457
rect 38066 219383 38122 219392
rect 38528 217168 38580 217174
rect 38528 217110 38580 217116
rect 38540 216873 38568 217110
rect 38526 216864 38582 216873
rect 38526 216799 38582 216808
rect 38528 214448 38580 214454
rect 38528 214390 38580 214396
rect 38540 214289 38568 214390
rect 38526 214280 38582 214289
rect 38526 214215 38582 214224
rect 34848 213904 34900 213910
rect 34768 213852 34848 213858
rect 34768 213846 34900 213852
rect 34768 213830 34888 213846
rect 34768 211682 34796 213830
rect 34768 211654 34980 211682
rect 34676 206906 34888 206922
rect 34676 206900 34900 206906
rect 34676 206894 34848 206900
rect 34848 206842 34900 206848
rect 16354 204896 16410 204905
rect 16354 204831 16410 204840
rect 16368 163250 16396 204831
rect 34848 204724 34900 204730
rect 34768 204684 34848 204712
rect 16448 202072 16500 202078
rect 16448 202014 16500 202020
rect 16460 189673 16488 202014
rect 17642 199728 17698 199737
rect 17642 199663 17698 199672
rect 17656 199358 17684 199663
rect 17644 199352 17696 199358
rect 17644 199294 17696 199300
rect 17458 195376 17514 195385
rect 17458 195311 17514 195320
rect 16446 189664 16502 189673
rect 16446 189599 16502 189608
rect 17472 189430 17500 195311
rect 34768 195226 34796 204684
rect 34848 204666 34900 204672
rect 34768 195198 34888 195226
rect 34860 189650 34888 195198
rect 34768 189622 34888 189650
rect 17460 189424 17512 189430
rect 17460 189366 17512 189372
rect 34768 189242 34796 189622
rect 34676 189214 34796 189242
rect 17460 185480 17512 185486
rect 17458 185448 17460 185457
rect 17512 185448 17514 185457
rect 17458 185383 17514 185392
rect 34388 183236 34440 183242
rect 34388 183178 34440 183184
rect 21258 182958 21640 182986
rect 23926 182958 24216 182986
rect 26594 182958 26976 182986
rect 29262 182958 29552 182986
rect 21612 181338 21640 182958
rect 21600 181332 21652 181338
rect 21600 181274 21652 181280
rect 24188 180658 24216 182958
rect 26948 180726 26976 182958
rect 29524 180794 29552 182958
rect 31824 182822 31930 182850
rect 31824 180862 31852 182822
rect 34400 181338 34428 183178
rect 34676 183122 34704 189214
rect 34952 183242 34980 211654
rect 38710 211560 38766 211569
rect 38710 211495 38766 211504
rect 38724 210986 38752 211495
rect 38712 210980 38764 210986
rect 38712 210922 38764 210928
rect 38528 209620 38580 209626
rect 38528 209562 38580 209568
rect 38540 209257 38568 209562
rect 38526 209248 38582 209257
rect 38526 209183 38582 209192
rect 38528 206832 38580 206838
rect 38528 206774 38580 206780
rect 38540 206673 38568 206774
rect 38526 206664 38582 206673
rect 38526 206599 38582 206608
rect 38528 204792 38580 204798
rect 38528 204734 38580 204740
rect 38540 204497 38568 204734
rect 38526 204488 38582 204497
rect 38526 204423 38582 204432
rect 38526 201496 38582 201505
rect 38526 201431 38582 201440
rect 38540 201330 38568 201431
rect 38528 201324 38580 201330
rect 38528 201266 38580 201272
rect 38528 199284 38580 199290
rect 38528 199226 38580 199232
rect 38540 199193 38568 199226
rect 38526 199184 38582 199193
rect 38526 199119 38582 199128
rect 38526 196464 38582 196473
rect 38526 196399 38582 196408
rect 38540 195822 38568 196399
rect 38528 195816 38580 195822
rect 38528 195758 38580 195764
rect 38804 195136 38856 195142
rect 38804 195078 38856 195084
rect 38816 194569 38844 195078
rect 38802 194560 38858 194569
rect 38802 194495 38858 194504
rect 38804 191668 38856 191674
rect 38804 191610 38856 191616
rect 38816 191577 38844 191610
rect 38802 191568 38858 191577
rect 38802 191503 38858 191512
rect 38068 189628 38120 189634
rect 38068 189570 38120 189576
rect 38080 189265 38108 189570
rect 38066 189256 38122 189265
rect 38066 189191 38122 189200
rect 38066 186536 38122 186545
rect 38066 186471 38122 186480
rect 38080 186166 38108 186471
rect 38068 186160 38120 186166
rect 38068 186102 38120 186108
rect 38802 184088 38858 184097
rect 38802 184023 38804 184032
rect 38856 184023 38858 184032
rect 38804 183994 38856 184000
rect 34940 183236 34992 183242
rect 34940 183178 34992 183184
rect 34676 183094 34796 183122
rect 34598 182958 34704 182986
rect 34572 182692 34624 182698
rect 34572 182634 34624 182640
rect 34388 181332 34440 181338
rect 34388 181274 34440 181280
rect 31812 180856 31864 180862
rect 31812 180798 31864 180804
rect 34584 180810 34612 182634
rect 34676 180930 34704 182958
rect 34768 182698 34796 183094
rect 34756 182692 34808 182698
rect 34756 182634 34808 182640
rect 34664 180924 34716 180930
rect 34664 180866 34716 180872
rect 46992 180924 47044 180930
rect 46992 180866 47044 180872
rect 45796 180856 45848 180862
rect 29512 180788 29564 180794
rect 34584 180782 34704 180810
rect 45796 180798 45848 180804
rect 29512 180730 29564 180736
rect 26936 180720 26988 180726
rect 26936 180662 26988 180668
rect 24176 180652 24228 180658
rect 24176 180594 24228 180600
rect 16356 163244 16408 163250
rect 16356 163186 16408 163192
rect 16264 149372 16316 149378
rect 16264 149314 16316 149320
rect 16172 123328 16224 123334
rect 16172 123270 16224 123276
rect 16170 120712 16226 120721
rect 16170 120647 16226 120656
rect 16184 29494 16212 120647
rect 16262 115136 16318 115145
rect 16262 115071 16318 115080
rect 16276 42618 16304 115071
rect 16354 111056 16410 111065
rect 16354 110991 16410 111000
rect 16368 55742 16396 110991
rect 18102 106296 18158 106305
rect 18102 106231 18158 106240
rect 18116 105518 18144 106231
rect 18104 105512 18156 105518
rect 18104 105454 18156 105460
rect 17458 101264 17514 101273
rect 17458 101199 17514 101208
rect 17472 99942 17500 101199
rect 17460 99936 17512 99942
rect 17460 99878 17512 99884
rect 18102 96232 18158 96241
rect 18102 96167 18158 96176
rect 18116 95862 18144 96167
rect 18104 95856 18156 95862
rect 18104 95798 18156 95804
rect 18104 91640 18156 91646
rect 18104 91582 18156 91588
rect 18116 91345 18144 91582
rect 18102 91336 18158 91345
rect 18102 91271 18158 91280
rect 21244 87158 21272 88860
rect 23912 87498 23940 88860
rect 23900 87492 23952 87498
rect 23900 87434 23952 87440
rect 21232 87152 21284 87158
rect 21232 87094 21284 87100
rect 26580 87090 26608 88860
rect 29248 87362 29276 88860
rect 29236 87356 29288 87362
rect 29236 87298 29288 87304
rect 31916 87294 31944 88860
rect 31904 87288 31956 87294
rect 31904 87230 31956 87236
rect 34584 87226 34612 88860
rect 34572 87220 34624 87226
rect 34572 87162 34624 87168
rect 34676 87158 34704 180782
rect 45808 175937 45836 180798
rect 46624 180788 46676 180794
rect 46624 180730 46676 180736
rect 46532 180720 46584 180726
rect 46532 180662 46584 180668
rect 46440 180652 46492 180658
rect 46440 180594 46492 180600
rect 45794 175928 45850 175937
rect 45794 175863 45850 175872
rect 46452 155809 46480 180594
rect 46544 158937 46572 180662
rect 46636 162065 46664 180730
rect 46898 176472 46954 176481
rect 46898 176407 46954 176416
rect 46912 175937 46940 176407
rect 46898 175928 46954 175937
rect 46898 175863 46954 175872
rect 46912 165193 46940 175863
rect 47004 168894 47032 180866
rect 46992 168888 47044 168894
rect 46992 168830 47044 168836
rect 46898 165184 46954 165193
rect 46898 165119 46954 165128
rect 46622 162056 46678 162065
rect 46622 161991 46678 162000
rect 46530 158928 46586 158937
rect 46530 158863 46586 158872
rect 46438 155800 46494 155809
rect 46438 155735 46494 155744
rect 47096 143433 47124 228330
rect 48568 186166 48596 235862
rect 49948 191674 49976 235862
rect 50580 222064 50632 222070
rect 50578 222032 50580 222041
rect 50632 222032 50634 222041
rect 50578 221967 50634 221976
rect 51222 200272 51278 200281
rect 51222 200207 51278 200216
rect 51236 199290 51264 200207
rect 51224 199284 51276 199290
rect 51224 199226 51276 199232
rect 51328 195822 51356 235862
rect 51406 215232 51462 215241
rect 51406 215167 51462 215176
rect 51420 214454 51448 215167
rect 51408 214448 51460 214454
rect 51408 214390 51460 214396
rect 51406 210200 51462 210209
rect 51406 210135 51462 210144
rect 51420 209626 51448 210135
rect 51408 209620 51460 209626
rect 51408 209562 51460 209568
rect 51408 206832 51460 206838
rect 51406 206800 51408 206809
rect 51460 206800 51462 206809
rect 51406 206735 51462 206744
rect 51406 205304 51462 205313
rect 51406 205239 51462 205248
rect 51420 204798 51448 205239
rect 51408 204792 51460 204798
rect 51408 204734 51460 204740
rect 51512 201330 51540 235862
rect 53536 232513 53564 235876
rect 54548 232513 54576 235876
rect 55364 233148 55416 233154
rect 55364 233090 55416 233096
rect 53522 232504 53578 232513
rect 53522 232439 53578 232448
rect 54534 232504 54590 232513
rect 54534 232439 54590 232448
rect 55376 222834 55404 233090
rect 55560 232513 55588 235876
rect 55546 232504 55602 232513
rect 55546 232439 55602 232448
rect 55744 228274 55772 235998
rect 56744 233284 56796 233290
rect 56744 233226 56796 233232
rect 55560 228246 55772 228274
rect 55560 226937 55588 228246
rect 55546 226928 55602 226937
rect 55546 226863 55602 226872
rect 56756 225334 56784 233226
rect 57676 232542 57704 235876
rect 58124 233352 58176 233358
rect 58124 233294 58176 233300
rect 57664 232536 57716 232542
rect 57664 232478 57716 232484
rect 56100 225328 56152 225334
rect 56100 225270 56152 225276
rect 56744 225328 56796 225334
rect 56744 225270 56796 225276
rect 55298 222806 55404 222834
rect 56112 222820 56140 225270
rect 57020 224784 57072 224790
rect 57020 224726 57072 224732
rect 57032 222820 57060 224726
rect 58136 222834 58164 233294
rect 58688 232678 58716 235876
rect 59504 232944 59556 232950
rect 59504 232886 59556 232892
rect 58676 232672 58728 232678
rect 58676 232614 58728 232620
rect 59516 225062 59544 232886
rect 59700 232610 59728 235876
rect 59688 232604 59740 232610
rect 59688 232546 59740 232552
rect 60712 232474 60740 235876
rect 61816 233630 61844 235876
rect 61804 233624 61856 233630
rect 61804 233566 61856 233572
rect 62828 233562 62856 235876
rect 63644 233760 63696 233766
rect 63644 233702 63696 233708
rect 62816 233556 62868 233562
rect 62816 233498 62868 233504
rect 62264 233216 62316 233222
rect 62264 233158 62316 233164
rect 60792 233080 60844 233086
rect 60792 233022 60844 233028
rect 60700 232468 60752 232474
rect 60700 232410 60752 232416
rect 59688 225328 59740 225334
rect 59688 225270 59740 225276
rect 58768 225056 58820 225062
rect 58768 224998 58820 225004
rect 59504 225056 59556 225062
rect 59504 224998 59556 225004
rect 57966 222806 58164 222834
rect 58780 222820 58808 224998
rect 59700 222820 59728 225270
rect 60804 222834 60832 233022
rect 60884 232876 60936 232882
rect 60884 232818 60936 232824
rect 60896 225334 60924 232818
rect 61620 232536 61672 232542
rect 61620 232478 61672 232484
rect 60884 225328 60936 225334
rect 60884 225270 60936 225276
rect 61436 225328 61488 225334
rect 61436 225270 61488 225276
rect 60634 222806 60832 222834
rect 61448 222820 61476 225270
rect 61632 224246 61660 232478
rect 62276 225334 62304 233158
rect 63092 232672 63144 232678
rect 63092 232614 63144 232620
rect 63000 232468 63052 232474
rect 63000 232410 63052 232416
rect 63012 225402 63040 232410
rect 63000 225396 63052 225402
rect 63000 225338 63052 225344
rect 62264 225328 62316 225334
rect 62264 225270 62316 225276
rect 62356 225328 62408 225334
rect 62356 225270 62408 225276
rect 61620 224240 61672 224246
rect 61620 224182 61672 224188
rect 62368 222820 62396 225270
rect 63104 225130 63132 232614
rect 63184 232604 63236 232610
rect 63184 232546 63236 232552
rect 63092 225124 63144 225130
rect 63092 225066 63144 225072
rect 63196 224314 63224 232546
rect 63656 225334 63684 233702
rect 63840 233426 63868 235876
rect 64852 233494 64880 235876
rect 65760 233624 65812 233630
rect 65760 233566 65812 233572
rect 64840 233488 64892 233494
rect 64840 233430 64892 233436
rect 63828 233420 63880 233426
rect 63828 233362 63880 233368
rect 65772 225334 65800 233566
rect 65852 233556 65904 233562
rect 65852 233498 65904 233504
rect 63644 225328 63696 225334
rect 63644 225270 63696 225276
rect 65760 225328 65812 225334
rect 65760 225270 65812 225276
rect 65864 225198 65892 233498
rect 65956 232542 65984 235876
rect 66968 233154 66996 235876
rect 67140 233488 67192 233494
rect 67140 233430 67192 233436
rect 66956 233148 67008 233154
rect 66956 233090 67008 233096
rect 65944 232536 65996 232542
rect 65944 232478 65996 232484
rect 67152 225402 67180 233430
rect 67232 233420 67284 233426
rect 67232 233362 67284 233368
rect 65944 225396 65996 225402
rect 65944 225338 65996 225344
rect 67140 225396 67192 225402
rect 67140 225338 67192 225344
rect 65852 225192 65904 225198
rect 65852 225134 65904 225140
rect 64104 225124 64156 225130
rect 64104 225066 64156 225072
rect 63184 224308 63236 224314
rect 63184 224250 63236 224256
rect 63276 224240 63328 224246
rect 63276 224182 63328 224188
rect 63288 222820 63316 224182
rect 64116 222820 64144 225066
rect 65024 224308 65076 224314
rect 65024 224250 65076 224256
rect 65036 222820 65064 224250
rect 65956 222820 65984 225338
rect 66772 225328 66824 225334
rect 66772 225270 66824 225276
rect 66784 222820 66812 225270
rect 67244 224314 67272 233362
rect 67980 233290 68008 235876
rect 67968 233284 68020 233290
rect 67968 233226 68020 233232
rect 68520 232536 68572 232542
rect 68520 232478 68572 232484
rect 67324 232468 67376 232474
rect 67324 232410 67376 232416
rect 67336 224790 67364 232410
rect 68532 225334 68560 232478
rect 68992 232474 69020 235876
rect 70096 233358 70124 235876
rect 70084 233352 70136 233358
rect 70084 233294 70136 233300
rect 71108 232950 71136 235876
rect 71096 232944 71148 232950
rect 71096 232886 71148 232892
rect 72120 232882 72148 235876
rect 73132 233086 73160 235876
rect 74130 233728 74186 233737
rect 74130 233663 74186 233672
rect 74144 233154 74172 233663
rect 74236 233222 74264 235876
rect 74682 235088 74738 235097
rect 74682 235023 74738 235032
rect 74224 233216 74276 233222
rect 74224 233158 74276 233164
rect 74132 233148 74184 233154
rect 74132 233090 74184 233096
rect 73120 233080 73172 233086
rect 73120 233022 73172 233028
rect 72108 232876 72160 232882
rect 72108 232818 72160 232824
rect 68980 232468 69032 232474
rect 68980 232410 69032 232416
rect 74040 228456 74092 228462
rect 74040 228398 74092 228404
rect 69440 225396 69492 225402
rect 69440 225338 69492 225344
rect 68520 225328 68572 225334
rect 68520 225270 68572 225276
rect 67692 225192 67744 225198
rect 67692 225134 67744 225140
rect 67324 224784 67376 224790
rect 67324 224726 67376 224732
rect 67232 224308 67284 224314
rect 67232 224250 67284 224256
rect 67704 222820 67732 225134
rect 68612 224308 68664 224314
rect 68612 224250 68664 224256
rect 68624 222820 68652 224250
rect 69452 222820 69480 225338
rect 70360 225328 70412 225334
rect 70360 225270 70412 225276
rect 70372 222820 70400 225270
rect 73946 224344 74002 224353
rect 73946 224279 74002 224288
rect 73960 223945 73988 224279
rect 73946 223936 74002 223945
rect 73946 223871 74002 223880
rect 53246 221352 53302 221361
rect 53246 221287 53302 221296
rect 52050 220264 52106 220273
rect 52050 220199 52106 220208
rect 52064 219962 52092 220199
rect 52052 219956 52104 219962
rect 52052 219898 52104 219904
rect 53260 217174 53288 221287
rect 53248 217168 53300 217174
rect 53248 217110 53300 217116
rect 54074 211016 54130 211025
rect 54074 210951 54076 210960
rect 54128 210951 54130 210960
rect 54076 210922 54128 210928
rect 70818 209520 70874 209529
rect 70818 209455 70874 209464
rect 70832 204769 70860 209455
rect 73854 205032 73910 205041
rect 73854 204967 73910 204976
rect 73868 204769 73896 204967
rect 70818 204760 70874 204769
rect 70818 204695 70874 204704
rect 73854 204760 73910 204769
rect 73854 204695 73910 204704
rect 51500 201324 51552 201330
rect 51500 201266 51552 201272
rect 51316 195816 51368 195822
rect 51316 195758 51368 195764
rect 51328 195362 51356 195758
rect 51236 195334 51356 195362
rect 51236 195090 51264 195334
rect 51314 195240 51370 195249
rect 51314 195175 51316 195184
rect 51368 195175 51370 195184
rect 51316 195146 51368 195152
rect 51236 195062 51356 195090
rect 49936 191668 49988 191674
rect 49936 191610 49988 191616
rect 48556 186160 48608 186166
rect 48556 186102 48608 186108
rect 48568 169930 48596 186102
rect 48568 169902 48964 169930
rect 48936 169658 48964 169902
rect 49948 169794 49976 191610
rect 51222 190208 51278 190217
rect 51222 190143 51278 190152
rect 51236 189634 51264 190143
rect 51224 189628 51276 189634
rect 51224 189570 51276 189576
rect 51328 169794 51356 195062
rect 51406 185312 51462 185321
rect 51406 185247 51462 185256
rect 51420 184058 51448 185247
rect 51408 184052 51460 184058
rect 51408 183994 51460 184000
rect 51512 179858 51540 201266
rect 73946 185584 74002 185593
rect 73946 185519 74002 185528
rect 73960 185457 73988 185519
rect 73946 185448 74002 185457
rect 73946 185383 74002 185392
rect 74052 185049 74080 228398
rect 74144 206537 74172 233090
rect 74222 220400 74278 220409
rect 74222 220335 74278 220344
rect 74130 206528 74186 206537
rect 74130 206463 74186 206472
rect 74144 204905 74172 206463
rect 74130 204896 74186 204905
rect 74130 204831 74186 204840
rect 74130 203536 74186 203545
rect 74130 203471 74186 203480
rect 74144 188041 74172 203471
rect 74236 203370 74264 220335
rect 74696 210209 74724 235023
rect 75248 233562 75276 235876
rect 76168 235862 76274 235890
rect 76064 235120 76116 235126
rect 76062 235088 76064 235097
rect 76116 235088 76118 235097
rect 76062 235023 76118 235032
rect 75236 233556 75288 233562
rect 75236 233498 75288 233504
rect 76168 219554 76196 235862
rect 76812 230910 76840 359706
rect 76892 357452 76944 357458
rect 76892 357394 76944 357400
rect 76904 331754 76932 357394
rect 76996 334338 77024 359774
rect 80204 357928 80256 357934
rect 80204 357870 80256 357876
rect 80216 357633 80244 357870
rect 80202 357624 80258 357633
rect 80202 357559 80258 357568
rect 80204 356568 80256 356574
rect 80204 356510 80256 356516
rect 80216 356409 80244 356510
rect 80202 356400 80258 356409
rect 80202 356335 80258 356344
rect 80204 355208 80256 355214
rect 80204 355150 80256 355156
rect 79284 355140 79336 355146
rect 79284 355082 79336 355088
rect 79296 354641 79324 355082
rect 80216 355049 80244 355150
rect 80202 355040 80258 355049
rect 80202 354975 80258 354984
rect 79282 354632 79338 354641
rect 79282 354567 79338 354576
rect 78916 353848 78968 353854
rect 78916 353790 78968 353796
rect 78928 353417 78956 353790
rect 78914 353408 78970 353417
rect 78914 353343 78970 353352
rect 80204 352420 80256 352426
rect 80204 352362 80256 352368
rect 80216 352193 80244 352362
rect 80202 352184 80258 352193
rect 80202 352119 80258 352128
rect 87194 351368 87250 351377
rect 87194 351303 87250 351312
rect 79100 351060 79152 351066
rect 79100 351002 79152 351008
rect 79112 350425 79140 351002
rect 80202 350688 80258 350697
rect 80202 350623 80258 350632
rect 79098 350416 79154 350425
rect 80216 350386 80244 350623
rect 79098 350351 79154 350360
rect 80204 350380 80256 350386
rect 80204 350322 80256 350328
rect 87208 349706 87236 351303
rect 89876 351066 89904 367662
rect 90060 367658 90088 370924
rect 92544 367726 92572 370924
rect 92532 367720 92584 367726
rect 92532 367662 92584 367668
rect 95028 367658 95056 370924
rect 90048 367652 90100 367658
rect 90048 367594 90100 367600
rect 91428 367652 91480 367658
rect 91428 367594 91480 367600
rect 95016 367652 95068 367658
rect 95016 367594 95068 367600
rect 96856 367652 96908 367658
rect 96856 367594 96908 367600
rect 91440 351898 91468 367594
rect 91440 351870 92112 351898
rect 92084 351762 92112 351870
rect 92084 351734 92420 351762
rect 96868 351626 96896 367594
rect 97512 367289 97540 370924
rect 99996 367658 100024 370924
rect 102388 370910 102494 370938
rect 99984 367652 100036 367658
rect 99984 367594 100036 367600
rect 100904 367652 100956 367658
rect 100904 367594 100956 367600
rect 97498 367280 97554 367289
rect 97498 367215 97554 367224
rect 100916 355078 100944 367594
rect 102388 358834 102416 370910
rect 105056 367658 105084 370924
rect 106528 370910 107554 370938
rect 105044 367652 105096 367658
rect 105044 367594 105096 367600
rect 102388 358806 102692 358834
rect 100904 355072 100956 355078
rect 100904 355014 100956 355020
rect 102376 355072 102428 355078
rect 102376 355014 102428 355020
rect 97314 352048 97370 352057
rect 97314 351983 97316 351992
rect 97368 351983 97370 351992
rect 97316 351954 97368 351960
rect 102388 351762 102416 355014
rect 102664 352426 102692 358806
rect 106528 353854 106556 370910
rect 110024 367658 110052 370924
rect 112140 370910 112522 370938
rect 106608 367652 106660 367658
rect 106608 367594 106660 367600
rect 110012 367652 110064 367658
rect 110012 367594 110064 367600
rect 112036 367652 112088 367658
rect 112036 367594 112088 367600
rect 106516 353848 106568 353854
rect 106516 353790 106568 353796
rect 102652 352420 102704 352426
rect 102652 352362 102704 352368
rect 102356 351734 102416 351762
rect 106620 351626 106648 367594
rect 112048 351762 112076 367594
rect 112140 355146 112168 370910
rect 114992 367658 115020 370924
rect 114980 367652 115032 367658
rect 114980 367594 115032 367600
rect 116176 367652 116228 367658
rect 116176 367594 116228 367600
rect 116188 363510 116216 367594
rect 116176 363504 116228 363510
rect 116176 363446 116228 363452
rect 117004 363504 117056 363510
rect 117004 363446 117056 363452
rect 112128 355140 112180 355146
rect 112128 355082 112180 355088
rect 117016 351762 117044 363446
rect 117568 355214 117596 370924
rect 120052 367658 120080 370924
rect 121800 370910 122550 370938
rect 125034 370910 125784 370938
rect 120040 367652 120092 367658
rect 120040 367594 120092 367600
rect 121696 367652 121748 367658
rect 121696 367594 121748 367600
rect 117556 355208 117608 355214
rect 117556 355150 117608 355156
rect 121708 351898 121736 367594
rect 121800 356574 121828 370910
rect 121788 356568 121840 356574
rect 121788 356510 121840 356516
rect 125756 355078 125784 370910
rect 127228 370910 127518 370938
rect 127228 357934 127256 370910
rect 127872 366230 127900 388538
rect 185372 386700 185400 388538
rect 190328 388528 190380 388534
rect 190328 388470 190380 388476
rect 190340 386700 190368 388470
rect 194848 386714 194876 389218
rect 205324 389208 205376 389214
rect 205324 389150 205376 389156
rect 200356 388936 200408 388942
rect 200356 388878 200408 388884
rect 194848 386686 195322 386714
rect 200368 386700 200396 388878
rect 205336 386700 205364 389150
rect 212788 389078 212816 393774
rect 210292 389072 210344 389078
rect 210292 389014 210344 389020
rect 212776 389072 212828 389078
rect 212776 389014 212828 389020
rect 210304 386700 210332 389014
rect 228600 388596 228652 388602
rect 228600 388538 228652 388544
rect 215352 388460 215404 388466
rect 215352 388402 215404 388408
rect 220320 388460 220372 388466
rect 220320 388402 220372 388408
rect 215364 386700 215392 388402
rect 220332 386700 220360 388402
rect 131354 384824 131410 384833
rect 131354 384759 131410 384768
rect 225194 384824 225250 384833
rect 225194 384759 225250 384768
rect 127860 366224 127912 366230
rect 127860 366166 127912 366172
rect 127216 357928 127268 357934
rect 127216 357870 127268 357876
rect 125744 355072 125796 355078
rect 125744 355014 125796 355020
rect 127216 355072 127268 355078
rect 127216 355014 127268 355020
rect 121708 351870 121920 351898
rect 112048 351734 112384 351762
rect 117016 351734 117352 351762
rect 121892 351626 121920 351870
rect 127228 351762 127256 355014
rect 127228 351734 127380 351762
rect 96868 351598 97388 351626
rect 106620 351598 107416 351626
rect 121892 351598 122412 351626
rect 89864 351060 89916 351066
rect 89864 351002 89916 351008
rect 87470 350416 87526 350425
rect 87470 350351 87526 350360
rect 80204 349700 80256 349706
rect 80204 349642 80256 349648
rect 87196 349700 87248 349706
rect 87196 349642 87248 349648
rect 80216 349337 80244 349642
rect 87286 349600 87342 349609
rect 87286 349535 87342 349544
rect 80202 349328 80258 349337
rect 80202 349263 80258 349272
rect 80204 348272 80256 348278
rect 80204 348214 80256 348220
rect 80216 348113 80244 348214
rect 80202 348104 80258 348113
rect 80202 348039 80258 348048
rect 87102 347832 87158 347841
rect 87102 347767 87158 347776
rect 80204 346912 80256 346918
rect 80204 346854 80256 346860
rect 79284 346844 79336 346850
rect 79284 346786 79336 346792
rect 79296 346345 79324 346786
rect 80216 346753 80244 346854
rect 80202 346744 80258 346753
rect 80202 346679 80258 346688
rect 79282 346336 79338 346345
rect 79282 346271 79338 346280
rect 79652 345620 79704 345626
rect 79652 345562 79704 345568
rect 79664 344033 79692 345562
rect 80202 344840 80258 344849
rect 87116 344810 87144 347767
rect 87300 346918 87328 349535
rect 87378 348648 87434 348657
rect 87378 348583 87434 348592
rect 87288 346912 87340 346918
rect 87194 346880 87250 346889
rect 87288 346854 87340 346860
rect 87392 346850 87420 348583
rect 87484 348278 87512 350351
rect 87472 348272 87524 348278
rect 87472 348214 87524 348220
rect 87194 346815 87250 346824
rect 87380 346844 87432 346850
rect 87208 345626 87236 346815
rect 87380 346786 87432 346792
rect 88114 346064 88170 346073
rect 88114 345999 88170 346008
rect 87196 345620 87248 345626
rect 87196 345562 87248 345568
rect 87378 345112 87434 345121
rect 87378 345047 87434 345056
rect 80202 344775 80204 344784
rect 80256 344775 80258 344784
rect 87104 344804 87156 344810
rect 80204 344746 80256 344752
rect 87104 344746 87156 344752
rect 87392 344674 87420 345047
rect 85816 344668 85868 344674
rect 85816 344610 85868 344616
rect 87380 344668 87432 344674
rect 87380 344610 87432 344616
rect 79650 344024 79706 344033
rect 79650 343959 79706 343968
rect 80202 342800 80258 342809
rect 80202 342735 80204 342744
rect 80256 342735 80258 342744
rect 80204 342706 80256 342712
rect 85828 342158 85856 344610
rect 87286 343344 87342 343353
rect 87286 343279 87342 343288
rect 80204 342152 80256 342158
rect 80204 342094 80256 342100
rect 85816 342152 85868 342158
rect 85816 342094 85868 342100
rect 80216 341857 80244 342094
rect 80202 341848 80258 341857
rect 80202 341783 80258 341792
rect 87194 341576 87250 341585
rect 87194 341511 87250 341520
rect 80204 341404 80256 341410
rect 80204 341346 80256 341352
rect 80216 341041 80244 341346
rect 80202 341032 80258 341041
rect 80202 340967 80258 340976
rect 80204 340044 80256 340050
rect 80204 339986 80256 339992
rect 80216 339817 80244 339986
rect 80202 339808 80258 339817
rect 80202 339743 80258 339752
rect 85080 338684 85132 338690
rect 85080 338626 85132 338632
rect 80204 338616 80256 338622
rect 80204 338558 80256 338564
rect 80112 338548 80164 338554
rect 80112 338490 80164 338496
rect 80124 338049 80152 338490
rect 80216 338457 80244 338558
rect 80202 338448 80258 338457
rect 80202 338383 80258 338392
rect 80110 338040 80166 338049
rect 80110 337975 80166 337984
rect 79836 337256 79888 337262
rect 79836 337198 79888 337204
rect 79848 336825 79876 337198
rect 79834 336816 79890 336825
rect 79834 336751 79890 336760
rect 80204 335896 80256 335902
rect 80204 335838 80256 335844
rect 80216 335737 80244 335838
rect 80202 335728 80258 335737
rect 80202 335663 80258 335672
rect 76984 334332 77036 334338
rect 76984 334274 77036 334280
rect 80110 334096 80166 334105
rect 80110 334031 80166 334040
rect 80204 334060 80256 334066
rect 80124 333930 80152 334031
rect 80204 334002 80256 334008
rect 80112 333924 80164 333930
rect 80112 333866 80164 333872
rect 80216 333697 80244 334002
rect 85092 333930 85120 338626
rect 87208 338554 87236 341511
rect 87300 340050 87328 343279
rect 88128 342770 88156 345999
rect 88482 344296 88538 344305
rect 88482 344231 88538 344240
rect 88116 342764 88168 342770
rect 88116 342706 88168 342712
rect 87562 342392 87618 342401
rect 87562 342327 87618 342336
rect 87378 340624 87434 340633
rect 87378 340559 87434 340568
rect 87288 340044 87340 340050
rect 87288 339986 87340 339992
rect 87286 339808 87342 339817
rect 87286 339743 87342 339752
rect 87196 338548 87248 338554
rect 87196 338490 87248 338496
rect 87194 338040 87250 338049
rect 87194 337975 87250 337984
rect 87208 337330 87236 337975
rect 85172 337324 85224 337330
rect 85172 337266 85224 337272
rect 87196 337324 87248 337330
rect 87196 337266 87248 337272
rect 85184 334066 85212 337266
rect 87194 336272 87250 336281
rect 87194 336207 87250 336216
rect 87208 335970 87236 336207
rect 85816 335964 85868 335970
rect 85816 335906 85868 335912
rect 87196 335964 87248 335970
rect 87196 335906 87248 335912
rect 85172 334060 85224 334066
rect 85172 334002 85224 334008
rect 85080 333924 85132 333930
rect 85080 333866 85132 333872
rect 80202 333688 80258 333697
rect 80202 333623 80258 333632
rect 80204 333108 80256 333114
rect 80204 333050 80256 333056
rect 80216 332745 80244 333050
rect 80202 332736 80258 332745
rect 80202 332671 80258 332680
rect 76892 331748 76944 331754
rect 76892 331690 76944 331696
rect 76904 305681 76932 331690
rect 80202 330968 80258 330977
rect 80202 330903 80258 330912
rect 80216 330802 80244 330903
rect 85828 330802 85856 335906
rect 87300 335902 87328 339743
rect 87392 337262 87420 340559
rect 87470 338856 87526 338865
rect 87470 338791 87526 338800
rect 87484 338690 87512 338791
rect 87472 338684 87524 338690
rect 87472 338626 87524 338632
rect 87576 338622 87604 342327
rect 88496 341410 88524 344231
rect 88484 341404 88536 341410
rect 88484 341346 88536 341352
rect 87564 338616 87616 338622
rect 87564 338558 87616 338564
rect 87380 337256 87432 337262
rect 87380 337198 87432 337204
rect 87562 337088 87618 337097
rect 87562 337023 87618 337032
rect 87288 335896 87340 335902
rect 87288 335838 87340 335844
rect 87576 333114 87604 337023
rect 91592 335822 91928 335850
rect 94904 335822 95240 335850
rect 98216 335822 98276 335850
rect 91244 333924 91296 333930
rect 91244 333866 91296 333872
rect 87564 333108 87616 333114
rect 87564 333050 87616 333056
rect 80204 330796 80256 330802
rect 80204 330738 80256 330744
rect 85816 330796 85868 330802
rect 85816 330738 85868 330744
rect 82318 329744 82374 329753
rect 82318 329679 82374 329688
rect 82332 329034 82360 329679
rect 82320 329028 82372 329034
rect 82320 328970 82372 328976
rect 76984 326308 77036 326314
rect 76984 326250 77036 326256
rect 76996 313598 77024 326250
rect 91256 321706 91284 333866
rect 91900 333794 91928 335822
rect 95212 333833 95240 335822
rect 98248 334338 98276 335822
rect 101008 335822 101528 335850
rect 104872 335822 104932 335850
rect 108244 335822 108304 335850
rect 98236 334332 98288 334338
rect 98236 334274 98288 334280
rect 98248 333862 98276 334274
rect 98236 333856 98288 333862
rect 95198 333824 95254 333833
rect 91888 333788 91940 333794
rect 98236 333798 98288 333804
rect 95198 333759 95254 333768
rect 91888 333730 91940 333736
rect 101008 327606 101036 335822
rect 104872 334406 104900 335822
rect 108276 334474 108304 335822
rect 111404 335822 111556 335850
rect 114808 335822 114868 335850
rect 118212 335822 118272 335850
rect 121248 335822 121584 335850
rect 124560 335822 124896 335850
rect 127872 335822 128208 335850
rect 108264 334468 108316 334474
rect 108264 334410 108316 334416
rect 104860 334400 104912 334406
rect 104860 334342 104912 334348
rect 111404 334338 111432 335822
rect 111392 334332 111444 334338
rect 111392 334274 111444 334280
rect 103664 333992 103716 333998
rect 103664 333934 103716 333940
rect 100996 327600 101048 327606
rect 100996 327542 101048 327548
rect 102284 327600 102336 327606
rect 102284 327542 102336 327548
rect 102296 326926 102324 327542
rect 102284 326920 102336 326926
rect 102284 326862 102336 326868
rect 103676 321706 103704 333934
rect 111404 331618 111432 334274
rect 114808 334270 114836 335822
rect 114796 334264 114848 334270
rect 114796 334206 114848 334212
rect 114808 331686 114836 334206
rect 118212 334202 118240 335822
rect 118200 334196 118252 334202
rect 118200 334138 118252 334144
rect 116084 334060 116136 334066
rect 116084 334002 116136 334008
rect 114796 331680 114848 331686
rect 114796 331622 114848 331628
rect 111392 331612 111444 331618
rect 111392 331554 111444 331560
rect 116096 321706 116124 334002
rect 118212 331754 118240 334138
rect 121248 333930 121276 335822
rect 124560 333998 124588 335822
rect 127872 334066 127900 335822
rect 131368 334202 131396 384759
rect 131446 382104 131502 382113
rect 131446 382039 131502 382048
rect 131460 334270 131488 382039
rect 131538 380200 131594 380209
rect 131538 380135 131594 380144
rect 131552 334338 131580 380135
rect 131630 377480 131686 377489
rect 131630 377415 131686 377424
rect 131644 334474 131672 377415
rect 131722 374760 131778 374769
rect 131722 374695 131778 374704
rect 131632 334468 131684 334474
rect 131632 334410 131684 334416
rect 131540 334332 131592 334338
rect 131540 334274 131592 334280
rect 131448 334264 131500 334270
rect 131448 334206 131500 334212
rect 131356 334196 131408 334202
rect 131356 334138 131408 334144
rect 127860 334060 127912 334066
rect 127860 334002 127912 334008
rect 124548 333992 124600 333998
rect 124548 333934 124600 333940
rect 131368 333930 131396 334138
rect 131460 333998 131488 334206
rect 131552 334134 131580 334274
rect 131540 334128 131592 334134
rect 131540 334070 131592 334076
rect 131644 334066 131672 334410
rect 131736 334406 131764 374695
rect 131814 372176 131870 372185
rect 131814 372111 131870 372120
rect 131828 371806 131856 372111
rect 131816 371800 131868 371806
rect 131816 371742 131868 371748
rect 134760 371800 134812 371806
rect 134760 371742 134812 371748
rect 131814 351368 131870 351377
rect 131814 351303 131870 351312
rect 131828 351134 131856 351303
rect 131816 351128 131868 351134
rect 131816 351070 131868 351076
rect 131814 350416 131870 350425
rect 131814 350351 131870 350360
rect 131828 349774 131856 350351
rect 131816 349768 131868 349774
rect 131816 349710 131868 349716
rect 131906 349600 131962 349609
rect 131906 349535 131962 349544
rect 131814 348648 131870 348657
rect 131814 348583 131870 348592
rect 131828 348346 131856 348583
rect 131920 348414 131948 349535
rect 131908 348408 131960 348414
rect 131908 348350 131960 348356
rect 131816 348340 131868 348346
rect 131816 348282 131868 348288
rect 132182 347832 132238 347841
rect 132182 347767 132238 347776
rect 132196 346986 132224 347767
rect 132184 346980 132236 346986
rect 132184 346922 132236 346928
rect 131906 346880 131962 346889
rect 131906 346815 131962 346824
rect 131814 346064 131870 346073
rect 131814 345999 131870 346008
rect 131828 345694 131856 345999
rect 131816 345688 131868 345694
rect 131816 345630 131868 345636
rect 131920 345626 131948 346815
rect 134116 345688 134168 345694
rect 134116 345630 134168 345636
rect 131908 345620 131960 345626
rect 131908 345562 131960 345568
rect 132366 345112 132422 345121
rect 132366 345047 132422 345056
rect 131814 344296 131870 344305
rect 131814 344231 131816 344240
rect 131868 344231 131870 344240
rect 131816 344202 131868 344208
rect 132380 344198 132408 345047
rect 132368 344192 132420 344198
rect 132368 344134 132420 344140
rect 131814 343344 131870 343353
rect 131814 343279 131870 343288
rect 131828 342838 131856 343279
rect 131816 342832 131868 342838
rect 131816 342774 131868 342780
rect 134128 342770 134156 345630
rect 134116 342764 134168 342770
rect 134116 342706 134168 342712
rect 131906 342392 131962 342401
rect 131906 342327 131962 342336
rect 131814 341576 131870 341585
rect 131920 341546 131948 342327
rect 131814 341511 131870 341520
rect 131908 341540 131960 341546
rect 131828 341478 131856 341511
rect 131908 341482 131960 341488
rect 131816 341472 131868 341478
rect 131816 341414 131868 341420
rect 131814 340624 131870 340633
rect 131814 340559 131870 340568
rect 131828 340118 131856 340559
rect 131816 340112 131868 340118
rect 131816 340054 131868 340060
rect 131906 339808 131962 339817
rect 131906 339743 131962 339752
rect 131814 338856 131870 338865
rect 131814 338791 131870 338800
rect 131828 338758 131856 338791
rect 131816 338752 131868 338758
rect 131816 338694 131868 338700
rect 131920 338690 131948 339743
rect 131908 338684 131960 338690
rect 131908 338626 131960 338632
rect 131814 338040 131870 338049
rect 131814 337975 131870 337984
rect 131828 337330 131856 337975
rect 131816 337324 131868 337330
rect 131816 337266 131868 337272
rect 131906 337088 131962 337097
rect 131906 337023 131962 337032
rect 131814 336272 131870 336281
rect 131814 336207 131870 336216
rect 131828 335970 131856 336207
rect 131920 336038 131948 337023
rect 131908 336032 131960 336038
rect 131908 335974 131960 335980
rect 131816 335964 131868 335970
rect 131816 335906 131868 335912
rect 131724 334400 131776 334406
rect 131724 334342 131776 334348
rect 131736 334202 131764 334342
rect 131724 334196 131776 334202
rect 131724 334138 131776 334144
rect 131632 334060 131684 334066
rect 131632 334002 131684 334008
rect 131448 333992 131500 333998
rect 131448 333934 131500 333940
rect 121236 333924 121288 333930
rect 121236 333866 121288 333872
rect 131356 333924 131408 333930
rect 131356 333866 131408 333872
rect 118200 331748 118252 331754
rect 118200 331690 118252 331696
rect 128504 329232 128556 329238
rect 128504 329174 128556 329180
rect 91086 321678 91284 321706
rect 103506 321678 103704 321706
rect 116018 321678 116124 321706
rect 128516 321692 128544 329174
rect 76984 313592 77036 313598
rect 81676 313592 81728 313598
rect 76984 313534 77036 313540
rect 81674 313560 81676 313569
rect 81728 313560 81730 313569
rect 76996 312510 77024 313534
rect 81674 313495 81730 313504
rect 76984 312504 77036 312510
rect 76984 312446 77036 312452
rect 76890 305672 76946 305681
rect 76890 305607 76946 305616
rect 81676 297204 81728 297210
rect 81676 297146 81728 297152
rect 81688 296841 81716 297146
rect 81674 296832 81730 296841
rect 81674 296767 81730 296776
rect 81676 280680 81728 280686
rect 81676 280622 81728 280628
rect 81688 280249 81716 280622
rect 81674 280240 81730 280249
rect 81674 280175 81730 280184
rect 88404 269670 88432 271916
rect 88392 269664 88444 269670
rect 88392 269606 88444 269612
rect 95488 269602 95516 271916
rect 102664 269602 102692 271916
rect 95476 269596 95528 269602
rect 95476 269538 95528 269544
rect 96764 269596 96816 269602
rect 96764 269538 96816 269544
rect 102652 269596 102704 269602
rect 102652 269538 102704 269544
rect 95568 269052 95620 269058
rect 95568 268994 95620 269000
rect 78916 264088 78968 264094
rect 78916 264030 78968 264036
rect 78928 263657 78956 264030
rect 78914 263648 78970 263657
rect 78914 263583 78970 263592
rect 78914 261744 78970 261753
rect 78914 261679 78970 261688
rect 78928 261442 78956 261679
rect 78916 261436 78968 261442
rect 78916 261378 78968 261384
rect 87196 261436 87248 261442
rect 87196 261378 87248 261384
rect 78914 260384 78970 260393
rect 78914 260319 78970 260328
rect 78928 260082 78956 260319
rect 78916 260076 78968 260082
rect 78916 260018 78968 260024
rect 85080 260076 85132 260082
rect 85080 260018 85132 260024
rect 78914 258888 78970 258897
rect 78914 258823 78970 258832
rect 78928 258722 78956 258823
rect 78916 258716 78968 258722
rect 78916 258658 78968 258664
rect 84436 258716 84488 258722
rect 84436 258658 84488 258664
rect 78914 257528 78970 257537
rect 78914 257463 78970 257472
rect 78928 257362 78956 257463
rect 78916 257356 78968 257362
rect 78916 257298 78968 257304
rect 81676 257356 81728 257362
rect 81676 257298 81728 257304
rect 78914 256168 78970 256177
rect 78914 256103 78970 256112
rect 78928 255934 78956 256103
rect 78916 255928 78968 255934
rect 78916 255870 78968 255876
rect 81688 255866 81716 257298
rect 81768 255928 81820 255934
rect 81768 255870 81820 255876
rect 81676 255860 81728 255866
rect 81676 255802 81728 255808
rect 78914 254672 78970 254681
rect 78914 254607 78970 254616
rect 78928 254506 78956 254607
rect 78916 254500 78968 254506
rect 78916 254442 78968 254448
rect 81780 254438 81808 255870
rect 84448 255798 84476 258658
rect 85092 256886 85120 260018
rect 87208 258081 87236 261378
rect 95580 261374 95608 268994
rect 96776 268990 96804 269538
rect 109748 269058 109776 271916
rect 109736 269052 109788 269058
rect 109736 268994 109788 269000
rect 96764 268984 96816 268990
rect 96764 268926 96816 268932
rect 116924 268582 116952 271916
rect 124008 271794 124036 271916
rect 123272 271766 124036 271794
rect 114796 268576 114848 268582
rect 114796 268518 114848 268524
rect 116912 268576 116964 268582
rect 116912 268518 116964 268524
rect 95568 261368 95620 261374
rect 95568 261310 95620 261316
rect 96212 261368 96264 261374
rect 96212 261310 96264 261316
rect 87194 258072 87250 258081
rect 87194 258007 87250 258016
rect 96224 257786 96252 261310
rect 114808 260490 114836 268518
rect 123272 264094 123300 271766
rect 131184 269398 131212 271916
rect 127768 269392 127820 269398
rect 127768 269334 127820 269340
rect 131172 269392 131224 269398
rect 131172 269334 131224 269340
rect 123260 264088 123312 264094
rect 123260 264030 123312 264036
rect 124364 264088 124416 264094
rect 124364 264030 124416 264036
rect 124376 263482 124404 264030
rect 124364 263476 124416 263482
rect 124364 263418 124416 263424
rect 127780 260626 127808 269334
rect 132000 262796 132052 262802
rect 132000 262738 132052 262744
rect 123536 260620 123588 260626
rect 123536 260562 123588 260568
rect 127768 260620 127820 260626
rect 127768 260562 127820 260568
rect 110196 260484 110248 260490
rect 110196 260426 110248 260432
rect 114796 260484 114848 260490
rect 114796 260426 114848 260432
rect 110208 257786 110236 260426
rect 123548 257786 123576 260562
rect 96224 257758 96560 257786
rect 109900 257758 110236 257786
rect 123240 257758 123576 257786
rect 131354 257392 131410 257401
rect 131354 257327 131410 257336
rect 131368 257294 131396 257327
rect 131356 257288 131408 257294
rect 131356 257230 131408 257236
rect 85080 256880 85132 256886
rect 87196 256880 87248 256886
rect 85080 256822 85132 256828
rect 87194 256848 87196 256857
rect 87248 256848 87250 256857
rect 87194 256783 87250 256792
rect 87196 255860 87248 255866
rect 87196 255802 87248 255808
rect 84436 255792 84488 255798
rect 84436 255734 84488 255740
rect 87208 255361 87236 255802
rect 87288 255792 87340 255798
rect 132012 255746 132040 262738
rect 132092 261436 132144 261442
rect 132092 261378 132144 261384
rect 87288 255734 87340 255740
rect 87300 255633 87328 255734
rect 131828 255718 132040 255746
rect 87286 255624 87342 255633
rect 87286 255559 87342 255568
rect 87194 255352 87250 255361
rect 87194 255287 87250 255296
rect 131354 254672 131410 254681
rect 131354 254607 131356 254616
rect 131408 254607 131410 254616
rect 131356 254578 131408 254584
rect 82688 254500 82740 254506
rect 82688 254442 82740 254448
rect 81768 254432 81820 254438
rect 81768 254374 81820 254380
rect 78914 253312 78970 253321
rect 78914 253247 78970 253256
rect 78928 253146 78956 253247
rect 78916 253140 78968 253146
rect 78916 253082 78968 253088
rect 82700 252942 82728 254442
rect 87196 254432 87248 254438
rect 87194 254400 87196 254409
rect 87248 254400 87250 254409
rect 87194 254335 87250 254344
rect 131354 253856 131410 253865
rect 131354 253791 131410 253800
rect 131368 253214 131396 253791
rect 131356 253208 131408 253214
rect 131356 253150 131408 253156
rect 87288 253004 87340 253010
rect 87288 252946 87340 252952
rect 82688 252936 82740 252942
rect 87196 252936 87248 252942
rect 82688 252878 82740 252884
rect 87194 252904 87196 252913
rect 87248 252904 87250 252913
rect 87194 252839 87250 252848
rect 87300 252777 87328 252946
rect 131354 252904 131410 252913
rect 131354 252839 131410 252848
rect 87286 252768 87342 252777
rect 87286 252703 87342 252712
rect 78914 251952 78970 251961
rect 78914 251887 78970 251896
rect 78928 251786 78956 251887
rect 131368 251854 131396 252839
rect 131356 251848 131408 251854
rect 131356 251790 131408 251796
rect 78916 251780 78968 251786
rect 78916 251722 78968 251728
rect 87196 251644 87248 251650
rect 87196 251586 87248 251592
rect 87208 251553 87236 251586
rect 87194 251544 87250 251553
rect 87194 251479 87250 251488
rect 79742 250592 79798 250601
rect 79742 250527 79798 250536
rect 79756 250358 79784 250527
rect 79744 250352 79796 250358
rect 87196 250352 87248 250358
rect 79744 250294 79796 250300
rect 87194 250320 87196 250329
rect 87248 250320 87250 250329
rect 87194 250255 87250 250264
rect 131828 250057 131856 255718
rect 131998 255624 132054 255633
rect 131998 255559 132054 255568
rect 132012 254574 132040 255559
rect 132000 254568 132052 254574
rect 132000 254510 132052 254516
rect 131998 250320 132054 250329
rect 131998 250255 132054 250264
rect 131814 250048 131870 250057
rect 131814 249983 131870 249992
rect 78916 249604 78968 249610
rect 78916 249546 78968 249552
rect 87196 249604 87248 249610
rect 87196 249546 87248 249552
rect 78928 249377 78956 249546
rect 87208 249377 87236 249546
rect 78914 249368 78970 249377
rect 78914 249303 78970 249312
rect 87194 249368 87250 249377
rect 87194 249303 87250 249312
rect 132012 248998 132040 250255
rect 132000 248992 132052 248998
rect 132104 248969 132132 261378
rect 132460 260076 132512 260082
rect 132460 260018 132512 260024
rect 132184 258648 132236 258654
rect 132184 258590 132236 258596
rect 132196 252346 132224 258590
rect 132276 257356 132328 257362
rect 132276 257298 132328 257304
rect 132288 252466 132316 257298
rect 132366 256440 132422 256449
rect 132366 256375 132422 256384
rect 132380 255934 132408 256375
rect 132368 255928 132420 255934
rect 132368 255870 132420 255876
rect 132276 252460 132328 252466
rect 132276 252402 132328 252408
rect 132196 252318 132408 252346
rect 132276 252256 132328 252262
rect 132276 252198 132328 252204
rect 132182 251136 132238 251145
rect 132182 251071 132238 251080
rect 132000 248934 132052 248940
rect 132090 248960 132146 248969
rect 132090 248895 132146 248904
rect 87194 248416 87250 248425
rect 87194 248351 87250 248360
rect 87208 248250 87236 248351
rect 78916 248244 78968 248250
rect 78916 248186 78968 248192
rect 87196 248244 87248 248250
rect 87196 248186 87248 248192
rect 78928 248017 78956 248186
rect 78914 248008 78970 248017
rect 78914 247943 78970 247952
rect 88482 247600 88538 247609
rect 78916 247564 78968 247570
rect 88482 247535 88484 247544
rect 78916 247506 78968 247512
rect 88536 247535 88538 247544
rect 88484 247506 88536 247512
rect 78928 246929 78956 247506
rect 78914 246920 78970 246929
rect 78914 246855 78970 246864
rect 87194 246648 87250 246657
rect 87194 246583 87250 246592
rect 87208 246210 87236 246583
rect 78916 246204 78968 246210
rect 78916 246146 78968 246152
rect 87196 246204 87248 246210
rect 87196 246146 87248 246152
rect 131356 246204 131408 246210
rect 131356 246146 131408 246152
rect 78928 245569 78956 246146
rect 87194 245832 87250 245841
rect 87194 245767 87250 245776
rect 78914 245560 78970 245569
rect 78914 245495 78970 245504
rect 87102 244880 87158 244889
rect 87102 244815 87158 244824
rect 78916 244776 78968 244782
rect 78916 244718 78968 244724
rect 78928 244209 78956 244718
rect 78914 244200 78970 244209
rect 78914 244135 78970 244144
rect 87010 244064 87066 244073
rect 87010 243999 87066 244008
rect 78916 243076 78968 243082
rect 78916 243018 78968 243024
rect 78928 242577 78956 243018
rect 78914 242568 78970 242577
rect 78914 242503 78970 242512
rect 79100 242192 79152 242198
rect 79100 242134 79152 242140
rect 79008 242124 79060 242130
rect 79008 242066 79060 242072
rect 78914 240664 78970 240673
rect 78914 240599 78970 240608
rect 78928 239682 78956 240599
rect 78916 239676 78968 239682
rect 78916 239618 78968 239624
rect 79020 239313 79048 242066
rect 79006 239304 79062 239313
rect 79006 239239 79062 239248
rect 79112 238633 79140 242134
rect 87024 239682 87052 243999
rect 87116 243082 87144 244815
rect 87208 244782 87236 245767
rect 131368 245569 131396 246146
rect 131354 245560 131410 245569
rect 131354 245495 131410 245504
rect 87196 244776 87248 244782
rect 87196 244718 87248 244724
rect 87286 243112 87342 243121
rect 87104 243076 87156 243082
rect 87286 243047 87342 243056
rect 87104 243018 87156 243024
rect 87194 242296 87250 242305
rect 87194 242231 87250 242240
rect 87208 242198 87236 242231
rect 87196 242192 87248 242198
rect 87196 242134 87248 242140
rect 87300 242130 87328 243047
rect 87288 242124 87340 242130
rect 87288 242066 87340 242072
rect 91670 241602 91698 241860
rect 95258 241738 95286 241860
rect 98938 241761 98966 241860
rect 95212 241710 95286 241738
rect 98924 241752 98980 241761
rect 91670 241574 91744 241602
rect 87012 239676 87064 239682
rect 87012 239618 87064 239624
rect 91716 239449 91744 241574
rect 95212 239721 95240 241710
rect 102526 241738 102554 241860
rect 106206 241738 106234 241860
rect 98924 241687 98980 241696
rect 102480 241710 102554 241738
rect 106160 241710 106234 241738
rect 95198 239712 95254 239721
rect 95198 239647 95254 239656
rect 91702 239440 91758 239449
rect 91702 239375 91758 239384
rect 79098 238624 79154 238633
rect 79098 238559 79154 238568
rect 102480 237953 102508 241710
rect 102466 237944 102522 237953
rect 102466 237879 102522 237888
rect 78916 236616 78968 236622
rect 78914 236584 78916 236593
rect 78968 236584 78970 236593
rect 78914 236519 78970 236528
rect 106160 235777 106188 241710
rect 109794 241602 109822 241860
rect 113474 241738 113502 241860
rect 117062 241738 117090 241860
rect 113474 241710 113548 241738
rect 117062 241710 117136 241738
rect 109288 241574 109822 241602
rect 106146 235768 106202 235777
rect 106146 235703 106202 235712
rect 109288 232814 109316 241574
rect 113520 235126 113548 241710
rect 117108 235913 117136 241710
rect 120742 241602 120770 241860
rect 124330 241654 124358 241860
rect 120328 241574 120770 241602
rect 123076 241648 123128 241654
rect 123076 241590 123128 241596
rect 124318 241648 124370 241654
rect 128010 241602 128038 241860
rect 124318 241590 124370 241596
rect 117094 235904 117150 235913
rect 117094 235839 117150 235848
rect 113508 235120 113560 235126
rect 113508 235062 113560 235068
rect 113876 235120 113928 235126
rect 113876 235062 113928 235068
rect 113888 234446 113916 235062
rect 113876 234440 113928 234446
rect 113876 234382 113928 234388
rect 109276 232808 109328 232814
rect 109276 232750 109328 232756
rect 76800 230904 76852 230910
rect 76800 230846 76852 230852
rect 115992 230428 116044 230434
rect 115992 230370 116044 230376
rect 103480 230360 103532 230366
rect 103480 230302 103532 230308
rect 91060 230292 91112 230298
rect 91060 230234 91112 230240
rect 91072 227716 91100 230234
rect 103492 227716 103520 230302
rect 116004 227716 116032 230370
rect 120328 230298 120356 241574
rect 123088 230366 123116 241590
rect 127228 241574 128038 241602
rect 127228 230434 127256 241574
rect 132196 239274 132224 251071
rect 132288 246113 132316 252198
rect 132380 247065 132408 252318
rect 132472 248289 132500 260018
rect 132552 254500 132604 254506
rect 132552 254442 132604 254448
rect 132458 248280 132514 248289
rect 132458 248215 132514 248224
rect 132366 247056 132422 247065
rect 132366 246991 132422 247000
rect 132274 246104 132330 246113
rect 132274 246039 132330 246048
rect 132564 244753 132592 254442
rect 133378 252088 133434 252097
rect 133378 252023 133434 252032
rect 132644 251780 132696 251786
rect 132644 251722 132696 251728
rect 132550 244744 132606 244753
rect 132550 244679 132606 244688
rect 132552 243212 132604 243218
rect 132552 243154 132604 243160
rect 132564 243121 132592 243154
rect 132550 243112 132606 243121
rect 132550 243047 132606 243056
rect 132656 242849 132684 251722
rect 132642 242840 132698 242849
rect 132642 242775 132698 242784
rect 133392 240634 133420 252023
rect 133380 240628 133432 240634
rect 133380 240570 133432 240576
rect 132184 239268 132236 239274
rect 132184 239210 132236 239216
rect 128136 237228 128188 237234
rect 128136 237170 128188 237176
rect 128148 236622 128176 237170
rect 128136 236616 128188 236622
rect 128136 236558 128188 236564
rect 127216 230428 127268 230434
rect 127216 230370 127268 230376
rect 123076 230360 123128 230366
rect 123076 230302 123128 230308
rect 120316 230292 120368 230298
rect 120316 230234 120368 230240
rect 128148 227730 128176 236558
rect 134772 230842 134800 371742
rect 184084 367658 184112 370924
rect 186280 368672 186332 368678
rect 186280 368614 186332 368620
rect 184072 367652 184124 367658
rect 184072 367594 184124 367600
rect 185176 367652 185228 367658
rect 185176 367594 185228 367600
rect 185268 367652 185320 367658
rect 185268 367594 185320 367600
rect 185188 358682 185216 367594
rect 185176 358676 185228 358682
rect 185176 358618 185228 358624
rect 139636 357928 139688 357934
rect 139636 357870 139688 357876
rect 174044 357928 174096 357934
rect 174044 357870 174096 357876
rect 139648 357769 139676 357870
rect 139634 357760 139690 357769
rect 139634 357695 139690 357704
rect 174056 357225 174084 357870
rect 174042 357216 174098 357225
rect 174042 357151 174098 357160
rect 139636 356568 139688 356574
rect 139634 356536 139636 356545
rect 173492 356568 173544 356574
rect 139688 356536 139690 356545
rect 173492 356510 173544 356516
rect 139634 356471 139690 356480
rect 173504 356137 173532 356510
rect 173490 356128 173546 356137
rect 173490 356063 173546 356072
rect 139636 355208 139688 355214
rect 139634 355176 139636 355185
rect 174044 355208 174096 355214
rect 139688 355176 139690 355185
rect 174042 355176 174044 355185
rect 174096 355176 174098 355185
rect 139634 355111 139690 355120
rect 139728 355140 139780 355146
rect 139728 355082 139780 355088
rect 173768 355140 173820 355146
rect 174042 355111 174098 355120
rect 173768 355082 173820 355088
rect 139740 354641 139768 355082
rect 139726 354632 139782 354641
rect 139726 354567 139782 354576
rect 173780 354097 173808 355082
rect 173766 354088 173822 354097
rect 173766 354023 173822 354032
rect 139636 353848 139688 353854
rect 139636 353790 139688 353796
rect 174044 353848 174096 353854
rect 174044 353790 174096 353796
rect 139648 353553 139676 353790
rect 139634 353544 139690 353553
rect 139634 353479 139690 353488
rect 174056 353009 174084 353790
rect 174042 353000 174098 353009
rect 174042 352935 174098 352944
rect 139636 352420 139688 352426
rect 139636 352362 139688 352368
rect 174044 352420 174096 352426
rect 174044 352362 174096 352368
rect 139648 352329 139676 352362
rect 139634 352320 139690 352329
rect 139634 352255 139690 352264
rect 174056 352057 174084 352362
rect 174042 352048 174098 352057
rect 174042 351983 174098 351992
rect 180850 351640 180906 351649
rect 180850 351575 180906 351584
rect 137428 351128 137480 351134
rect 137428 351070 137480 351076
rect 137440 349706 137468 351070
rect 139636 351060 139688 351066
rect 139636 351002 139688 351008
rect 173768 351060 173820 351066
rect 173768 351002 173820 351008
rect 139648 350561 139676 351002
rect 139726 350960 139782 350969
rect 139726 350895 139782 350904
rect 139634 350552 139690 350561
rect 139634 350487 139690 350496
rect 139740 350386 139768 350895
rect 139728 350380 139780 350386
rect 139728 350322 139780 350328
rect 173780 349881 173808 351002
rect 174044 350992 174096 350998
rect 174042 350960 174044 350969
rect 174096 350960 174098 350969
rect 174042 350895 174098 350904
rect 173766 349872 173822 349881
rect 173766 349807 173822 349816
rect 137520 349768 137572 349774
rect 137520 349710 137572 349716
rect 137428 349700 137480 349706
rect 137428 349642 137480 349648
rect 137428 348408 137480 348414
rect 137428 348350 137480 348356
rect 137440 346918 137468 348350
rect 137532 348278 137560 349710
rect 139636 349700 139688 349706
rect 139636 349642 139688 349648
rect 139648 349609 139676 349642
rect 139634 349600 139690 349609
rect 139634 349535 139690 349544
rect 180864 349094 180892 351575
rect 185280 351066 185308 367594
rect 186004 358676 186056 358682
rect 186004 358618 186056 358624
rect 186016 351762 186044 358618
rect 186292 351882 186320 368614
rect 186568 367658 186596 370924
rect 189066 370910 189264 370938
rect 186556 367652 186608 367658
rect 186556 367594 186608 367600
rect 189236 354058 189264 370910
rect 191536 368678 191564 370924
rect 194034 370910 194784 370938
rect 191524 368672 191576 368678
rect 191524 368614 191576 368620
rect 194756 355078 194784 370910
rect 196228 370910 196518 370938
rect 194744 355072 194796 355078
rect 194744 355014 194796 355020
rect 189224 354052 189276 354058
rect 189224 353994 189276 354000
rect 191340 354052 191392 354058
rect 191340 353994 191392 354000
rect 186280 351876 186332 351882
rect 186280 351818 186332 351824
rect 186016 351734 186398 351762
rect 191352 351748 191380 353994
rect 196228 352426 196256 370910
rect 199080 367658 199108 370924
rect 200368 370910 201578 370938
rect 199068 367652 199120 367658
rect 199068 367594 199120 367600
rect 200264 367652 200316 367658
rect 200264 367594 200316 367600
rect 196308 355072 196360 355078
rect 196308 355014 196360 355020
rect 196216 352420 196268 352426
rect 196216 352362 196268 352368
rect 196320 351748 196348 355014
rect 200276 354058 200304 367594
rect 200264 354052 200316 354058
rect 200264 353994 200316 354000
rect 200368 353854 200396 370910
rect 204048 367658 204076 370924
rect 205980 370910 206546 370938
rect 204036 367652 204088 367658
rect 204036 367594 204088 367600
rect 205876 367652 205928 367658
rect 205876 367594 205928 367600
rect 201368 354052 201420 354058
rect 201368 353994 201420 354000
rect 200356 353848 200408 353854
rect 200356 353790 200408 353796
rect 201380 351748 201408 353994
rect 205888 351762 205916 367594
rect 205980 355146 206008 370910
rect 209016 368610 209044 370924
rect 211408 370910 211606 370938
rect 209004 368604 209056 368610
rect 209004 368546 209056 368552
rect 210016 368604 210068 368610
rect 210016 368546 210068 368552
rect 210028 363510 210056 368546
rect 210016 363504 210068 363510
rect 210016 363446 210068 363452
rect 211028 363504 211080 363510
rect 211028 363446 211080 363452
rect 205968 355140 206020 355146
rect 205968 355082 206020 355088
rect 211040 351762 211068 363446
rect 211408 355214 211436 370910
rect 214076 367658 214104 370924
rect 215640 370910 216574 370938
rect 219058 370910 219624 370938
rect 214064 367652 214116 367658
rect 214064 367594 214116 367600
rect 215536 367652 215588 367658
rect 215536 367594 215588 367600
rect 211396 355208 211448 355214
rect 211396 355150 211448 355156
rect 215548 351898 215576 367594
rect 215640 356574 215668 370910
rect 215628 356568 215680 356574
rect 215628 356510 215680 356516
rect 219596 353922 219624 370910
rect 221068 370910 221542 370938
rect 221068 357934 221096 370910
rect 221056 357928 221108 357934
rect 221056 357870 221108 357876
rect 219584 353916 219636 353922
rect 219584 353858 219636 353864
rect 221332 353916 221384 353922
rect 221332 353858 221384 353864
rect 215548 351870 215852 351898
rect 205888 351734 206362 351762
rect 211040 351734 211330 351762
rect 215824 351626 215852 351870
rect 221344 351748 221372 353858
rect 215824 351598 216390 351626
rect 185268 351060 185320 351066
rect 185268 351002 185320 351008
rect 180942 350008 180998 350017
rect 180942 349943 180998 349952
rect 173032 349088 173084 349094
rect 173032 349030 173084 349036
rect 180852 349088 180904 349094
rect 180852 349030 180904 349036
rect 173044 348929 173072 349030
rect 173030 348920 173086 348929
rect 173030 348855 173086 348864
rect 137612 348340 137664 348346
rect 137612 348282 137664 348288
rect 137520 348272 137572 348278
rect 137520 348214 137572 348220
rect 137428 346912 137480 346918
rect 137428 346854 137480 346860
rect 137624 346850 137652 348282
rect 139636 348272 139688 348278
rect 139634 348240 139636 348249
rect 139688 348240 139690 348249
rect 139634 348175 139690 348184
rect 180956 348006 180984 349943
rect 182322 349600 182378 349609
rect 182322 349535 182378 349544
rect 182138 348648 182194 348657
rect 182138 348583 182194 348592
rect 172940 348000 172992 348006
rect 172940 347942 172992 347948
rect 180944 348000 180996 348006
rect 180944 347942 180996 347948
rect 172952 347841 172980 347942
rect 172938 347832 172994 347841
rect 172938 347767 172994 347776
rect 180942 347288 180998 347297
rect 180942 347223 180998 347232
rect 139820 346980 139872 346986
rect 139820 346922 139872 346928
rect 139636 346912 139688 346918
rect 139634 346880 139636 346889
rect 139688 346880 139690 346889
rect 137612 346844 137664 346850
rect 139634 346815 139690 346824
rect 139728 346844 139780 346850
rect 137612 346786 137664 346792
rect 139728 346786 139780 346792
rect 139740 346345 139768 346786
rect 139726 346336 139782 346345
rect 139726 346271 139782 346280
rect 139636 345620 139688 345626
rect 139636 345562 139688 345568
rect 139648 344169 139676 345562
rect 139832 345393 139860 346922
rect 174044 346912 174096 346918
rect 174042 346880 174044 346889
rect 174096 346880 174098 346889
rect 173768 346844 173820 346850
rect 174042 346815 174098 346824
rect 173768 346786 173820 346792
rect 173780 345801 173808 346786
rect 173766 345792 173822 345801
rect 173766 345727 173822 345736
rect 172848 345688 172900 345694
rect 172848 345630 172900 345636
rect 139818 345384 139874 345393
rect 139818 345319 139874 345328
rect 172756 344804 172808 344810
rect 172756 344746 172808 344752
rect 172768 344713 172796 344746
rect 172754 344704 172810 344713
rect 172754 344639 172810 344648
rect 139820 344260 139872 344266
rect 139820 344202 139872 344208
rect 139728 344192 139780 344198
rect 139634 344160 139690 344169
rect 139728 344134 139780 344140
rect 139634 344095 139690 344104
rect 137520 342832 137572 342838
rect 137520 342774 137572 342780
rect 135404 341540 135456 341546
rect 135404 341482 135456 341488
rect 135312 341472 135364 341478
rect 135312 341414 135364 341420
rect 135324 338554 135352 341414
rect 135416 338622 135444 341482
rect 137532 340050 137560 342774
rect 139636 342764 139688 342770
rect 139636 342706 139688 342712
rect 139648 342673 139676 342706
rect 139634 342664 139690 342673
rect 139634 342599 139690 342608
rect 139740 342265 139768 344134
rect 139726 342256 139782 342265
rect 139726 342191 139782 342200
rect 139832 341313 139860 344202
rect 172860 343761 172888 345630
rect 172940 345620 172992 345626
rect 172940 345562 172992 345568
rect 172846 343752 172902 343761
rect 172846 343687 172902 343696
rect 172756 342764 172808 342770
rect 172756 342706 172808 342712
rect 172768 341585 172796 342706
rect 172952 342673 172980 345562
rect 180956 344810 180984 347223
rect 181586 346880 181642 346889
rect 182152 346850 182180 348583
rect 182336 346918 182364 349535
rect 182324 346912 182376 346918
rect 182324 346854 182376 346860
rect 181586 346815 181642 346824
rect 182140 346844 182192 346850
rect 181600 345694 181628 346815
rect 182140 346786 182192 346792
rect 182322 346064 182378 346073
rect 182322 345999 182378 346008
rect 181588 345688 181640 345694
rect 181588 345630 181640 345636
rect 182336 345626 182364 345999
rect 182324 345620 182376 345626
rect 182324 345562 182376 345568
rect 180944 344804 180996 344810
rect 180944 344746 180996 344752
rect 180942 344704 180998 344713
rect 180942 344639 180998 344648
rect 173124 344192 173176 344198
rect 173124 344134 173176 344140
rect 172938 342664 172994 342673
rect 172938 342599 172994 342608
rect 172754 341576 172810 341585
rect 172754 341511 172810 341520
rect 139818 341304 139874 341313
rect 139818 341239 139874 341248
rect 173136 340633 173164 344134
rect 173952 342832 174004 342838
rect 173952 342774 174004 342780
rect 173768 341540 173820 341546
rect 173768 341482 173820 341488
rect 173122 340624 173178 340633
rect 173122 340559 173178 340568
rect 139544 340112 139596 340118
rect 139544 340054 139596 340060
rect 137520 340044 137572 340050
rect 137520 339986 137572 339992
rect 136140 338752 136192 338758
rect 136140 338694 136192 338700
rect 135404 338616 135456 338622
rect 135404 338558 135456 338564
rect 135312 338548 135364 338554
rect 135312 338490 135364 338496
rect 136152 334474 136180 338694
rect 136232 337324 136284 337330
rect 136232 337266 136284 337272
rect 136140 334468 136192 334474
rect 136140 334410 136192 334416
rect 136244 334270 136272 337266
rect 139556 336825 139584 340054
rect 139636 340044 139688 340050
rect 139636 339986 139688 339992
rect 139648 339953 139676 339986
rect 139634 339944 139690 339953
rect 139634 339879 139690 339888
rect 139636 338684 139688 338690
rect 139636 338626 139688 338632
rect 173492 338684 173544 338690
rect 173492 338626 173544 338632
rect 139542 336816 139598 336825
rect 139542 336751 139598 336760
rect 137612 336032 137664 336038
rect 137612 335974 137664 335980
rect 136232 334264 136284 334270
rect 136232 334206 136284 334212
rect 136876 334196 136928 334202
rect 136876 334138 136928 334144
rect 134852 333788 134904 333794
rect 134852 333730 134904 333736
rect 134864 232406 134892 333730
rect 136888 332201 136916 334138
rect 137060 334128 137112 334134
rect 137060 334070 137112 334076
rect 136874 332192 136930 332201
rect 136874 332127 136930 332136
rect 136888 307857 136916 332127
rect 137072 331521 137100 334070
rect 137336 334060 137388 334066
rect 137336 334002 137388 334008
rect 137058 331512 137114 331521
rect 137058 331447 137114 331456
rect 136968 326920 137020 326926
rect 136968 326862 137020 326868
rect 136980 326518 137008 326862
rect 136968 326512 137020 326518
rect 136968 326454 137020 326460
rect 136874 307848 136930 307857
rect 136874 307783 136930 307792
rect 136980 304185 137008 326454
rect 137072 314113 137100 331447
rect 137348 327606 137376 334002
rect 137520 333992 137572 333998
rect 137520 333934 137572 333940
rect 137532 328778 137560 333934
rect 137624 333114 137652 335974
rect 139648 335873 139676 338626
rect 139728 338616 139780 338622
rect 139726 338584 139728 338593
rect 139780 338584 139782 338593
rect 139726 338519 139782 338528
rect 139820 338548 139872 338554
rect 139820 338490 139872 338496
rect 139832 338049 139860 338490
rect 139818 338040 139874 338049
rect 139818 337975 139874 337984
rect 172848 336032 172900 336038
rect 172848 335974 172900 335980
rect 139820 335964 139872 335970
rect 139820 335906 139872 335912
rect 139634 335864 139690 335873
rect 139634 335799 139690 335808
rect 139636 334468 139688 334474
rect 139636 334410 139688 334416
rect 139648 334377 139676 334410
rect 139634 334368 139690 334377
rect 139634 334303 139690 334312
rect 139636 334264 139688 334270
rect 139636 334206 139688 334212
rect 139648 333969 139676 334206
rect 139634 333960 139690 333969
rect 137704 333924 137756 333930
rect 139634 333895 139690 333904
rect 137704 333866 137756 333872
rect 137612 333108 137664 333114
rect 137612 333050 137664 333056
rect 137716 329034 137744 333866
rect 137796 333856 137848 333862
rect 137796 333798 137848 333804
rect 137704 329028 137756 329034
rect 137704 328970 137756 328976
rect 137532 328750 137744 328778
rect 137716 327606 137744 328750
rect 137336 327600 137388 327606
rect 137336 327542 137388 327548
rect 137520 327600 137572 327606
rect 137520 327542 137572 327548
rect 137704 327600 137756 327606
rect 137704 327542 137756 327548
rect 137058 314104 137114 314113
rect 137058 314039 137114 314048
rect 137532 310985 137560 327542
rect 137612 326988 137664 326994
rect 137612 326930 137664 326936
rect 137518 310976 137574 310985
rect 137518 310911 137574 310920
rect 136966 304176 137022 304185
rect 136966 304111 137022 304120
rect 137518 304176 137574 304185
rect 137518 304111 137574 304120
rect 136874 301592 136930 301601
rect 136874 301527 136930 301536
rect 136888 284873 136916 301527
rect 136874 284864 136930 284873
rect 136874 284799 136930 284808
rect 136888 279433 136916 284799
rect 136874 279424 136930 279433
rect 136874 279359 136930 279368
rect 137532 275178 137560 304111
rect 137624 298609 137652 326930
rect 137716 317241 137744 327542
rect 137808 327470 137836 333798
rect 139636 333108 139688 333114
rect 139636 333050 139688 333056
rect 139648 333017 139676 333050
rect 139634 333008 139690 333017
rect 139634 332943 139690 332952
rect 139832 331657 139860 335906
rect 172860 332337 172888 335974
rect 172940 335964 172992 335970
rect 172940 335906 172992 335912
rect 172846 332328 172902 332337
rect 172846 332263 172902 332272
rect 139818 331648 139874 331657
rect 139818 331583 139874 331592
rect 172952 331249 172980 335906
rect 173504 335465 173532 338626
rect 173780 337505 173808 341482
rect 173860 340112 173912 340118
rect 173860 340054 173912 340060
rect 173766 337496 173822 337505
rect 173766 337431 173822 337440
rect 173676 337324 173728 337330
rect 173676 337266 173728 337272
rect 173490 335456 173546 335465
rect 173490 335391 173546 335400
rect 173688 333289 173716 337266
rect 173872 336417 173900 340054
rect 173964 339545 173992 342774
rect 180956 342770 180984 344639
rect 182322 344296 182378 344305
rect 182322 344231 182378 344240
rect 182336 344198 182364 344231
rect 182324 344192 182376 344198
rect 182324 344134 182376 344140
rect 181402 343344 181458 343353
rect 181402 343279 181458 343288
rect 181416 342838 181444 343279
rect 181404 342832 181456 342838
rect 181404 342774 181456 342780
rect 180944 342764 180996 342770
rect 180944 342706 180996 342712
rect 181402 342392 181458 342401
rect 181402 342327 181458 342336
rect 181416 341478 181444 342327
rect 182322 341576 182378 341585
rect 182322 341511 182324 341520
rect 182376 341511 182378 341520
rect 182324 341482 182376 341488
rect 174044 341472 174096 341478
rect 174044 341414 174096 341420
rect 181404 341472 181456 341478
rect 181404 341414 181456 341420
rect 173950 339536 174006 339545
rect 173950 339471 174006 339480
rect 174056 338593 174084 341414
rect 181402 340624 181458 340633
rect 181402 340559 181458 340568
rect 181416 340118 181444 340559
rect 181404 340112 181456 340118
rect 181404 340054 181456 340060
rect 181586 339808 181642 339817
rect 181586 339743 181642 339752
rect 180298 339400 180354 339409
rect 180298 339335 180354 339344
rect 174042 338584 174098 338593
rect 174042 338519 174098 338528
rect 173858 336408 173914 336417
rect 173858 336343 173914 336352
rect 180312 334406 180340 339335
rect 181600 338690 181628 339743
rect 181588 338684 181640 338690
rect 181588 338626 181640 338632
rect 181770 338040 181826 338049
rect 181770 337975 181826 337984
rect 181784 337330 181812 337975
rect 181772 337324 181824 337330
rect 181772 337266 181824 337272
rect 181586 337088 181642 337097
rect 181586 337023 181642 337032
rect 181600 336038 181628 337023
rect 181770 336272 181826 336281
rect 181770 336207 181826 336216
rect 181588 336032 181640 336038
rect 181588 335974 181640 335980
rect 181784 335970 181812 336207
rect 181772 335964 181824 335970
rect 181772 335906 181824 335912
rect 187948 335958 188882 335986
rect 192088 335958 192194 335986
rect 194848 335958 195506 335986
rect 198804 335958 198910 335986
rect 218584 335958 218874 335986
rect 221896 335958 222186 335986
rect 185570 335822 185952 335850
rect 174044 334400 174096 334406
rect 174042 334368 174044 334377
rect 180300 334400 180352 334406
rect 174096 334368 174098 334377
rect 180300 334342 180352 334348
rect 174042 334303 174098 334312
rect 185084 333856 185136 333862
rect 185084 333798 185136 333804
rect 173674 333280 173730 333289
rect 173674 333215 173730 333224
rect 172938 331240 172994 331249
rect 172938 331175 172994 331184
rect 140554 330288 140610 330297
rect 140554 330223 140610 330232
rect 173398 330288 173454 330297
rect 173398 330223 173454 330232
rect 140568 329238 140596 330223
rect 159598 330152 159654 330161
rect 159654 330110 159764 330138
rect 159598 330087 159654 330096
rect 155900 329974 155960 330002
rect 156820 329974 156880 330002
rect 142408 329838 143388 329866
rect 144308 329838 144644 329866
rect 145228 329838 145564 329866
rect 140556 329232 140608 329238
rect 140556 329174 140608 329180
rect 137888 329028 137940 329034
rect 137888 328970 137940 328976
rect 137796 327464 137848 327470
rect 137796 327406 137848 327412
rect 137702 317232 137758 317241
rect 137702 317167 137758 317176
rect 137704 309716 137756 309722
rect 137704 309658 137756 309664
rect 137610 298600 137666 298609
rect 137610 298535 137666 298544
rect 137610 285272 137666 285281
rect 137610 285207 137666 285216
rect 137520 275172 137572 275178
rect 137520 275114 137572 275120
rect 137532 273857 137560 275114
rect 137518 273848 137574 273857
rect 137518 273783 137574 273792
rect 136140 254636 136192 254642
rect 136140 254578 136192 254584
rect 136152 246210 136180 254578
rect 136232 254568 136284 254574
rect 136232 254510 136284 254516
rect 136244 247298 136272 254510
rect 137520 253140 137572 253146
rect 137520 253082 137572 253088
rect 136232 247292 136284 247298
rect 136232 247234 136284 247240
rect 136140 246204 136192 246210
rect 136140 246146 136192 246152
rect 137532 243218 137560 253082
rect 137520 243212 137572 243218
rect 137520 243154 137572 243160
rect 136874 235904 136930 235913
rect 136874 235839 136930 235848
rect 136888 235330 136916 235839
rect 137058 235768 137114 235777
rect 137058 235703 137114 235712
rect 136876 235324 136928 235330
rect 136876 235266 136928 235272
rect 137072 235262 137100 235703
rect 137244 235324 137296 235330
rect 137244 235266 137296 235272
rect 137060 235256 137112 235262
rect 137060 235198 137112 235204
rect 136874 235088 136930 235097
rect 136874 235023 136930 235032
rect 134852 232400 134904 232406
rect 134852 232342 134904 232348
rect 134760 230836 134812 230842
rect 134760 230778 134812 230784
rect 128148 227702 128530 227730
rect 76800 226960 76852 226966
rect 76800 226902 76852 226908
rect 76156 219548 76208 219554
rect 76156 219490 76208 219496
rect 75418 217408 75474 217417
rect 75418 217343 75474 217352
rect 74682 210200 74738 210209
rect 74682 210135 74738 210144
rect 74406 204896 74462 204905
rect 74406 204831 74462 204840
rect 74420 204769 74448 204831
rect 74406 204760 74462 204769
rect 74406 204695 74462 204704
rect 74224 203364 74276 203370
rect 74224 203306 74276 203312
rect 74222 195240 74278 195249
rect 74222 195175 74278 195184
rect 74498 195240 74554 195249
rect 74498 195175 74554 195184
rect 74236 195113 74264 195175
rect 74512 195113 74540 195175
rect 74222 195104 74278 195113
rect 74222 195039 74278 195048
rect 74498 195104 74554 195113
rect 74498 195039 74554 195048
rect 74130 188032 74186 188041
rect 74186 187990 74264 188018
rect 74130 187967 74186 187976
rect 74236 185593 74264 187990
rect 75432 186846 75460 217343
rect 75420 186840 75472 186846
rect 75420 186782 75472 186788
rect 74314 185720 74370 185729
rect 74314 185655 74370 185664
rect 74222 185584 74278 185593
rect 74222 185519 74278 185528
rect 74038 185040 74094 185049
rect 74038 184975 74094 184984
rect 55298 182822 55404 182850
rect 56126 182822 56784 182850
rect 51512 179830 51632 179858
rect 51604 170338 51632 179830
rect 53522 172936 53578 172945
rect 53522 172871 53578 172880
rect 54534 172936 54590 172945
rect 54534 172871 54590 172880
rect 51604 170310 52000 170338
rect 51972 169794 52000 170310
rect 49948 169766 50422 169794
rect 51328 169766 51434 169794
rect 51972 169766 52446 169794
rect 53536 169780 53564 172871
rect 54548 169780 54576 172871
rect 55376 172498 55404 182822
rect 55546 172936 55602 172945
rect 55546 172871 55602 172880
rect 55364 172492 55416 172498
rect 55364 172434 55416 172440
rect 55560 169780 55588 172871
rect 56558 172800 56614 172809
rect 56558 172735 56614 172744
rect 56572 169780 56600 172735
rect 56756 172430 56784 182822
rect 57032 180658 57060 182836
rect 57966 182822 58072 182850
rect 58794 182822 59544 182850
rect 57020 180652 57072 180658
rect 57020 180594 57072 180600
rect 58044 172566 58072 182822
rect 59516 172634 59544 182822
rect 59700 181338 59728 182836
rect 59688 181332 59740 181338
rect 59688 181274 59740 181280
rect 59688 172900 59740 172906
rect 59688 172842 59740 172848
rect 59504 172628 59556 172634
rect 59504 172570 59556 172576
rect 58032 172560 58084 172566
rect 58032 172502 58084 172508
rect 56744 172424 56796 172430
rect 56744 172366 56796 172372
rect 58676 172084 58728 172090
rect 58676 172026 58728 172032
rect 57664 171948 57716 171954
rect 57664 171890 57716 171896
rect 57676 169780 57704 171890
rect 58688 169780 58716 172026
rect 59700 169780 59728 172842
rect 60620 172362 60648 182836
rect 61448 181338 61476 182836
rect 60884 181332 60936 181338
rect 60884 181274 60936 181280
rect 61436 181332 61488 181338
rect 61436 181274 61488 181280
rect 62264 181332 62316 181338
rect 62264 181274 62316 181280
rect 60700 173036 60752 173042
rect 60700 172978 60752 172984
rect 60608 172356 60660 172362
rect 60608 172298 60660 172304
rect 60712 169780 60740 172978
rect 60896 172770 60924 181274
rect 60884 172764 60936 172770
rect 60884 172706 60936 172712
rect 62276 172702 62304 181274
rect 62368 180522 62396 182836
rect 63000 181332 63052 181338
rect 63000 181274 63052 181280
rect 62356 180516 62408 180522
rect 62356 180458 62408 180464
rect 62264 172696 62316 172702
rect 62264 172638 62316 172644
rect 63012 172090 63040 181274
rect 63000 172084 63052 172090
rect 63000 172026 63052 172032
rect 63288 171954 63316 182836
rect 64116 181338 64144 182836
rect 64104 181332 64156 181338
rect 64104 181274 64156 181280
rect 63644 180516 63696 180522
rect 63644 180458 63696 180464
rect 63656 172838 63684 180458
rect 64840 172968 64892 172974
rect 64840 172910 64892 172916
rect 63644 172832 63696 172838
rect 63644 172774 63696 172780
rect 63828 172288 63880 172294
rect 63828 172230 63880 172236
rect 63276 171948 63328 171954
rect 63276 171890 63328 171896
rect 62816 171880 62868 171886
rect 62816 171822 62868 171828
rect 61804 171744 61856 171750
rect 61804 171686 61856 171692
rect 61816 169780 61844 171686
rect 62828 169780 62856 171822
rect 63840 169780 63868 172230
rect 64852 169780 64880 172910
rect 65036 172906 65064 182836
rect 65760 181332 65812 181338
rect 65760 181274 65812 181280
rect 65024 172900 65076 172906
rect 65024 172842 65076 172848
rect 65772 171750 65800 181274
rect 65956 173042 65984 182836
rect 66784 181338 66812 182836
rect 66772 181332 66824 181338
rect 66772 181274 66824 181280
rect 65944 173036 65996 173042
rect 65944 172978 65996 172984
rect 66956 172492 67008 172498
rect 66956 172434 67008 172440
rect 65944 172084 65996 172090
rect 65944 172026 65996 172032
rect 65760 171744 65812 171750
rect 65760 171686 65812 171692
rect 65956 169780 65984 172026
rect 66968 169780 66996 172434
rect 67704 171886 67732 182836
rect 68060 180652 68112 180658
rect 68060 180594 68112 180600
rect 67968 172424 68020 172430
rect 67968 172366 68020 172372
rect 67692 171880 67744 171886
rect 67692 171822 67744 171828
rect 67980 169780 68008 172366
rect 68072 169930 68100 180594
rect 68520 180516 68572 180522
rect 68520 180458 68572 180464
rect 68532 172974 68560 180458
rect 68520 172968 68572 172974
rect 68520 172910 68572 172916
rect 68624 172294 68652 182836
rect 69452 180522 69480 182836
rect 70386 182822 70492 182850
rect 69440 180516 69492 180522
rect 69440 180458 69492 180464
rect 70084 172560 70136 172566
rect 70084 172502 70136 172508
rect 68612 172288 68664 172294
rect 68612 172230 68664 172236
rect 68072 169902 68652 169930
rect 68624 169794 68652 169902
rect 68624 169766 69006 169794
rect 70096 169780 70124 172502
rect 70464 172090 70492 182822
rect 74328 173761 74356 185655
rect 74314 173752 74370 173761
rect 74314 173687 74370 173696
rect 75236 172832 75288 172838
rect 75236 172774 75288 172780
rect 72108 172764 72160 172770
rect 72108 172706 72160 172712
rect 71096 172628 71148 172634
rect 71096 172570 71148 172576
rect 70452 172084 70504 172090
rect 70452 172026 70504 172032
rect 71108 169780 71136 172570
rect 72120 169780 72148 172706
rect 74224 172696 74276 172702
rect 74224 172638 74276 172644
rect 73120 172356 73172 172362
rect 73120 172298 73172 172304
rect 73132 169780 73160 172298
rect 74236 169780 74264 172638
rect 75248 169780 75276 172774
rect 76168 169794 76196 219490
rect 76168 169766 76274 169794
rect 48936 169630 49410 169658
rect 71646 169536 71702 169545
rect 71646 169471 71702 169480
rect 71660 169438 71688 169471
rect 71648 169432 71700 169438
rect 71648 169374 71700 169380
rect 49200 168888 49252 168894
rect 49198 168856 49200 168865
rect 49252 168856 49254 168865
rect 49198 168791 49254 168800
rect 47082 143424 47138 143433
rect 47082 143359 47138 143368
rect 73946 142200 74002 142209
rect 73946 142135 74002 142144
rect 75418 142200 75474 142209
rect 75418 142135 75474 142144
rect 48568 141886 49410 141914
rect 49948 141886 50422 141914
rect 51328 141886 51434 141914
rect 51512 141886 52446 141914
rect 38802 127512 38858 127521
rect 38802 127447 38858 127456
rect 38816 126802 38844 127447
rect 48462 127240 48518 127249
rect 48462 127175 48518 127184
rect 48476 126802 48504 127175
rect 38804 126796 38856 126802
rect 38804 126738 38856 126744
rect 48464 126796 48516 126802
rect 48464 126738 48516 126744
rect 38252 126116 38304 126122
rect 38252 126058 38304 126064
rect 38264 125617 38292 126058
rect 38250 125608 38306 125617
rect 38250 125543 38306 125552
rect 38802 122752 38858 122761
rect 38802 122687 38858 122696
rect 38816 122654 38844 122687
rect 38804 122648 38856 122654
rect 38804 122590 38856 122596
rect 38804 120608 38856 120614
rect 38804 120550 38856 120556
rect 38816 120313 38844 120550
rect 38802 120304 38858 120313
rect 38802 120239 38858 120248
rect 38250 117584 38306 117593
rect 38250 117519 38306 117528
rect 38264 117146 38292 117519
rect 38252 117140 38304 117146
rect 38252 117082 38304 117088
rect 38804 115100 38856 115106
rect 38804 115042 38856 115048
rect 38816 115009 38844 115042
rect 38802 115000 38858 115009
rect 38802 114935 38858 114944
rect 38804 112992 38856 112998
rect 38804 112934 38856 112940
rect 38816 112833 38844 112934
rect 38802 112824 38858 112833
rect 38802 112759 38858 112768
rect 38252 110952 38304 110958
rect 38252 110894 38304 110900
rect 38264 110521 38292 110894
rect 38250 110512 38306 110521
rect 38250 110447 38306 110456
rect 38802 107520 38858 107529
rect 38802 107455 38804 107464
rect 38856 107455 38858 107464
rect 38804 107426 38856 107432
rect 38804 105444 38856 105450
rect 38804 105386 38856 105392
rect 38816 105353 38844 105386
rect 38802 105344 38858 105353
rect 38802 105279 38858 105288
rect 38618 102488 38674 102497
rect 38618 102423 38674 102432
rect 38632 101370 38660 102423
rect 38620 101364 38672 101370
rect 38620 101306 38672 101312
rect 38804 100616 38856 100622
rect 38804 100558 38856 100564
rect 38816 100321 38844 100558
rect 38802 100312 38858 100321
rect 38802 100247 38858 100256
rect 38802 97864 38858 97873
rect 38802 97799 38804 97808
rect 38856 97799 38858 97808
rect 38804 97770 38856 97776
rect 38068 95788 38120 95794
rect 38068 95730 38120 95736
rect 38080 95425 38108 95730
rect 38066 95416 38122 95425
rect 38066 95351 38122 95360
rect 37606 92560 37662 92569
rect 37606 92495 37662 92504
rect 37620 92326 37648 92495
rect 48568 92326 48596 141886
rect 49948 97834 49976 141886
rect 51328 101574 51356 141886
rect 51512 134418 51540 141886
rect 53536 139625 53564 141900
rect 54548 139625 54576 141900
rect 53522 139616 53578 139625
rect 53522 139551 53578 139560
rect 54534 139616 54590 139625
rect 54534 139551 54590 139560
rect 55364 139308 55416 139314
rect 55364 139250 55416 139256
rect 51500 134412 51552 134418
rect 51500 134354 51552 134360
rect 51592 134412 51644 134418
rect 51592 134354 51644 134360
rect 51604 127362 51632 134354
rect 55376 128722 55404 139250
rect 55560 134457 55588 141900
rect 56112 141886 56586 141914
rect 55546 134448 55602 134457
rect 55546 134383 55602 134392
rect 56112 132417 56140 141886
rect 56744 139444 56796 139450
rect 56744 139386 56796 139392
rect 56098 132408 56154 132417
rect 56098 132343 56154 132352
rect 56756 131630 56784 139386
rect 57676 138634 57704 141900
rect 58124 139376 58176 139382
rect 58124 139318 58176 139324
rect 57664 138628 57716 138634
rect 57664 138570 57716 138576
rect 56100 131624 56152 131630
rect 56100 131566 56152 131572
rect 56744 131624 56796 131630
rect 56744 131566 56796 131572
rect 55298 128694 55404 128722
rect 56112 128708 56140 131566
rect 57020 130604 57072 130610
rect 57020 130546 57072 130552
rect 57032 128708 57060 130546
rect 58136 128722 58164 139318
rect 58688 138974 58716 141900
rect 59504 139512 59556 139518
rect 59504 139454 59556 139460
rect 58676 138968 58728 138974
rect 58676 138910 58728 138916
rect 59516 128858 59544 139454
rect 59700 138838 59728 141900
rect 59688 138832 59740 138838
rect 59688 138774 59740 138780
rect 60712 138702 60740 141900
rect 60884 139580 60936 139586
rect 60884 139522 60936 139528
rect 60792 139240 60844 139246
rect 60792 139182 60844 139188
rect 60700 138696 60752 138702
rect 60700 138638 60752 138644
rect 60804 131630 60832 139182
rect 59688 131624 59740 131630
rect 59688 131566 59740 131572
rect 60792 131624 60844 131630
rect 60792 131566 60844 131572
rect 59148 128830 59544 128858
rect 59148 128722 59176 128830
rect 57966 128694 58164 128722
rect 58794 128694 59176 128722
rect 59700 128708 59728 131566
rect 60896 128722 60924 139522
rect 61816 138770 61844 141900
rect 62264 139648 62316 139654
rect 62264 139590 62316 139596
rect 61804 138764 61856 138770
rect 61804 138706 61856 138712
rect 61620 138628 61672 138634
rect 61620 138570 61672 138576
rect 61632 130474 61660 138570
rect 61620 130468 61672 130474
rect 61620 130410 61672 130416
rect 62276 130338 62304 139590
rect 62828 138906 62856 141900
rect 63644 139716 63696 139722
rect 63644 139658 63696 139664
rect 63000 138968 63052 138974
rect 63000 138910 63052 138916
rect 62816 138900 62868 138906
rect 62816 138842 62868 138848
rect 62356 130400 62408 130406
rect 62356 130342 62408 130348
rect 61436 130332 61488 130338
rect 61436 130274 61488 130280
rect 62264 130332 62316 130338
rect 62264 130274 62316 130280
rect 60634 128694 60924 128722
rect 61448 128708 61476 130274
rect 62368 128708 62396 130342
rect 63012 130338 63040 138910
rect 63092 138832 63144 138838
rect 63092 138774 63144 138780
rect 63104 130542 63132 138774
rect 63184 138696 63236 138702
rect 63184 138638 63236 138644
rect 63196 130746 63224 138638
rect 63184 130740 63236 130746
rect 63184 130682 63236 130688
rect 63092 130536 63144 130542
rect 63092 130478 63144 130484
rect 63276 130468 63328 130474
rect 63276 130410 63328 130416
rect 63000 130332 63052 130338
rect 63000 130274 63052 130280
rect 63288 128708 63316 130410
rect 63656 130406 63684 139658
rect 63840 139110 63868 141900
rect 64852 139790 64880 141900
rect 64840 139784 64892 139790
rect 64840 139726 64892 139732
rect 63828 139104 63880 139110
rect 63828 139046 63880 139052
rect 64380 138968 64432 138974
rect 64380 138910 64432 138916
rect 64392 130610 64420 138910
rect 65760 138764 65812 138770
rect 65760 138706 65812 138712
rect 64380 130604 64432 130610
rect 64380 130546 64432 130552
rect 65024 130536 65076 130542
rect 65024 130478 65076 130484
rect 63644 130400 63696 130406
rect 63644 130342 63696 130348
rect 64104 130332 64156 130338
rect 64104 130274 64156 130280
rect 64116 128708 64144 130274
rect 65036 128708 65064 130478
rect 65772 130338 65800 138706
rect 65956 138634 65984 141900
rect 66968 139314 66996 141900
rect 67980 139450 68008 141900
rect 67968 139444 68020 139450
rect 67968 139386 68020 139392
rect 66956 139308 67008 139314
rect 66956 139250 67008 139256
rect 68612 139104 68664 139110
rect 68612 139046 68664 139052
rect 67692 138900 67744 138906
rect 67692 138842 67744 138848
rect 65944 138628 65996 138634
rect 65944 138570 65996 138576
rect 65944 130740 65996 130746
rect 65944 130682 65996 130688
rect 65760 130332 65812 130338
rect 65760 130274 65812 130280
rect 65956 128708 65984 130682
rect 66772 130332 66824 130338
rect 66772 130274 66824 130280
rect 66784 128708 66812 130274
rect 67704 128708 67732 138842
rect 68624 128708 68652 139046
rect 68992 138974 69020 141900
rect 70096 139382 70124 141900
rect 70452 139784 70504 139790
rect 70452 139726 70504 139732
rect 70084 139376 70136 139382
rect 70084 139318 70136 139324
rect 68980 138968 69032 138974
rect 68980 138910 69032 138916
rect 70464 129674 70492 139726
rect 71108 139518 71136 141900
rect 71096 139512 71148 139518
rect 71096 139454 71148 139460
rect 72120 139246 72148 141900
rect 73132 139586 73160 141900
rect 73960 140606 73988 142135
rect 74132 141280 74184 141286
rect 74132 141222 74184 141228
rect 73948 140600 74000 140606
rect 73948 140542 74000 140548
rect 73120 139580 73172 139586
rect 73120 139522 73172 139528
rect 72108 139240 72160 139246
rect 72108 139182 72160 139188
rect 70544 138628 70596 138634
rect 70544 138570 70596 138576
rect 69820 129646 70492 129674
rect 69820 128722 69848 129646
rect 70556 128722 70584 138570
rect 69466 128694 69848 128722
rect 70386 128694 70584 128722
rect 73960 127498 73988 140542
rect 73960 127470 74080 127498
rect 51604 127334 51724 127362
rect 51696 115174 51724 127334
rect 52602 126288 52658 126297
rect 52602 126223 52658 126232
rect 52616 126122 52644 126223
rect 52604 126116 52656 126122
rect 52604 126058 52656 126064
rect 54076 122648 54128 122654
rect 54076 122590 54128 122596
rect 54088 122081 54116 122590
rect 54074 122072 54130 122081
rect 54074 122007 54130 122016
rect 52602 121256 52658 121265
rect 52602 121191 52658 121200
rect 52616 120614 52644 121191
rect 52604 120608 52656 120614
rect 52604 120550 52656 120556
rect 73394 120576 73450 120585
rect 73394 120511 73450 120520
rect 73408 119769 73436 120511
rect 73394 119760 73450 119769
rect 73394 119695 73450 119704
rect 54074 117176 54130 117185
rect 54074 117111 54076 117120
rect 54128 117111 54130 117120
rect 54076 117082 54128 117088
rect 52142 116224 52198 116233
rect 52142 116159 52198 116168
rect 51684 115168 51736 115174
rect 51684 115110 51736 115116
rect 52156 115106 52184 116159
rect 52144 115100 52196 115106
rect 52144 115042 52196 115048
rect 51592 113740 51644 113746
rect 51592 113682 51644 113688
rect 51604 108306 51632 113682
rect 51866 113096 51922 113105
rect 51866 113031 51922 113040
rect 51880 112998 51908 113031
rect 51868 112992 51920 112998
rect 51868 112934 51920 112940
rect 52602 111328 52658 111337
rect 52602 111263 52658 111272
rect 52616 111026 52644 111263
rect 52604 111020 52656 111026
rect 52604 110962 52656 110968
rect 51592 108300 51644 108306
rect 51592 108242 51644 108248
rect 52602 106296 52658 106305
rect 52602 106231 52658 106240
rect 52616 105450 52644 106231
rect 52604 105444 52656 105450
rect 52604 105386 52656 105392
rect 51684 104084 51736 104090
rect 51684 104026 51736 104032
rect 50028 101568 50080 101574
rect 50028 101510 50080 101516
rect 51316 101568 51368 101574
rect 51316 101510 51368 101516
rect 50040 101370 50068 101510
rect 50028 101364 50080 101370
rect 50028 101306 50080 101312
rect 49936 97828 49988 97834
rect 49936 97770 49988 97776
rect 37608 92320 37660 92326
rect 37608 92262 37660 92268
rect 48556 92320 48608 92326
rect 48556 92262 48608 92268
rect 38804 90212 38856 90218
rect 38804 90154 38856 90160
rect 38816 90121 38844 90154
rect 38802 90112 38858 90121
rect 38802 90047 38858 90056
rect 36044 87424 36096 87430
rect 36044 87366 36096 87372
rect 34664 87152 34716 87158
rect 34664 87094 34716 87100
rect 36056 87090 36084 87366
rect 26568 87084 26620 87090
rect 26568 87026 26620 87032
rect 36044 87084 36096 87090
rect 36044 87026 36096 87032
rect 48568 75818 48596 92262
rect 48568 75790 48950 75818
rect 49948 75804 49976 97770
rect 50040 75682 50068 101306
rect 51696 89062 51724 104026
rect 52602 101264 52658 101273
rect 52602 101199 52658 101208
rect 52616 100622 52644 101199
rect 52604 100616 52656 100622
rect 52604 100558 52656 100564
rect 52602 96232 52658 96241
rect 52602 96167 52658 96176
rect 52616 95862 52644 96167
rect 52604 95856 52656 95862
rect 52604 95798 52656 95804
rect 73408 93754 73436 119695
rect 73486 115136 73542 115145
rect 73486 115071 73542 115080
rect 73396 93748 73448 93754
rect 73396 93690 73448 93696
rect 73396 91504 73448 91510
rect 73396 91446 73448 91452
rect 52602 91336 52658 91345
rect 52602 91271 52658 91280
rect 52616 90218 52644 91271
rect 73408 91209 73436 91446
rect 73394 91200 73450 91209
rect 73394 91135 73450 91144
rect 52604 90212 52656 90218
rect 52604 90154 52656 90160
rect 51684 89056 51736 89062
rect 51684 88998 51736 89004
rect 69544 88982 70386 89010
rect 55298 88846 55404 88874
rect 51500 86132 51552 86138
rect 51500 86074 51552 86080
rect 51512 75682 51540 86074
rect 55376 78522 55404 88846
rect 56112 86818 56140 88860
rect 57032 86886 57060 88860
rect 57966 88846 58164 88874
rect 58794 88846 59544 88874
rect 57020 86880 57072 86886
rect 57020 86822 57072 86828
rect 56100 86812 56152 86818
rect 56100 86754 56152 86760
rect 57204 79060 57256 79066
rect 57204 79002 57256 79008
rect 55364 78516 55416 78522
rect 55364 78458 55416 78464
rect 54074 78008 54130 78017
rect 54074 77943 54130 77952
rect 53062 77872 53118 77881
rect 53062 77807 53118 77816
rect 53076 75804 53104 77807
rect 54088 75804 54116 77943
rect 55086 77872 55142 77881
rect 55086 77807 55142 77816
rect 56098 77872 56154 77881
rect 56098 77807 56154 77816
rect 55100 75804 55128 77807
rect 56112 75804 56140 77807
rect 57216 75804 57244 79002
rect 58136 78930 58164 88846
rect 58124 78924 58176 78930
rect 58124 78866 58176 78872
rect 59228 78652 59280 78658
rect 59228 78594 59280 78600
rect 58216 78380 58268 78386
rect 58216 78322 58268 78328
rect 58228 75804 58256 78322
rect 59240 75804 59268 78594
rect 59516 78590 59544 88846
rect 59700 87022 59728 88860
rect 60634 88846 60924 88874
rect 59688 87016 59740 87022
rect 59688 86958 59740 86964
rect 60240 79196 60292 79202
rect 60240 79138 60292 79144
rect 59504 78584 59556 78590
rect 59504 78526 59556 78532
rect 60252 75804 60280 79138
rect 60896 78726 60924 88846
rect 61448 86138 61476 88860
rect 61620 86200 61672 86206
rect 61620 86142 61672 86148
rect 61436 86132 61488 86138
rect 61436 86074 61488 86080
rect 61632 79066 61660 86142
rect 62368 86138 62396 88860
rect 63288 86206 63316 88860
rect 63840 88846 64130 88874
rect 64760 88846 65050 88874
rect 63276 86200 63328 86206
rect 63276 86142 63328 86148
rect 62264 86132 62316 86138
rect 62264 86074 62316 86080
rect 62356 86132 62408 86138
rect 62356 86074 62408 86080
rect 63644 86132 63696 86138
rect 63644 86074 63696 86080
rect 63736 86132 63788 86138
rect 63736 86074 63788 86080
rect 61620 79060 61672 79066
rect 61620 79002 61672 79008
rect 62276 78794 62304 86074
rect 62356 78992 62408 78998
rect 62356 78934 62408 78940
rect 62264 78788 62316 78794
rect 62264 78730 62316 78736
rect 60884 78720 60936 78726
rect 60884 78662 60936 78668
rect 61344 78108 61396 78114
rect 61344 78050 61396 78056
rect 61356 75804 61384 78050
rect 62368 75804 62396 78934
rect 63656 78862 63684 86074
rect 63644 78856 63696 78862
rect 63644 78798 63696 78804
rect 63748 78658 63776 86074
rect 63736 78652 63788 78658
rect 63736 78594 63788 78600
rect 63368 78448 63420 78454
rect 63368 78390 63420 78396
rect 63380 75804 63408 78390
rect 63840 78386 63868 88846
rect 64380 87152 64432 87158
rect 64380 87094 64432 87100
rect 64392 79202 64420 87094
rect 64760 86138 64788 88846
rect 65956 87158 65984 88860
rect 65944 87152 65996 87158
rect 65944 87094 65996 87100
rect 66680 86812 66732 86818
rect 66680 86754 66732 86760
rect 64748 86132 64800 86138
rect 64748 86074 64800 86080
rect 65760 86132 65812 86138
rect 65760 86074 65812 86080
rect 64380 79196 64432 79202
rect 64380 79138 64432 79144
rect 65484 79128 65536 79134
rect 65484 79070 65536 79076
rect 64380 78924 64432 78930
rect 64380 78866 64432 78872
rect 63828 78380 63880 78386
rect 63828 78322 63880 78328
rect 64392 75804 64420 78866
rect 65496 75804 65524 79070
rect 65772 78114 65800 86074
rect 66588 86064 66640 86070
rect 66588 86006 66640 86012
rect 66600 79202 66628 86006
rect 66588 79196 66640 79202
rect 66588 79138 66640 79144
rect 66496 78516 66548 78522
rect 66496 78458 66548 78464
rect 65760 78108 65812 78114
rect 65760 78050 65812 78056
rect 66508 75804 66536 78458
rect 66692 75682 66720 86754
rect 66784 86138 66812 88860
rect 67336 88846 67718 88874
rect 67140 87016 67192 87022
rect 67140 86958 67192 86964
rect 66772 86132 66824 86138
rect 66772 86074 66824 86080
rect 67152 78794 67180 86958
rect 67232 86200 67284 86206
rect 67232 86142 67284 86148
rect 67140 78788 67192 78794
rect 67140 78730 67192 78736
rect 67244 78454 67272 86142
rect 67336 86070 67364 88846
rect 67876 86880 67928 86886
rect 67876 86822 67928 86828
rect 67324 86064 67376 86070
rect 67324 86006 67376 86012
rect 67232 78448 67284 78454
rect 67232 78390 67284 78396
rect 67888 75682 67916 86822
rect 68624 86206 68652 88860
rect 68612 86200 68664 86206
rect 68612 86142 68664 86148
rect 69452 86138 69480 88860
rect 68520 86132 68572 86138
rect 68520 86074 68572 86080
rect 69440 86132 69492 86138
rect 69440 86074 69492 86080
rect 68532 78930 68560 86074
rect 69544 86018 69572 88982
rect 72014 87528 72070 87537
rect 72014 87463 72016 87472
rect 72068 87463 72070 87472
rect 72016 87434 72068 87440
rect 73500 87294 73528 115071
rect 73578 112824 73634 112833
rect 73578 112759 73634 112768
rect 73592 87362 73620 112759
rect 73670 109560 73726 109569
rect 73670 109495 73726 109504
rect 73684 108889 73712 109495
rect 73670 108880 73726 108889
rect 73670 108815 73726 108824
rect 73684 94042 73712 108815
rect 74052 105217 74080 127470
rect 74144 116233 74172 141222
rect 74236 139654 74264 141900
rect 75248 139722 75276 141900
rect 75432 141286 75460 142135
rect 76064 142096 76116 142102
rect 76062 142064 76064 142073
rect 76116 142064 76118 142073
rect 76062 141999 76118 142008
rect 76168 141886 76274 141914
rect 75420 141280 75472 141286
rect 75420 141222 75472 141228
rect 76064 140192 76116 140198
rect 76064 140134 76116 140140
rect 75236 139716 75288 139722
rect 75236 139658 75288 139664
rect 74224 139648 74276 139654
rect 74224 139590 74276 139596
rect 74222 139480 74278 139489
rect 74222 139415 74278 139424
rect 75142 139480 75198 139489
rect 75142 139415 75198 139424
rect 74236 120585 74264 139415
rect 75156 139382 75184 139415
rect 75144 139376 75196 139382
rect 75144 139318 75196 139324
rect 76076 137177 76104 140134
rect 76062 137168 76118 137177
rect 76062 137103 76118 137112
rect 74314 126424 74370 126433
rect 74314 126359 74370 126368
rect 74222 120576 74278 120585
rect 74222 120511 74278 120520
rect 74130 116224 74186 116233
rect 74130 116159 74186 116168
rect 74144 115145 74172 116159
rect 74130 115136 74186 115145
rect 74130 115071 74186 115080
rect 74328 109530 74356 126359
rect 76168 125102 76196 141886
rect 76156 125096 76208 125102
rect 76156 125038 76208 125044
rect 75418 122752 75474 122761
rect 75418 122687 75474 122696
rect 74316 109524 74368 109530
rect 74316 109466 74368 109472
rect 74038 105208 74094 105217
rect 74038 105143 74094 105152
rect 73684 94014 73896 94042
rect 73672 93748 73724 93754
rect 73672 93690 73724 93696
rect 73580 87356 73632 87362
rect 73580 87298 73632 87304
rect 73488 87288 73540 87294
rect 73488 87230 73540 87236
rect 73500 86177 73528 87230
rect 73592 86313 73620 87298
rect 73684 87226 73712 93690
rect 73868 87430 73896 94014
rect 74052 89849 74080 105143
rect 75432 92734 75460 122687
rect 75420 92728 75472 92734
rect 75420 92670 75472 92676
rect 76812 91510 76840 226902
rect 134760 225532 134812 225538
rect 134760 225474 134812 225480
rect 81674 219584 81730 219593
rect 81674 219519 81676 219528
rect 81728 219519 81730 219528
rect 81676 219490 81728 219496
rect 81676 203364 81728 203370
rect 81676 203306 81728 203312
rect 81688 202865 81716 203306
rect 81674 202856 81730 202865
rect 81674 202791 81730 202800
rect 81676 186840 81728 186846
rect 81676 186782 81728 186788
rect 81688 186273 81716 186782
rect 81674 186264 81730 186273
rect 81674 186199 81730 186208
rect 88404 175830 88432 177940
rect 88392 175824 88444 175830
rect 88392 175766 88444 175772
rect 95488 175762 95516 177940
rect 95476 175756 95528 175762
rect 95476 175698 95528 175704
rect 96764 175212 96816 175218
rect 96764 175154 96816 175160
rect 79744 170248 79796 170254
rect 79744 170190 79796 170196
rect 79756 169137 79784 170190
rect 79742 169128 79798 169137
rect 79742 169063 79798 169072
rect 77258 167700 77314 167709
rect 77258 167635 77314 167644
rect 77272 167602 77300 167635
rect 77260 167596 77312 167602
rect 77260 167538 77312 167544
rect 87196 167596 87248 167602
rect 87196 167538 87248 167544
rect 77258 166340 77314 166349
rect 77258 166275 77314 166284
rect 77272 166242 77300 166275
rect 77260 166236 77312 166242
rect 77260 166178 77312 166184
rect 85724 166236 85776 166242
rect 85724 166178 85776 166184
rect 79742 164912 79798 164921
rect 79742 164847 79744 164856
rect 79796 164847 79798 164856
rect 85632 164876 85684 164882
rect 79744 164818 79796 164824
rect 85632 164818 85684 164824
rect 77258 163484 77314 163493
rect 77258 163419 77314 163428
rect 77166 162124 77222 162133
rect 77166 162059 77222 162068
rect 77180 160598 77208 162059
rect 77272 162026 77300 163419
rect 77260 162020 77312 162026
rect 77260 161962 77312 161968
rect 85644 161958 85672 164818
rect 85736 163386 85764 166178
rect 87208 164105 87236 167538
rect 87194 164096 87250 164105
rect 87194 164031 87250 164040
rect 96776 163810 96804 175154
rect 102664 175150 102692 177940
rect 109748 175218 109776 177940
rect 109736 175212 109788 175218
rect 109736 175154 109788 175160
rect 102652 175144 102704 175150
rect 102652 175086 102704 175092
rect 116924 166854 116952 177940
rect 124008 170254 124036 177940
rect 131184 174470 131212 177940
rect 124364 174464 124416 174470
rect 124364 174406 124416 174412
rect 131172 174464 131224 174470
rect 131172 174406 131224 174412
rect 123996 170248 124048 170254
rect 123996 170190 124048 170196
rect 124008 169574 124036 170190
rect 123996 169568 124048 169574
rect 123996 169510 124048 169516
rect 110196 166848 110248 166854
rect 110196 166790 110248 166796
rect 116912 166848 116964 166854
rect 116912 166790 116964 166796
rect 110208 163810 110236 166790
rect 124376 166378 124404 174406
rect 132184 168956 132236 168962
rect 132184 168898 132236 168904
rect 128136 168548 128188 168554
rect 128136 168490 128188 168496
rect 123536 166372 123588 166378
rect 123536 166314 123588 166320
rect 124364 166372 124416 166378
rect 124364 166314 124416 166320
rect 123548 163810 123576 166314
rect 96560 163782 96804 163810
rect 109900 163782 110236 163810
rect 123240 163782 123576 163810
rect 85724 163380 85776 163386
rect 85724 163322 85776 163328
rect 87196 163380 87248 163386
rect 87196 163322 87248 163328
rect 87208 163153 87236 163322
rect 87194 163144 87250 163153
rect 87194 163079 87250 163088
rect 87196 162020 87248 162026
rect 87196 161962 87248 161968
rect 85632 161952 85684 161958
rect 85632 161894 85684 161900
rect 87208 161385 87236 161962
rect 87288 161952 87340 161958
rect 87286 161920 87288 161929
rect 87340 161920 87342 161929
rect 87286 161855 87342 161864
rect 87194 161376 87250 161385
rect 87194 161311 87250 161320
rect 77168 160592 77220 160598
rect 77168 160534 77220 160540
rect 87196 160592 87248 160598
rect 87196 160534 87248 160540
rect 87208 160433 87236 160534
rect 87194 160424 87250 160433
rect 87194 160359 87250 160368
rect 81674 160016 81730 160025
rect 81674 159951 81730 159960
rect 79282 159336 79338 159345
rect 79282 159271 79284 159280
rect 79336 159271 79338 159280
rect 79284 159242 79336 159248
rect 81688 159102 81716 159951
rect 87288 159164 87340 159170
rect 87288 159106 87340 159112
rect 81676 159096 81728 159102
rect 81676 159038 81728 159044
rect 87196 159096 87248 159102
rect 87196 159038 87248 159044
rect 87208 158937 87236 159038
rect 87194 158928 87250 158937
rect 87194 158863 87250 158872
rect 87300 158665 87328 159106
rect 87286 158656 87342 158665
rect 87286 158591 87342 158600
rect 79742 157976 79798 157985
rect 79742 157911 79744 157920
rect 79796 157911 79798 157920
rect 87196 157940 87248 157946
rect 79744 157882 79796 157888
rect 87196 157882 87248 157888
rect 87208 157849 87236 157882
rect 87194 157840 87250 157849
rect 87194 157775 87250 157784
rect 77258 156548 77314 156557
rect 77258 156483 77260 156492
rect 77312 156483 77314 156492
rect 77260 156454 77312 156460
rect 87196 156444 87248 156450
rect 87196 156386 87248 156392
rect 87208 156353 87236 156386
rect 87194 156344 87250 156353
rect 87194 156279 87250 156288
rect 87194 155392 87250 155401
rect 87194 155327 87250 155336
rect 79742 155120 79798 155129
rect 87208 155090 87236 155327
rect 79742 155055 79744 155064
rect 79796 155055 79798 155064
rect 87196 155084 87248 155090
rect 79744 155026 79796 155032
rect 87196 155026 87248 155032
rect 87194 154440 87250 154449
rect 79744 154404 79796 154410
rect 87194 154375 87196 154384
rect 79744 154346 79796 154352
rect 87248 154375 87250 154384
rect 87196 154346 87248 154352
rect 79756 153769 79784 154346
rect 79742 153760 79798 153769
rect 79742 153695 79798 153704
rect 87194 153624 87250 153633
rect 87194 153559 87250 153568
rect 87208 153050 87236 153559
rect 79744 153044 79796 153050
rect 79744 152986 79796 152992
rect 87196 153044 87248 153050
rect 87196 152986 87248 152992
rect 79756 152409 79784 152986
rect 87194 152672 87250 152681
rect 87194 152607 87250 152616
rect 87208 152438 87236 152607
rect 85816 152432 85868 152438
rect 79742 152400 79798 152409
rect 85816 152374 85868 152380
rect 87196 152432 87248 152438
rect 87196 152374 87248 152380
rect 79742 152335 79798 152344
rect 77258 150836 77314 150845
rect 77258 150771 77314 150780
rect 77272 149854 77300 150771
rect 85828 149854 85856 152374
rect 87470 151856 87526 151865
rect 87470 151791 87526 151800
rect 87484 151418 87512 151791
rect 85908 151412 85960 151418
rect 85908 151354 85960 151360
rect 87472 151412 87524 151418
rect 87472 151354 87524 151360
rect 77260 149848 77312 149854
rect 77260 149790 77312 149796
rect 85816 149848 85868 149854
rect 85816 149790 85868 149796
rect 80112 149644 80164 149650
rect 80112 149586 80164 149592
rect 78914 149000 78970 149009
rect 78914 148935 78970 148944
rect 76982 148592 77038 148601
rect 76982 148527 77038 148536
rect 76890 145872 76946 145881
rect 76890 145807 76946 145816
rect 76904 143394 76932 145807
rect 76996 144113 77024 148527
rect 78928 148494 78956 148935
rect 78916 148488 78968 148494
rect 78916 148430 78968 148436
rect 78914 147912 78970 147921
rect 78914 147847 78970 147856
rect 78928 147746 78956 147847
rect 78916 147740 78968 147746
rect 78916 147682 78968 147688
rect 80124 146697 80152 149586
rect 85920 148494 85948 151354
rect 87010 150904 87066 150913
rect 87010 150839 87066 150848
rect 85908 148488 85960 148494
rect 85908 148430 85960 148436
rect 87024 147746 87052 150839
rect 87194 150088 87250 150097
rect 87194 150023 87250 150032
rect 87208 149650 87236 150023
rect 87196 149644 87248 149650
rect 87196 149586 87248 149592
rect 87194 149136 87250 149145
rect 87194 149071 87250 149080
rect 87102 148320 87158 148329
rect 87102 148255 87158 148264
rect 87012 147740 87064 147746
rect 87012 147682 87064 147688
rect 80110 146688 80166 146697
rect 80110 146623 80166 146632
rect 79376 145428 79428 145434
rect 79376 145370 79428 145376
rect 79388 145337 79416 145370
rect 79374 145328 79430 145337
rect 79374 145263 79430 145272
rect 76982 144104 77038 144113
rect 76982 144039 77038 144048
rect 78914 143560 78970 143569
rect 78914 143495 78970 143504
rect 76892 143388 76944 143394
rect 76892 143330 76944 143336
rect 78928 143258 78956 143495
rect 87116 143258 87144 148255
rect 87208 145434 87236 149071
rect 91670 147626 91698 147884
rect 95258 147626 95286 147884
rect 98938 147762 98966 147884
rect 98892 147734 98966 147762
rect 91670 147598 91744 147626
rect 95258 147598 95332 147626
rect 91716 145434 91744 147598
rect 87196 145428 87248 145434
rect 87196 145370 87248 145376
rect 91704 145428 91756 145434
rect 91704 145370 91756 145376
rect 91244 144748 91296 144754
rect 91244 144690 91296 144696
rect 88576 143388 88628 143394
rect 88576 143330 88628 143336
rect 78916 143252 78968 143258
rect 78916 143194 78968 143200
rect 87104 143252 87156 143258
rect 87104 143194 87156 143200
rect 88588 142889 88616 143330
rect 88574 142880 88630 142889
rect 88574 142815 88630 142824
rect 78914 141928 78970 141937
rect 78914 141863 78970 141872
rect 78928 141354 78956 141863
rect 78916 141348 78968 141354
rect 78916 141290 78968 141296
rect 91256 133754 91284 144690
rect 95304 144113 95332 147598
rect 98892 144249 98920 147734
rect 102526 147626 102554 147884
rect 106206 147762 106234 147884
rect 109794 147762 109822 147884
rect 102388 147598 102554 147626
rect 106160 147734 106234 147762
rect 109748 147734 109822 147762
rect 98878 144240 98934 144249
rect 98878 144175 98934 144184
rect 95290 144104 95346 144113
rect 95290 144039 95346 144048
rect 95304 143938 95332 144039
rect 95292 143932 95344 143938
rect 95292 143874 95344 143880
rect 102388 140606 102416 147598
rect 103664 144816 103716 144822
rect 103664 144758 103716 144764
rect 102376 140600 102428 140606
rect 102376 140542 102428 140548
rect 103676 133754 103704 144758
rect 106160 141937 106188 147734
rect 109748 143297 109776 147734
rect 113474 147626 113502 147884
rect 117062 147626 117090 147884
rect 120742 147626 120770 147884
rect 124330 147626 124358 147884
rect 128024 147870 128084 147898
rect 113428 147598 113502 147626
rect 116188 147598 117090 147626
rect 120696 147598 120770 147626
rect 124284 147598 124358 147626
rect 109734 143288 109790 143297
rect 109734 143223 109790 143232
rect 106146 141928 106202 141937
rect 106146 141863 106202 141872
rect 113428 141286 113456 147598
rect 116084 144884 116136 144890
rect 116084 144826 116136 144832
rect 113416 141280 113468 141286
rect 113416 141222 113468 141228
rect 113876 141280 113928 141286
rect 113876 141222 113928 141228
rect 113888 140674 113916 141222
rect 113876 140668 113928 140674
rect 113876 140610 113928 140616
rect 116096 133754 116124 144826
rect 116188 139518 116216 147598
rect 120696 144754 120724 147598
rect 124284 144822 124312 147598
rect 128056 144890 128084 147870
rect 128148 145434 128176 168490
rect 132092 166236 132144 166242
rect 132092 166178 132144 166184
rect 131356 163448 131408 163454
rect 131354 163416 131356 163425
rect 131408 163416 131410 163425
rect 131354 163351 131410 163360
rect 131998 162464 132054 162473
rect 131998 162399 132054 162408
rect 132012 162162 132040 162399
rect 132000 162156 132052 162162
rect 132000 162098 132052 162104
rect 131908 162088 131960 162094
rect 131908 162030 131960 162036
rect 131538 161648 131594 161657
rect 131538 161583 131594 161592
rect 131356 160728 131408 160734
rect 131354 160696 131356 160705
rect 131408 160696 131410 160705
rect 131354 160631 131410 160640
rect 131354 158928 131410 158937
rect 131354 158863 131410 158872
rect 131368 158014 131396 158863
rect 131356 158008 131408 158014
rect 131356 157950 131408 157956
rect 131552 153730 131580 161583
rect 131724 160660 131776 160666
rect 131724 160602 131776 160608
rect 131632 157940 131684 157946
rect 131632 157882 131684 157888
rect 131540 153724 131592 153730
rect 131540 153666 131592 153672
rect 131356 149508 131408 149514
rect 131356 149450 131408 149456
rect 131368 149145 131396 149450
rect 131354 149136 131410 149145
rect 131354 149071 131410 149080
rect 131644 148873 131672 157882
rect 131736 150505 131764 160602
rect 131814 159880 131870 159889
rect 131814 159815 131870 159824
rect 131722 150496 131778 150505
rect 131722 150431 131778 150440
rect 131828 149582 131856 159815
rect 131920 150913 131948 162030
rect 132000 162020 132052 162026
rect 132000 161962 132052 161968
rect 132012 155129 132040 161962
rect 131998 155120 132054 155129
rect 131998 155055 132054 155064
rect 132104 153633 132132 166178
rect 132196 156081 132224 168898
rect 132276 167596 132328 167602
rect 132276 167538 132328 167544
rect 132288 162026 132316 167538
rect 132552 164808 132604 164814
rect 132552 164750 132604 164756
rect 132276 162020 132328 162026
rect 132276 161962 132328 161968
rect 132274 158112 132330 158121
rect 132274 158047 132330 158056
rect 132182 156072 132238 156081
rect 132182 156007 132238 156016
rect 132090 153624 132146 153633
rect 132090 153559 132146 153568
rect 131906 150904 131962 150913
rect 131906 150839 131962 150848
rect 131816 149576 131868 149582
rect 131816 149518 131868 149524
rect 131630 148864 131686 148873
rect 131630 148799 131686 148808
rect 132288 146794 132316 158047
rect 132458 157160 132514 157169
rect 132458 157095 132514 157104
rect 132366 156344 132422 156353
rect 132366 156279 132422 156288
rect 132276 146788 132328 146794
rect 132276 146730 132328 146736
rect 128136 145428 128188 145434
rect 128136 145370 128188 145376
rect 128044 144884 128096 144890
rect 128044 144826 128096 144832
rect 124272 144816 124324 144822
rect 124272 144758 124324 144764
rect 120684 144748 120736 144754
rect 120684 144690 120736 144696
rect 132380 144074 132408 156279
rect 132472 145434 132500 157095
rect 132564 153361 132592 164750
rect 132644 163516 132696 163522
rect 132644 163458 132696 163464
rect 132550 153352 132606 153361
rect 132550 153287 132606 153296
rect 132656 152273 132684 163458
rect 132642 152264 132698 152273
rect 132642 152199 132698 152208
rect 132460 145428 132512 145434
rect 132460 145370 132512 145376
rect 132368 144068 132420 144074
rect 132368 144010 132420 144016
rect 127584 142028 127636 142034
rect 127584 141970 127636 141976
rect 127596 141354 127624 141970
rect 127216 141348 127268 141354
rect 127216 141290 127268 141296
rect 127584 141348 127636 141354
rect 127584 141290 127636 141296
rect 116176 139512 116228 139518
rect 116176 139454 116228 139460
rect 127228 134434 127256 141290
rect 127228 134406 128084 134434
rect 91086 133726 91284 133754
rect 103506 133726 103704 133754
rect 116018 133726 116124 133754
rect 128056 133618 128084 134406
rect 128056 133590 128530 133618
rect 84710 127512 84766 127521
rect 85828 127482 88156 127498
rect 84710 127447 84712 127456
rect 84764 127447 84766 127456
rect 85816 127476 88156 127482
rect 84712 127418 84764 127424
rect 85868 127470 88156 127476
rect 85816 127418 85868 127424
rect 76892 125504 76944 125510
rect 82688 125504 82740 125510
rect 76892 125446 76944 125452
rect 82686 125472 82688 125481
rect 82740 125472 82742 125481
rect 76904 125102 76932 125446
rect 82686 125407 82742 125416
rect 76892 125096 76944 125102
rect 76892 125038 76944 125044
rect 76800 91504 76852 91510
rect 76800 91446 76852 91452
rect 74038 89840 74094 89849
rect 74038 89775 74094 89784
rect 73856 87424 73908 87430
rect 73856 87366 73908 87372
rect 73672 87220 73724 87226
rect 73672 87162 73724 87168
rect 73578 86304 73634 86313
rect 73578 86239 73634 86248
rect 73684 86177 73712 87162
rect 73868 86449 73896 87366
rect 73854 86440 73910 86449
rect 73854 86375 73910 86384
rect 73486 86168 73542 86177
rect 73486 86103 73542 86112
rect 73670 86168 73726 86177
rect 73670 86103 73726 86112
rect 69360 85990 69572 86018
rect 69360 79134 69388 85990
rect 76904 79202 76932 125038
rect 88128 117842 88156 127470
rect 88128 117814 88340 117842
rect 84710 109832 84766 109841
rect 88312 109818 88340 117814
rect 84710 109767 84712 109776
rect 84764 109767 84766 109776
rect 85816 109796 85868 109802
rect 84712 109738 84764 109744
rect 85816 109738 85868 109744
rect 87208 109790 88432 109818
rect 85828 109682 85856 109738
rect 87208 109682 87236 109790
rect 85828 109654 87236 109682
rect 82596 109524 82648 109530
rect 82596 109466 82648 109472
rect 82608 108889 82636 109466
rect 82594 108880 82650 108889
rect 82594 108815 82650 108824
rect 88404 98530 88432 109790
rect 88220 98502 88432 98530
rect 84802 93512 84858 93521
rect 85828 93482 87420 93498
rect 84802 93447 84804 93456
rect 84856 93447 84858 93456
rect 85816 93476 87420 93482
rect 84804 93418 84856 93424
rect 85868 93470 87420 93476
rect 85816 93418 85868 93424
rect 87392 93226 87420 93470
rect 88220 93362 88248 98502
rect 88128 93334 88248 93362
rect 88128 93226 88156 93334
rect 87392 93198 88156 93226
rect 82688 92728 82740 92734
rect 82688 92670 82740 92676
rect 82700 92297 82728 92670
rect 82686 92288 82742 92297
rect 82686 92223 82742 92232
rect 87392 88738 87420 93198
rect 87392 88710 88432 88738
rect 88404 84386 88432 88710
rect 88220 84358 88432 84386
rect 75788 79196 75840 79202
rect 75788 79138 75840 79144
rect 76892 79196 76944 79202
rect 76892 79138 76944 79144
rect 69348 79128 69400 79134
rect 69348 79070 69400 79076
rect 68520 78924 68572 78930
rect 68520 78866 68572 78872
rect 74776 78856 74828 78862
rect 74776 78798 74828 78804
rect 71648 78788 71700 78794
rect 71648 78730 71700 78736
rect 70636 78652 70688 78658
rect 70636 78594 70688 78600
rect 69624 78584 69676 78590
rect 69624 78526 69676 78532
rect 69636 75804 69664 78526
rect 70648 75804 70676 78594
rect 71660 75804 71688 78730
rect 72660 78720 72712 78726
rect 72660 78662 72712 78668
rect 72672 75804 72700 78662
rect 73764 78516 73816 78522
rect 73764 78458 73816 78464
rect 73776 75804 73804 78458
rect 74788 75804 74816 78798
rect 75800 75804 75828 79138
rect 88220 76482 88248 84358
rect 88418 83814 88524 83842
rect 95502 83814 95792 83842
rect 102678 83814 102968 83842
rect 109762 83814 109868 83842
rect 116938 83814 117136 83842
rect 124022 83814 124128 83842
rect 131198 83814 131304 83842
rect 88496 81990 88524 83814
rect 88484 81984 88536 81990
rect 88484 81926 88536 81932
rect 95764 81922 95792 83814
rect 95752 81916 95804 81922
rect 95752 81858 95804 81864
rect 102940 81854 102968 83814
rect 102928 81848 102980 81854
rect 102928 81790 102980 81796
rect 109840 81310 109868 83814
rect 96764 81304 96816 81310
rect 96764 81246 96816 81252
rect 109828 81304 109880 81310
rect 109828 81246 109880 81252
rect 88024 76476 88076 76482
rect 88024 76418 88076 76424
rect 88208 76476 88260 76482
rect 88208 76418 88260 76424
rect 79468 76408 79520 76414
rect 79468 76350 79520 76356
rect 79480 75841 79508 76350
rect 79466 75832 79522 75841
rect 79466 75767 79522 75776
rect 50040 75654 50974 75682
rect 51512 75654 51986 75682
rect 66692 75654 67534 75682
rect 67888 75654 68546 75682
rect 80202 73928 80258 73937
rect 80202 73863 80258 73872
rect 80216 73762 80244 73863
rect 80204 73756 80256 73762
rect 80204 73698 80256 73704
rect 87932 73756 87984 73762
rect 87932 73698 87984 73704
rect 79834 72840 79890 72849
rect 79834 72775 79890 72784
rect 79848 72402 79876 72775
rect 79836 72396 79888 72402
rect 79836 72338 79888 72344
rect 85724 72396 85776 72402
rect 85724 72338 85776 72344
rect 78914 71616 78970 71625
rect 78914 71551 78970 71560
rect 78928 71042 78956 71551
rect 80202 71208 80258 71217
rect 80258 71166 80336 71194
rect 80202 71143 80258 71152
rect 78916 71036 78968 71042
rect 78916 70978 78968 70984
rect 80202 69848 80258 69857
rect 80202 69783 80258 69792
rect 80216 69614 80244 69783
rect 80204 69608 80256 69614
rect 80204 69550 80256 69556
rect 79282 68624 79338 68633
rect 79282 68559 79338 68568
rect 79296 68254 79324 68559
rect 79284 68248 79336 68254
rect 79284 68190 79336 68196
rect 79560 67568 79612 67574
rect 79560 67510 79612 67516
rect 79466 64544 79522 64553
rect 79466 64479 79468 64488
rect 79520 64479 79522 64488
rect 79468 64450 79520 64456
rect 78914 56112 78970 56121
rect 78914 56047 78970 56056
rect 78928 55810 78956 56047
rect 78916 55804 78968 55810
rect 78916 55746 78968 55752
rect 16356 55736 16408 55742
rect 79572 55713 79600 67510
rect 80202 67400 80258 67409
rect 80202 67335 80258 67344
rect 80216 67234 80244 67335
rect 80204 67228 80256 67234
rect 80204 67170 80256 67176
rect 80202 66856 80258 66865
rect 80202 66791 80204 66800
rect 80256 66791 80258 66800
rect 80204 66762 80256 66768
rect 80308 66758 80336 71166
rect 85632 71036 85684 71042
rect 85632 70978 85684 70984
rect 85080 68248 85132 68254
rect 85080 68190 85132 68196
rect 82780 67228 82832 67234
rect 82780 67170 82832 67176
rect 80296 66752 80348 66758
rect 80296 66694 80348 66700
rect 80202 65632 80258 65641
rect 80202 65567 80258 65576
rect 80216 65466 80244 65567
rect 80204 65460 80256 65466
rect 80204 65402 80256 65408
rect 82792 65398 82820 67170
rect 82780 65392 82832 65398
rect 82780 65334 82832 65340
rect 85092 65330 85120 68190
rect 85644 68186 85672 70978
rect 85736 69002 85764 72338
rect 87288 69608 87340 69614
rect 87288 69550 87340 69556
rect 85724 68996 85776 69002
rect 85724 68938 85776 68944
rect 85632 68180 85684 68186
rect 85632 68122 85684 68128
rect 87196 66752 87248 66758
rect 87194 66720 87196 66729
rect 87248 66720 87250 66729
rect 87194 66655 87250 66664
rect 87300 65913 87328 69550
rect 87944 69449 87972 73698
rect 88036 69562 88064 76418
rect 96776 69834 96804 81246
rect 117108 79354 117136 83814
rect 124100 83706 124128 83814
rect 131276 83706 131304 83814
rect 116924 79326 117136 79354
rect 124008 83678 124128 83706
rect 131092 83678 131304 83706
rect 116924 79218 116952 79326
rect 116832 79190 116952 79218
rect 116832 73490 116860 79190
rect 124008 76414 124036 83678
rect 131092 79218 131120 83678
rect 131000 79190 131120 79218
rect 123996 76408 124048 76414
rect 123996 76350 124048 76356
rect 110196 73484 110248 73490
rect 110196 73426 110248 73432
rect 116820 73484 116872 73490
rect 116820 73426 116872 73432
rect 110208 69834 110236 73426
rect 131000 72402 131028 79190
rect 123536 72396 123588 72402
rect 123536 72338 123588 72344
rect 130988 72396 131040 72402
rect 130988 72338 131040 72344
rect 123548 69834 123576 72338
rect 132552 70968 132604 70974
rect 132552 70910 132604 70916
rect 96560 69806 96804 69834
rect 109900 69806 110236 69834
rect 123240 69806 123576 69834
rect 88036 69534 88248 69562
rect 87930 69440 87986 69449
rect 87930 69375 87986 69384
rect 87656 68996 87708 69002
rect 87656 68938 87708 68944
rect 87668 68497 87696 68938
rect 87654 68488 87710 68497
rect 87654 68423 87710 68432
rect 87840 68180 87892 68186
rect 87840 68122 87892 68128
rect 87852 67681 87880 68122
rect 87838 67672 87894 67681
rect 87838 67607 87894 67616
rect 87380 66820 87432 66826
rect 87380 66762 87432 66768
rect 87286 65904 87342 65913
rect 87286 65839 87342 65848
rect 87288 65460 87340 65466
rect 87288 65402 87340 65408
rect 87196 65392 87248 65398
rect 87196 65334 87248 65340
rect 85080 65324 85132 65330
rect 85080 65266 85132 65272
rect 82412 64508 82464 64514
rect 82412 64450 82464 64456
rect 80202 63320 80258 63329
rect 80202 63255 80258 63264
rect 80216 63018 80244 63255
rect 80204 63012 80256 63018
rect 80204 62954 80256 62960
rect 80202 62912 80258 62921
rect 80202 62847 80258 62856
rect 80216 62746 80244 62847
rect 80204 62740 80256 62746
rect 80204 62682 80256 62688
rect 82424 62610 82452 64450
rect 87208 64145 87236 65334
rect 87194 64136 87250 64145
rect 87194 64071 87250 64080
rect 82596 63012 82648 63018
rect 82596 62954 82648 62960
rect 82412 62604 82464 62610
rect 82412 62546 82464 62552
rect 80202 61416 80258 61425
rect 80202 61351 80204 61360
rect 80256 61351 80258 61360
rect 81676 61380 81728 61386
rect 80204 61322 80256 61328
rect 81676 61322 81728 61328
rect 80202 60192 80258 60201
rect 80202 60127 80204 60136
rect 80256 60127 80258 60136
rect 80204 60098 80256 60104
rect 81688 59550 81716 61322
rect 82608 61250 82636 62954
rect 85724 62740 85776 62746
rect 85724 62682 85776 62688
rect 82596 61244 82648 61250
rect 82596 61186 82648 61192
rect 81768 60156 81820 60162
rect 81768 60098 81820 60104
rect 81676 59544 81728 59550
rect 81676 59486 81728 59492
rect 79650 59104 79706 59113
rect 79650 59039 79706 59048
rect 79664 58666 79692 59039
rect 79652 58660 79704 58666
rect 79652 58602 79704 58608
rect 80204 58592 80256 58598
rect 80202 58560 80204 58569
rect 80256 58560 80258 58569
rect 81780 58530 81808 60098
rect 85736 59754 85764 62682
rect 87196 62604 87248 62610
rect 87196 62546 87248 62552
rect 87208 61425 87236 62546
rect 87300 62377 87328 65402
rect 87392 63193 87420 66762
rect 88220 66758 88248 69534
rect 131356 69540 131408 69546
rect 131356 69482 131408 69488
rect 131368 69449 131396 69482
rect 131816 69472 131868 69478
rect 131354 69440 131410 69449
rect 131816 69414 131868 69420
rect 131354 69375 131410 69384
rect 131828 68497 131856 69414
rect 131814 68488 131870 68497
rect 131814 68423 131870 68432
rect 132368 68180 132420 68186
rect 132368 68122 132420 68128
rect 132380 67681 132408 68122
rect 132366 67672 132422 67681
rect 132366 67607 132422 67616
rect 129424 67568 129476 67574
rect 129424 67510 129476 67516
rect 88208 66752 88260 66758
rect 88208 66694 88260 66700
rect 87472 65324 87524 65330
rect 87472 65266 87524 65272
rect 87484 64961 87512 65266
rect 87470 64952 87526 64961
rect 87470 64887 87526 64896
rect 87378 63184 87434 63193
rect 87378 63119 87434 63128
rect 87286 62368 87342 62377
rect 87286 62303 87342 62312
rect 87194 61416 87250 61425
rect 87194 61351 87250 61360
rect 87196 61244 87248 61250
rect 87196 61186 87248 61192
rect 87208 60473 87236 61186
rect 87194 60464 87250 60473
rect 87194 60399 87250 60408
rect 85724 59748 85776 59754
rect 85724 59690 85776 59696
rect 87840 59748 87892 59754
rect 87840 59690 87892 59696
rect 87852 59657 87880 59690
rect 87838 59648 87894 59657
rect 87838 59583 87894 59592
rect 87196 59544 87248 59550
rect 87196 59486 87248 59492
rect 87208 58705 87236 59486
rect 87194 58696 87250 58705
rect 82964 58660 83016 58666
rect 87194 58631 87250 58640
rect 82964 58602 83016 58608
rect 82412 58592 82464 58598
rect 82412 58534 82464 58540
rect 80202 58495 80258 58504
rect 81768 58524 81820 58530
rect 81768 58466 81820 58472
rect 80202 57200 80258 57209
rect 80202 57135 80204 57144
rect 80256 57135 80258 57144
rect 81860 57164 81912 57170
rect 80204 57106 80256 57112
rect 81860 57106 81912 57112
rect 81872 55742 81900 57106
rect 82424 57034 82452 58534
rect 82976 57102 83004 58602
rect 87196 58524 87248 58530
rect 87196 58466 87248 58472
rect 87208 57889 87236 58466
rect 87194 57880 87250 57889
rect 87194 57815 87250 57824
rect 88300 57164 88352 57170
rect 88300 57106 88352 57112
rect 82964 57096 83016 57102
rect 82964 57038 83016 57044
rect 87196 57096 87248 57102
rect 87196 57038 87248 57044
rect 82412 57028 82464 57034
rect 82412 56970 82464 56976
rect 87208 56937 87236 57038
rect 87288 57028 87340 57034
rect 87288 56970 87340 56976
rect 87194 56928 87250 56937
rect 87194 56863 87250 56872
rect 87300 56121 87328 56970
rect 87286 56112 87342 56121
rect 87286 56047 87342 56056
rect 82964 55804 83016 55810
rect 82964 55746 83016 55752
rect 81860 55736 81912 55742
rect 16356 55678 16408 55684
rect 79558 55704 79614 55713
rect 81860 55678 81912 55684
rect 79558 55639 79614 55648
rect 80202 54616 80258 54625
rect 80202 54551 80258 54560
rect 80216 54450 80244 54551
rect 80204 54444 80256 54450
rect 80204 54386 80256 54392
rect 82976 54314 83004 55746
rect 87196 55736 87248 55742
rect 87196 55678 87248 55684
rect 87208 55169 87236 55678
rect 87194 55160 87250 55169
rect 87194 55095 87250 55104
rect 87194 54344 87250 54353
rect 82964 54308 83016 54314
rect 87194 54279 87196 54288
rect 82964 54250 83016 54256
rect 87248 54279 87250 54288
rect 87196 54250 87248 54256
rect 80204 53696 80256 53702
rect 80202 53664 80204 53673
rect 80256 53664 80258 53673
rect 80202 53599 80258 53608
rect 80204 53016 80256 53022
rect 80204 52958 80256 52964
rect 80216 52721 80244 52958
rect 80202 52712 80258 52721
rect 80202 52647 80258 52656
rect 88312 51526 88340 57106
rect 129436 55062 129464 67510
rect 132368 66752 132420 66758
rect 132564 66729 132592 70910
rect 132368 66694 132420 66700
rect 132550 66720 132606 66729
rect 132380 65913 132408 66694
rect 132550 66655 132606 66664
rect 132366 65904 132422 65913
rect 132366 65839 132422 65848
rect 131356 65392 131408 65398
rect 131356 65334 131408 65340
rect 131368 64961 131396 65334
rect 132184 65324 132236 65330
rect 132184 65266 132236 65272
rect 131354 64952 131410 64961
rect 131354 64887 131410 64896
rect 132196 64145 132224 65266
rect 132182 64136 132238 64145
rect 132182 64071 132238 64080
rect 132368 64032 132420 64038
rect 132368 63974 132420 63980
rect 132380 63193 132408 63974
rect 132366 63184 132422 63193
rect 132366 63119 132422 63128
rect 131724 62604 131776 62610
rect 131724 62546 131776 62552
rect 131356 62536 131408 62542
rect 131356 62478 131408 62484
rect 131368 62377 131396 62478
rect 131354 62368 131410 62377
rect 131354 62303 131410 62312
rect 131736 61425 131764 62546
rect 131722 61416 131778 61425
rect 131722 61351 131778 61360
rect 131356 61244 131408 61250
rect 131356 61186 131408 61192
rect 131368 60473 131396 61186
rect 131354 60464 131410 60473
rect 131354 60399 131410 60408
rect 131356 59884 131408 59890
rect 131356 59826 131408 59832
rect 131368 59657 131396 59826
rect 131448 59816 131500 59822
rect 131448 59758 131500 59764
rect 131354 59648 131410 59657
rect 131354 59583 131410 59592
rect 131460 58705 131488 59758
rect 131446 58696 131502 58705
rect 131446 58631 131502 58640
rect 131356 58524 131408 58530
rect 131356 58466 131408 58472
rect 131368 57889 131396 58466
rect 131354 57880 131410 57889
rect 131354 57815 131410 57824
rect 132184 57096 132236 57102
rect 132184 57038 132236 57044
rect 131356 57028 131408 57034
rect 131356 56970 131408 56976
rect 131368 56937 131396 56970
rect 131354 56928 131410 56937
rect 131354 56863 131410 56872
rect 132196 56121 132224 57038
rect 132182 56112 132238 56121
rect 132182 56047 132238 56056
rect 131356 55736 131408 55742
rect 131356 55678 131408 55684
rect 131368 55169 131396 55678
rect 131354 55160 131410 55169
rect 131354 55095 131410 55104
rect 129424 55056 129476 55062
rect 129424 54998 129476 55004
rect 123536 54172 123588 54178
rect 123536 54114 123588 54120
rect 100424 54030 100484 54058
rect 91040 53894 91284 53922
rect 93340 53894 93676 53922
rect 95732 53894 95792 53922
rect 98032 53894 98092 53922
rect 91256 51594 91284 53894
rect 91244 51588 91296 51594
rect 91244 51530 91296 51536
rect 93648 51526 93676 53894
rect 88300 51520 88352 51526
rect 88300 51462 88352 51468
rect 93636 51520 93688 51526
rect 93636 51462 93688 51468
rect 91244 50908 91296 50914
rect 91244 50850 91296 50856
rect 78914 50808 78970 50817
rect 78914 50743 78970 50752
rect 78928 50370 78956 50743
rect 78916 50364 78968 50370
rect 78916 50306 78968 50312
rect 80204 50296 80256 50302
rect 80202 50264 80204 50273
rect 80256 50264 80258 50273
rect 80202 50199 80258 50208
rect 88392 49548 88444 49554
rect 88392 49490 88444 49496
rect 88404 49321 88432 49490
rect 88390 49312 88446 49321
rect 88390 49247 88446 49256
rect 80202 49176 80258 49185
rect 80202 49111 80258 49120
rect 80216 48942 80244 49111
rect 80204 48936 80256 48942
rect 80204 48878 80256 48884
rect 88298 48632 88354 48641
rect 88298 48567 88354 48576
rect 88312 48097 88340 48567
rect 67874 48088 67930 48097
rect 67718 48046 67874 48074
rect 67874 48023 67930 48032
rect 74314 48088 74370 48097
rect 80202 48088 80258 48097
rect 74370 48060 74710 48074
rect 74370 48046 74724 48060
rect 74314 48023 74370 48032
rect 50224 45746 50252 47924
rect 53720 46018 53748 47924
rect 53708 46012 53760 46018
rect 53708 45954 53760 45960
rect 57216 45950 57244 47924
rect 60712 47446 60740 47924
rect 60700 47440 60752 47446
rect 60700 47382 60752 47388
rect 57204 45944 57256 45950
rect 64208 45921 64236 47924
rect 71214 47910 71504 47938
rect 71476 47417 71504 47910
rect 74224 47440 74276 47446
rect 71462 47408 71518 47417
rect 71462 47343 71518 47352
rect 73118 47408 73174 47417
rect 74224 47382 74276 47388
rect 73118 47343 73174 47352
rect 73132 46222 73160 47343
rect 73120 46216 73172 46222
rect 74236 46193 74264 47382
rect 74696 46834 74724 48046
rect 80202 48023 80258 48032
rect 88298 48088 88354 48097
rect 88298 48023 88354 48032
rect 80216 47718 80244 48023
rect 80204 47712 80256 47718
rect 80204 47654 80256 47660
rect 74684 46828 74736 46834
rect 74684 46770 74736 46776
rect 88116 46828 88168 46834
rect 88116 46770 88168 46776
rect 88024 46760 88076 46766
rect 88024 46702 88076 46708
rect 73120 46158 73172 46164
rect 74222 46184 74278 46193
rect 88036 46154 88064 46702
rect 88128 46154 88156 46770
rect 88208 46216 88260 46222
rect 88208 46158 88260 46164
rect 74222 46119 74224 46128
rect 74276 46119 74278 46128
rect 88024 46148 88076 46154
rect 74224 46090 74276 46096
rect 88024 46090 88076 46096
rect 88116 46148 88168 46154
rect 88116 46090 88168 46096
rect 57204 45886 57256 45892
rect 64194 45912 64250 45921
rect 64194 45847 64250 45856
rect 50212 45740 50264 45746
rect 50212 45682 50264 45688
rect 16264 42612 16316 42618
rect 16264 42554 16316 42560
rect 16172 29488 16224 29494
rect 16172 29430 16224 29436
rect 88036 23345 88064 46090
rect 88128 33681 88156 46090
rect 88114 33672 88170 33681
rect 88114 33607 88170 33616
rect 88220 30825 88248 46158
rect 88206 30816 88262 30825
rect 88206 30751 88262 30760
rect 88312 28105 88340 48023
rect 88298 28096 88354 28105
rect 88298 28031 88354 28040
rect 88404 26065 88432 49247
rect 91256 34746 91284 50850
rect 93648 50681 93676 51462
rect 93634 50672 93690 50681
rect 93634 50607 93690 50616
rect 93728 47576 93780 47582
rect 93648 47536 93728 47564
rect 93648 34746 93676 47536
rect 93728 47518 93780 47524
rect 95476 46012 95528 46018
rect 95476 45954 95528 45960
rect 95488 45882 95516 45954
rect 95764 45882 95792 53894
rect 96764 48528 96816 48534
rect 96764 48470 96816 48476
rect 95476 45876 95528 45882
rect 95476 45818 95528 45824
rect 95752 45876 95804 45882
rect 95752 45818 95804 45824
rect 96776 37518 96804 48470
rect 98064 45950 98092 53894
rect 98604 48936 98656 48942
rect 98604 48878 98656 48884
rect 98052 45944 98104 45950
rect 98052 45886 98104 45892
rect 96396 37512 96448 37518
rect 96396 37454 96448 37460
rect 96764 37512 96816 37518
rect 96764 37454 96816 37460
rect 96408 34746 96436 37454
rect 98616 34746 98644 48878
rect 100456 47514 100484 54030
rect 102388 53894 102724 53922
rect 105116 53894 105176 53922
rect 107508 53894 107568 53922
rect 102388 51361 102416 53894
rect 102374 51352 102430 51361
rect 102374 51287 102430 51296
rect 102284 51044 102336 51050
rect 102284 50986 102336 50992
rect 100260 47508 100312 47514
rect 100260 47450 100312 47456
rect 100444 47508 100496 47514
rect 100444 47450 100496 47456
rect 100272 46766 100300 47450
rect 100260 46760 100312 46766
rect 100260 46702 100312 46708
rect 102296 37790 102324 50986
rect 102388 49554 102416 51287
rect 103572 50296 103624 50302
rect 103572 50238 103624 50244
rect 102376 49548 102428 49554
rect 102376 49490 102428 49496
rect 101364 37784 101416 37790
rect 101364 37726 101416 37732
rect 102284 37784 102336 37790
rect 102284 37726 102336 37732
rect 101376 34746 101404 37726
rect 103584 34746 103612 50238
rect 105148 49321 105176 53894
rect 106424 51112 106476 51118
rect 106424 51054 106476 51060
rect 105134 49312 105190 49321
rect 105134 49247 105190 49256
rect 105148 48097 105176 49247
rect 105134 48088 105190 48097
rect 105134 48023 105190 48032
rect 106436 34746 106464 51054
rect 107540 50273 107568 53894
rect 109472 53894 109808 53922
rect 112048 53894 112200 53922
rect 114164 53894 114500 53922
rect 116556 53894 116892 53922
rect 119132 53894 119284 53922
rect 121248 53894 121584 53922
rect 108632 50364 108684 50370
rect 108632 50306 108684 50312
rect 107526 50264 107582 50273
rect 107526 50199 107582 50208
rect 106606 47408 106662 47417
rect 106606 47343 106662 47352
rect 106620 46222 106648 47343
rect 106608 46216 106660 46222
rect 106608 46158 106660 46164
rect 108644 34746 108672 50306
rect 109472 50273 109500 53894
rect 111944 51180 111996 51186
rect 111944 51122 111996 51128
rect 109458 50264 109514 50273
rect 109458 50199 109514 50208
rect 109458 47272 109514 47281
rect 109458 47207 109514 47216
rect 109472 46154 109500 47207
rect 109460 46148 109512 46154
rect 109460 46090 109512 46096
rect 111956 36702 111984 51122
rect 112048 50914 112076 53894
rect 113966 53120 114022 53129
rect 113966 53055 114022 53064
rect 113980 53022 114008 53055
rect 113968 53016 114020 53022
rect 113968 52958 114020 52964
rect 114164 50982 114192 53894
rect 116556 51050 116584 53894
rect 118660 53696 118712 53702
rect 118660 53638 118712 53644
rect 118672 53129 118700 53638
rect 118658 53120 118714 53129
rect 118658 53055 118714 53064
rect 119132 51118 119160 53894
rect 121248 51186 121276 53894
rect 121236 51180 121288 51186
rect 121236 51122 121288 51128
rect 119120 51112 119172 51118
rect 119120 51054 119172 51060
rect 116544 51044 116596 51050
rect 116544 50986 116596 50992
rect 114152 50976 114204 50982
rect 114152 50918 114204 50924
rect 112036 50908 112088 50914
rect 112036 50850 112088 50856
rect 116084 50908 116136 50914
rect 116084 50850 116136 50856
rect 113598 43328 113654 43337
rect 113598 43263 113654 43272
rect 111392 36696 111444 36702
rect 111392 36638 111444 36644
rect 111944 36696 111996 36702
rect 111944 36638 111996 36644
rect 111404 34746 111432 36638
rect 113612 34746 113640 43263
rect 116096 34746 116124 50850
rect 123548 50794 123576 54114
rect 123640 53894 123976 53922
rect 125940 53894 126276 53922
rect 128668 53894 128728 53922
rect 123640 50914 123668 53894
rect 125940 51322 125968 53894
rect 125100 51316 125152 51322
rect 125100 51258 125152 51264
rect 125928 51316 125980 51322
rect 125928 51258 125980 51264
rect 123628 50908 123680 50914
rect 123628 50850 123680 50856
rect 123548 50766 123760 50794
rect 123732 50114 123760 50766
rect 123732 50086 123852 50114
rect 118658 46184 118714 46193
rect 118658 46119 118714 46128
rect 118672 34746 118700 46119
rect 121420 37172 121472 37178
rect 121420 37114 121472 37120
rect 121432 34746 121460 37114
rect 123824 34746 123852 50086
rect 125112 37178 125140 51258
rect 128700 50438 128728 53894
rect 127124 50432 127176 50438
rect 127124 50374 127176 50380
rect 128688 50432 128740 50438
rect 128688 50374 128740 50380
rect 125100 37172 125152 37178
rect 125100 37114 125152 37120
rect 127136 36634 127164 50374
rect 129436 40730 129464 54998
rect 134116 54444 134168 54450
rect 134116 54386 134168 54392
rect 131356 54376 131408 54382
rect 131354 54344 131356 54353
rect 131408 54344 131410 54353
rect 134128 54314 134156 54386
rect 131354 54279 131410 54288
rect 134116 54308 134168 54314
rect 134116 54250 134168 54256
rect 134772 51594 134800 225474
rect 136888 213881 136916 235023
rect 136966 234952 137022 234961
rect 136966 234887 137022 234896
rect 136874 213872 136930 213881
rect 136874 213807 136930 213816
rect 136980 210753 137008 234887
rect 137072 217009 137100 235198
rect 137152 233148 137204 233154
rect 137152 233090 137204 233096
rect 137164 220137 137192 233090
rect 137256 226393 137284 235266
rect 137336 234440 137388 234446
rect 137336 234382 137388 234388
rect 137348 234281 137376 234382
rect 137334 234272 137390 234281
rect 137334 234207 137390 234216
rect 137242 226384 137298 226393
rect 137242 226319 137298 226328
rect 137348 223265 137376 234207
rect 137624 226150 137652 285207
rect 137716 279705 137744 309658
rect 137808 301601 137836 327406
rect 137900 320369 137928 328970
rect 137886 320360 137942 320369
rect 137886 320295 137942 320304
rect 137794 301592 137850 301601
rect 137794 301527 137850 301536
rect 137796 295912 137848 295918
rect 137796 295854 137848 295860
rect 137702 279696 137758 279705
rect 137702 279631 137758 279640
rect 137808 276577 137836 295854
rect 137888 283536 137940 283542
rect 137888 283478 137940 283484
rect 137794 276568 137850 276577
rect 137794 276503 137850 276512
rect 137900 273449 137928 283478
rect 142408 283406 142436 329838
rect 144616 326722 144644 329838
rect 144604 326716 144656 326722
rect 144604 326658 144656 326664
rect 145536 326382 145564 329838
rect 145904 329838 146240 329866
rect 147160 329838 147496 329866
rect 148172 329838 148508 329866
rect 145524 326376 145576 326382
rect 145524 326318 145576 326324
rect 145904 326314 145932 329838
rect 147468 326654 147496 329838
rect 147456 326648 147508 326654
rect 147456 326590 147508 326596
rect 148480 326586 148508 329838
rect 148756 329838 149092 329866
rect 150104 329838 150440 329866
rect 151024 329838 151360 329866
rect 152036 329838 152188 329866
rect 152956 329838 153292 329866
rect 153968 329838 154304 329866
rect 148468 326580 148520 326586
rect 148468 326522 148520 326528
rect 148756 326314 148784 329838
rect 149388 327260 149440 327266
rect 149388 327202 149440 327208
rect 145340 326308 145392 326314
rect 145340 326250 145392 326256
rect 145892 326308 145944 326314
rect 145892 326250 145944 326256
rect 147916 326308 147968 326314
rect 147916 326250 147968 326256
rect 148744 326308 148796 326314
rect 148744 326250 148796 326256
rect 145352 319990 145380 326250
rect 147928 320058 147956 326250
rect 149296 320120 149348 320126
rect 149296 320062 149348 320068
rect 147916 320052 147968 320058
rect 147916 319994 147968 320000
rect 145340 319984 145392 319990
rect 145340 319926 145392 319932
rect 149308 316796 149336 320062
rect 149400 316946 149428 327202
rect 150412 326518 150440 329838
rect 150860 327328 150912 327334
rect 150860 327270 150912 327276
rect 150768 327056 150820 327062
rect 150768 326998 150820 327004
rect 150400 326512 150452 326518
rect 150400 326454 150452 326460
rect 149400 316918 149796 316946
rect 149768 316810 149796 316918
rect 150780 316810 150808 326998
rect 150872 320670 150900 327270
rect 151332 326314 151360 329838
rect 152160 326450 152188 329838
rect 152240 327192 152292 327198
rect 152240 327134 152292 327140
rect 152148 326444 152200 326450
rect 152148 326386 152200 326392
rect 151320 326308 151372 326314
rect 151320 326250 151372 326256
rect 150860 320664 150912 320670
rect 150860 320606 150912 320612
rect 151964 320664 152016 320670
rect 151964 320606 152016 320612
rect 149768 316782 150150 316810
rect 150780 316782 151070 316810
rect 151976 316796 152004 320606
rect 152252 316946 152280 327134
rect 152332 326376 152384 326382
rect 153264 326353 153292 329838
rect 154080 327124 154132 327130
rect 154080 327066 154132 327072
rect 153528 326784 153580 326790
rect 153528 326726 153580 326732
rect 152332 326318 152384 326324
rect 153250 326344 153306 326353
rect 152344 319514 152372 326318
rect 153250 326279 153306 326288
rect 152332 319508 152384 319514
rect 152332 319450 152384 319456
rect 152252 316918 152464 316946
rect 152436 316810 152464 316918
rect 153540 316810 153568 326726
rect 152436 316782 152818 316810
rect 153540 316782 153738 316810
rect 154092 316674 154120 327066
rect 154276 326926 154304 329838
rect 154874 329594 154902 329852
rect 154828 329566 154902 329594
rect 154828 327402 154856 329566
rect 155932 327470 155960 329974
rect 155920 327464 155972 327470
rect 155920 327406 155972 327412
rect 154816 327396 154868 327402
rect 154816 327338 154868 327344
rect 154828 326994 154856 327338
rect 154816 326988 154868 326994
rect 154816 326930 154868 326936
rect 156288 326988 156340 326994
rect 156288 326930 156340 326936
rect 154264 326920 154316 326926
rect 154264 326862 154316 326868
rect 154908 326852 154960 326858
rect 154908 326794 154960 326800
rect 154816 326308 154868 326314
rect 154816 326250 154868 326256
rect 154828 320602 154856 326250
rect 154816 320596 154868 320602
rect 154816 320538 154868 320544
rect 154920 316810 154948 326794
rect 156196 326716 156248 326722
rect 156196 326658 156248 326664
rect 155644 326308 155696 326314
rect 155644 326250 155696 326256
rect 155656 320126 155684 326250
rect 156208 320670 156236 326658
rect 156196 320664 156248 320670
rect 156196 320606 156248 320612
rect 155644 320120 155696 320126
rect 155644 320062 155696 320068
rect 156300 316810 156328 326930
rect 156852 326382 156880 329974
rect 157832 329838 158168 329866
rect 158140 327441 158168 329838
rect 158416 329838 158752 329866
rect 160684 329838 161020 329866
rect 161696 329838 161756 329866
rect 158416 327538 158444 329838
rect 160992 327606 161020 329838
rect 161728 329481 161756 329838
rect 162280 329838 162616 329866
rect 163292 329838 163628 329866
rect 164548 329838 164608 329866
rect 161714 329472 161770 329481
rect 161714 329407 161770 329416
rect 161728 329034 161756 329407
rect 161716 329028 161768 329034
rect 161716 328970 161768 328976
rect 160980 327600 161032 327606
rect 160980 327542 161032 327548
rect 158404 327532 158456 327538
rect 158404 327474 158456 327480
rect 158126 327432 158182 327441
rect 158126 327367 158182 327376
rect 159048 326648 159100 326654
rect 159048 326590 159100 326596
rect 158956 326512 159008 326518
rect 158956 326454 159008 326460
rect 156840 326376 156892 326382
rect 156840 326318 156892 326324
rect 158968 320670 158996 326454
rect 156932 320664 156984 320670
rect 156932 320606 156984 320612
rect 158956 320664 159008 320670
rect 158956 320606 159008 320612
rect 156944 316810 156972 320606
rect 159060 320074 159088 326590
rect 160244 326580 160296 326586
rect 160244 326522 160296 326528
rect 159060 320046 159456 320074
rect 159048 319984 159100 319990
rect 159048 319926 159100 319932
rect 158128 319508 158180 319514
rect 158128 319450 158180 319456
rect 154920 316782 155486 316810
rect 156300 316782 156406 316810
rect 156944 316782 157326 316810
rect 158140 316796 158168 319450
rect 159060 316796 159088 319926
rect 159428 316674 159456 320046
rect 160256 319394 160284 326522
rect 162280 326314 162308 329838
rect 163292 327266 163320 329838
rect 163280 327260 163332 327266
rect 163280 327202 163332 327208
rect 164580 327062 164608 329838
rect 165224 329838 165560 329866
rect 166144 329838 166480 329866
rect 167340 329838 167492 329866
rect 168076 329838 168412 329866
rect 169088 329838 169424 329866
rect 170008 329838 170344 329866
rect 165224 327334 165252 329838
rect 165212 327328 165264 327334
rect 165212 327270 165264 327276
rect 166144 327198 166172 329838
rect 166132 327192 166184 327198
rect 166132 327134 166184 327140
rect 164568 327056 164620 327062
rect 164568 326998 164620 327004
rect 167340 326790 167368 329838
rect 168076 327130 168104 329838
rect 168064 327124 168116 327130
rect 168064 327066 168116 327072
rect 169088 326858 169116 329838
rect 170008 326994 170036 329838
rect 173412 329102 173440 330223
rect 173400 329096 173452 329102
rect 173400 329038 173452 329044
rect 169996 326988 170048 326994
rect 169996 326930 170048 326936
rect 169076 326852 169128 326858
rect 169076 326794 169128 326800
rect 167328 326784 167380 326790
rect 167328 326726 167380 326732
rect 163004 326444 163056 326450
rect 163004 326386 163056 326392
rect 162268 326308 162320 326314
rect 162268 326250 162320 326256
rect 162636 320664 162688 320670
rect 162636 320606 162688 320612
rect 161716 320052 161768 320058
rect 161716 319994 161768 320000
rect 160256 319366 160376 319394
rect 160348 316810 160376 319366
rect 160348 316782 160822 316810
rect 161728 316796 161756 319994
rect 162648 316796 162676 320606
rect 163016 319990 163044 326386
rect 185096 321692 185124 333798
rect 185924 333794 185952 335822
rect 185912 333788 185964 333794
rect 185912 333730 185964 333736
rect 187948 327402 187976 335958
rect 192088 327470 192116 335958
rect 192076 327464 192128 327470
rect 192076 327406 192128 327412
rect 187936 327396 187988 327402
rect 187936 327338 187988 327344
rect 189224 327396 189276 327402
rect 189224 327338 189276 327344
rect 189236 326994 189264 327338
rect 192088 327062 192116 327406
rect 194848 327130 194876 335958
rect 197504 333924 197556 333930
rect 197504 333866 197556 333872
rect 194836 327124 194888 327130
rect 194836 327066 194888 327072
rect 192076 327056 192128 327062
rect 192076 326998 192128 327004
rect 189224 326988 189276 326994
rect 189224 326930 189276 326936
rect 194848 326314 194876 327066
rect 194836 326308 194888 326314
rect 194836 326250 194888 326256
rect 197516 321692 197544 333866
rect 198804 332978 198832 335958
rect 202222 335822 202512 335850
rect 205534 335822 205640 335850
rect 208846 335822 209320 335850
rect 212250 335822 212356 335850
rect 215562 335822 215668 335850
rect 202484 334474 202512 335822
rect 202472 334468 202524 334474
rect 202472 334410 202524 334416
rect 198792 332972 198844 332978
rect 198792 332914 198844 332920
rect 198804 332201 198832 332914
rect 198790 332192 198846 332201
rect 198790 332127 198846 332136
rect 205612 331657 205640 335822
rect 205598 331648 205654 331657
rect 205598 331583 205654 331592
rect 209292 328966 209320 335822
rect 212328 334406 212356 335822
rect 212316 334400 212368 334406
rect 212316 334342 212368 334348
rect 211304 333992 211356 333998
rect 211304 333934 211356 333940
rect 209280 328960 209332 328966
rect 209280 328902 209332 328908
rect 209292 327606 209320 328902
rect 209280 327600 209332 327606
rect 209280 327542 209332 327548
rect 211316 324206 211344 333934
rect 212328 333561 212356 334342
rect 215640 333862 215668 335822
rect 218584 333930 218612 335958
rect 221896 333998 221924 335958
rect 225208 334406 225236 384759
rect 226484 382816 226536 382822
rect 226482 382784 226484 382793
rect 227220 382816 227272 382822
rect 226536 382784 226538 382793
rect 227220 382758 227272 382764
rect 226482 382719 226538 382728
rect 225286 380200 225342 380209
rect 225286 380135 225342 380144
rect 225196 334400 225248 334406
rect 225196 334342 225248 334348
rect 221884 333992 221936 333998
rect 221884 333934 221936 333940
rect 218572 333924 218624 333930
rect 218572 333866 218624 333872
rect 215628 333856 215680 333862
rect 215628 333798 215680 333804
rect 225208 333590 225236 334342
rect 225196 333584 225248 333590
rect 212314 333552 212370 333561
rect 225196 333526 225248 333532
rect 212314 333487 212370 333496
rect 225300 331657 225328 380135
rect 225378 377480 225434 377489
rect 225378 377415 225434 377424
rect 225392 334474 225420 377415
rect 226484 375200 226536 375206
rect 226484 375142 226536 375148
rect 226496 374769 226524 375142
rect 226482 374760 226538 374769
rect 226482 374695 226538 374704
rect 225838 372176 225894 372185
rect 225838 372111 225894 372120
rect 225852 371806 225880 372111
rect 225840 371800 225892 371806
rect 225840 371742 225892 371748
rect 226298 351368 226354 351377
rect 226298 351303 226300 351312
rect 226352 351303 226354 351312
rect 226300 351274 226352 351280
rect 226390 350416 226446 350425
rect 226390 350351 226446 350360
rect 226404 349774 226432 350351
rect 226392 349768 226444 349774
rect 226392 349710 226444 349716
rect 226482 349600 226538 349609
rect 226482 349535 226538 349544
rect 226390 348648 226446 348657
rect 226390 348583 226446 348592
rect 226404 348414 226432 348583
rect 226392 348408 226444 348414
rect 226392 348350 226444 348356
rect 226496 348346 226524 349535
rect 226484 348340 226536 348346
rect 226484 348282 226536 348288
rect 226390 347832 226446 347841
rect 226390 347767 226446 347776
rect 226404 346986 226432 347767
rect 226392 346980 226444 346986
rect 226392 346922 226444 346928
rect 226298 346880 226354 346889
rect 226298 346815 226354 346824
rect 226312 345694 226340 346815
rect 226390 346064 226446 346073
rect 226390 345999 226446 346008
rect 226300 345688 226352 345694
rect 226300 345630 226352 345636
rect 226404 345626 226432 345999
rect 226392 345620 226444 345626
rect 226392 345562 226444 345568
rect 226482 345112 226538 345121
rect 226482 345047 226538 345056
rect 226390 344296 226446 344305
rect 226496 344266 226524 345047
rect 226390 344231 226446 344240
rect 226484 344260 226536 344266
rect 226404 344198 226432 344231
rect 226484 344202 226536 344208
rect 226392 344192 226444 344198
rect 226392 344134 226444 344140
rect 226390 343344 226446 343353
rect 226390 343279 226446 343288
rect 226404 342838 226432 343279
rect 226392 342832 226444 342838
rect 226392 342774 226444 342780
rect 226482 342392 226538 342401
rect 226482 342327 226538 342336
rect 226390 341576 226446 341585
rect 226496 341546 226524 342327
rect 226390 341511 226446 341520
rect 226484 341540 226536 341546
rect 226404 341478 226432 341511
rect 226484 341482 226536 341488
rect 226392 341472 226444 341478
rect 226392 341414 226444 341420
rect 226390 340624 226446 340633
rect 226390 340559 226446 340568
rect 226404 340118 226432 340559
rect 226392 340112 226444 340118
rect 226392 340054 226444 340060
rect 226482 339808 226538 339817
rect 226482 339743 226538 339752
rect 226390 338856 226446 338865
rect 226390 338791 226446 338800
rect 226404 338690 226432 338791
rect 226496 338758 226524 339743
rect 226484 338752 226536 338758
rect 226484 338694 226536 338700
rect 226392 338684 226444 338690
rect 226392 338626 226444 338632
rect 226390 338040 226446 338049
rect 226390 337975 226446 337984
rect 226404 337670 226432 337975
rect 226392 337664 226444 337670
rect 226392 337606 226444 337612
rect 226390 337088 226446 337097
rect 226390 337023 226446 337032
rect 226404 335970 226432 337023
rect 226574 336272 226630 336281
rect 226574 336207 226630 336216
rect 226392 335964 226444 335970
rect 226392 335906 226444 335912
rect 225380 334468 225432 334474
rect 225380 334410 225432 334416
rect 225392 333182 225420 334410
rect 225380 333176 225432 333182
rect 225380 333118 225432 333124
rect 226588 331754 226616 336207
rect 226576 331748 226628 331754
rect 226576 331690 226628 331696
rect 225286 331648 225342 331657
rect 225286 331583 225342 331592
rect 225300 330666 225328 331583
rect 225288 330660 225340 330666
rect 225288 330602 225340 330608
rect 222528 329232 222580 329238
rect 222528 329174 222580 329180
rect 210016 324200 210068 324206
rect 210016 324142 210068 324148
rect 211304 324200 211356 324206
rect 211304 324142 211356 324148
rect 210028 321692 210056 324142
rect 222540 321692 222568 329174
rect 227232 328966 227260 382758
rect 228416 346980 228468 346986
rect 228416 346922 228468 346928
rect 227956 345688 228008 345694
rect 227956 345630 228008 345636
rect 227968 344130 227996 345630
rect 228428 345558 228456 346922
rect 228416 345552 228468 345558
rect 228416 345494 228468 345500
rect 227956 344124 228008 344130
rect 227956 344066 228008 344072
rect 227220 328960 227272 328966
rect 227220 328902 227272 328908
rect 163464 320596 163516 320602
rect 163464 320538 163516 320544
rect 163004 319984 163056 319990
rect 163004 319926 163056 319932
rect 163476 316796 163504 320538
rect 164384 319984 164436 319990
rect 164384 319926 164436 319932
rect 164396 316796 164424 319926
rect 154092 316646 154658 316674
rect 159428 316646 159994 316674
rect 165118 315872 165174 315881
rect 165118 315807 165174 315816
rect 165132 313122 165160 315807
rect 175514 313560 175570 313569
rect 175514 313495 175570 313504
rect 175528 313122 175556 313495
rect 165120 313116 165172 313122
rect 165120 313058 165172 313064
rect 175516 313116 175568 313122
rect 175516 313058 175568 313064
rect 145522 310160 145578 310169
rect 145522 310095 145578 310104
rect 145536 309722 145564 310095
rect 145524 309716 145576 309722
rect 145524 309658 145576 309664
rect 145430 296832 145486 296841
rect 145430 296767 145486 296776
rect 145444 295918 145472 296767
rect 145432 295912 145484 295918
rect 145432 295854 145484 295860
rect 145156 283536 145208 283542
rect 145154 283504 145156 283513
rect 145208 283504 145210 283513
rect 145154 283439 145210 283448
rect 142396 283400 142448 283406
rect 142396 283342 142448 283348
rect 143040 283400 143092 283406
rect 143040 283342 143092 283348
rect 138162 282552 138218 282561
rect 138162 282487 138218 282496
rect 138176 282386 138204 282487
rect 143052 282386 143080 283342
rect 138164 282380 138216 282386
rect 138164 282322 138216 282328
rect 143040 282380 143092 282386
rect 143040 282322 143092 282328
rect 138438 279288 138494 279297
rect 138438 279223 138494 279232
rect 138452 275110 138480 279223
rect 138440 275104 138492 275110
rect 138440 275046 138492 275052
rect 137886 273440 137942 273449
rect 137886 273375 137942 273384
rect 138452 269913 138480 275046
rect 138438 269904 138494 269913
rect 138438 269839 138494 269848
rect 143052 266542 143080 282322
rect 149216 275042 149244 276948
rect 149204 275036 149256 275042
rect 149204 274978 149256 274984
rect 149768 274974 149796 276948
rect 150426 276934 150532 276962
rect 149756 274968 149808 274974
rect 149756 274910 149808 274916
rect 149204 274764 149256 274770
rect 149204 274706 149256 274712
rect 147824 274696 147876 274702
rect 147824 274638 147876 274644
rect 145064 274628 145116 274634
rect 145064 274570 145116 274576
rect 143684 274492 143736 274498
rect 143684 274434 143736 274440
rect 143040 266536 143092 266542
rect 143040 266478 143092 266484
rect 143696 263770 143724 274434
rect 145076 263770 145104 274570
rect 146444 274560 146496 274566
rect 146444 274502 146496 274508
rect 146456 263770 146484 274502
rect 147836 263770 147864 274638
rect 149216 263770 149244 274706
rect 150504 266610 150532 276934
rect 150584 274900 150636 274906
rect 150584 274842 150636 274848
rect 150492 266604 150544 266610
rect 150492 266546 150544 266552
rect 150596 263770 150624 274842
rect 151056 273886 151084 276948
rect 151622 276934 151820 276962
rect 151044 273880 151096 273886
rect 151044 273822 151096 273828
rect 151792 266406 151820 276934
rect 151872 274832 151924 274838
rect 151872 274774 151924 274780
rect 151780 266400 151832 266406
rect 151780 266342 151832 266348
rect 151884 264042 151912 274774
rect 151964 273880 152016 273886
rect 151964 273822 152016 273828
rect 151976 266678 152004 273822
rect 152252 273818 152280 276948
rect 152910 276934 153384 276962
rect 152240 273812 152292 273818
rect 152240 273754 152292 273760
rect 153252 273812 153304 273818
rect 153252 273754 153304 273760
rect 153160 266808 153212 266814
rect 153160 266750 153212 266756
rect 151964 266672 152016 266678
rect 151964 266614 152016 266620
rect 151884 264014 151958 264042
rect 143572 263742 143724 263770
rect 144952 263742 145104 263770
rect 146332 263742 146484 263770
rect 147712 263742 147864 263770
rect 149092 263742 149244 263770
rect 150564 263742 150624 263770
rect 151930 263756 151958 264014
rect 153172 263770 153200 266750
rect 153264 266474 153292 273754
rect 153356 266898 153384 276934
rect 153448 273818 153476 276948
rect 154106 276934 154672 276962
rect 153436 273812 153488 273818
rect 153436 273754 153488 273760
rect 154644 268122 154672 276934
rect 154736 273857 154764 276948
rect 155288 275110 155316 276948
rect 155932 275178 155960 276948
rect 155920 275172 155972 275178
rect 155920 275114 155972 275120
rect 155276 275104 155328 275110
rect 155276 275046 155328 275052
rect 156576 274401 156604 276948
rect 157220 274537 157248 276948
rect 157772 274809 157800 276948
rect 158220 275036 158272 275042
rect 158220 274978 158272 274984
rect 157758 274800 157814 274809
rect 157758 274735 157814 274744
rect 157206 274528 157262 274537
rect 157206 274463 157262 274472
rect 156562 274392 156618 274401
rect 156562 274327 156618 274336
rect 154722 273848 154778 273857
rect 154722 273783 154778 273792
rect 154724 273744 154776 273750
rect 154724 273686 154776 273692
rect 154552 268094 154672 268122
rect 153356 266870 153476 266898
rect 153448 266762 153476 266870
rect 153356 266734 153476 266762
rect 153252 266468 153304 266474
rect 153252 266410 153304 266416
rect 153356 266270 153384 266734
rect 153344 266264 153396 266270
rect 153344 266206 153396 266212
rect 154552 266202 154580 268094
rect 154736 267986 154764 273686
rect 154644 267958 154764 267986
rect 154644 266338 154672 267958
rect 158232 266882 158260 274978
rect 158416 274673 158444 276948
rect 159060 274945 159088 276948
rect 159046 274936 159102 274945
rect 159046 274871 159102 274880
rect 158402 274664 158458 274673
rect 158402 274599 158458 274608
rect 159612 274498 159640 276948
rect 160256 274634 160284 276948
rect 160520 274968 160572 274974
rect 160520 274910 160572 274916
rect 160244 274628 160296 274634
rect 160244 274570 160296 274576
rect 159600 274492 159652 274498
rect 159600 274434 159652 274440
rect 158220 266876 158272 266882
rect 158220 266818 158272 266824
rect 158956 266876 159008 266882
rect 158956 266818 159008 266824
rect 154724 266740 154776 266746
rect 154724 266682 154776 266688
rect 154632 266332 154684 266338
rect 154632 266274 154684 266280
rect 154540 266196 154592 266202
rect 154540 266138 154592 266144
rect 154736 263770 154764 266682
rect 155736 266536 155788 266542
rect 155736 266478 155788 266484
rect 153172 263742 153324 263770
rect 154704 263742 154764 263770
rect 155748 263770 155776 266478
rect 157852 265720 157904 265726
rect 157852 265662 157904 265668
rect 157864 263770 157892 265662
rect 158968 263770 158996 266818
rect 160532 263770 160560 274910
rect 160900 274566 160928 276948
rect 161452 274702 161480 276948
rect 162096 274770 162124 276948
rect 162740 274906 162768 276948
rect 162728 274900 162780 274906
rect 162728 274842 162780 274848
rect 163292 274838 163320 276948
rect 163280 274832 163332 274838
rect 163280 274774 163332 274780
rect 162084 274764 162136 274770
rect 162084 274706 162136 274712
rect 161440 274696 161492 274702
rect 161440 274638 161492 274644
rect 160888 274560 160940 274566
rect 160888 274502 160940 274508
rect 163936 273818 163964 276948
rect 164488 276934 164594 276962
rect 162360 273812 162412 273818
rect 162360 273754 162412 273760
rect 163924 273812 163976 273818
rect 163924 273754 163976 273760
rect 162372 266814 162400 273754
rect 162360 266808 162412 266814
rect 162360 266750 162412 266756
rect 164488 266746 164516 276934
rect 164476 266740 164528 266746
rect 164476 266682 164528 266688
rect 161716 266672 161768 266678
rect 161716 266614 161768 266620
rect 161728 263770 161756 266614
rect 164568 266400 164620 266406
rect 164568 266342 164620 266348
rect 163096 266128 163148 266134
rect 163096 266070 163148 266076
rect 163108 263770 163136 266070
rect 164580 263770 164608 266342
rect 165132 265726 165160 313058
rect 167878 306216 167934 306225
rect 167878 306151 167934 306160
rect 167892 297210 167920 306151
rect 167880 297204 167932 297210
rect 167880 297146 167932 297152
rect 175516 297204 175568 297210
rect 175516 297146 175568 297152
rect 175528 296841 175556 297146
rect 175514 296832 175570 296841
rect 175514 296767 175570 296776
rect 168062 286360 168118 286369
rect 168062 286295 168118 286304
rect 168076 286262 168104 286295
rect 168064 286256 168116 286262
rect 168064 286198 168116 286204
rect 175424 286256 175476 286262
rect 175424 286198 175476 286204
rect 175436 280249 175464 286198
rect 175422 280240 175478 280249
rect 175422 280175 175478 280184
rect 182428 269670 182456 271916
rect 189512 270162 189540 271916
rect 189420 270134 189540 270162
rect 182416 269664 182468 269670
rect 182416 269606 182468 269612
rect 182968 269664 183020 269670
rect 182968 269606 183020 269612
rect 182980 269505 183008 269606
rect 189420 269534 189448 270134
rect 196688 269602 196716 271916
rect 196676 269596 196728 269602
rect 196676 269538 196728 269544
rect 189408 269528 189460 269534
rect 182966 269496 183022 269505
rect 189408 269470 189460 269476
rect 182966 269431 183022 269440
rect 189316 269052 189368 269058
rect 189316 268994 189368 269000
rect 170640 268984 170692 268990
rect 170640 268926 170692 268932
rect 165948 266468 166000 266474
rect 165948 266410 166000 266416
rect 165120 265720 165172 265726
rect 165120 265662 165172 265668
rect 165960 263770 165988 266410
rect 168708 266332 168760 266338
rect 168708 266274 168760 266280
rect 167328 266264 167380 266270
rect 167328 266206 167380 266212
rect 167340 263770 167368 266206
rect 168720 263770 168748 266274
rect 170088 266196 170140 266202
rect 170088 266138 170140 266144
rect 170100 263770 170128 266138
rect 155748 263742 156084 263770
rect 157556 263742 157892 263770
rect 158936 263742 158996 263770
rect 160316 263742 160560 263770
rect 161696 263742 161756 263770
rect 163076 263742 163136 263770
rect 164548 263742 164608 263770
rect 165928 263742 165988 263770
rect 167308 263742 167368 263770
rect 168688 263742 168748 263770
rect 170068 263742 170128 263770
rect 140280 263476 140332 263482
rect 140280 263418 140332 263424
rect 139818 263104 139874 263113
rect 139818 263039 139874 263048
rect 139832 262802 139860 263039
rect 139820 262796 139872 262802
rect 139820 262738 139872 262744
rect 138806 259976 138862 259985
rect 138806 259911 138862 259920
rect 137704 253208 137756 253214
rect 137704 253150 137756 253156
rect 137716 244782 137744 253150
rect 138820 250601 138848 259911
rect 139728 255928 139780 255934
rect 139728 255870 139780 255876
rect 138992 251848 139044 251854
rect 138992 251790 139044 251796
rect 138806 250592 138862 250601
rect 138806 250527 138862 250536
rect 138900 248992 138952 248998
rect 138900 248934 138952 248940
rect 138438 245560 138494 245569
rect 138438 245495 138494 245504
rect 137704 244776 137756 244782
rect 137704 244718 137756 244724
rect 138452 240945 138480 245495
rect 138438 240936 138494 240945
rect 138438 240871 138494 240880
rect 138912 238633 138940 248934
rect 139004 242849 139032 251790
rect 139740 248425 139768 255870
rect 139818 253312 139874 253321
rect 139818 253247 139874 253256
rect 139832 253146 139860 253247
rect 139820 253140 139872 253146
rect 139820 253082 139872 253088
rect 139726 248416 139782 248425
rect 139726 248351 139782 248360
rect 140096 244776 140148 244782
rect 140096 244718 140148 244724
rect 140108 244073 140136 244718
rect 140094 244064 140150 244073
rect 140094 243999 140150 244008
rect 138990 242840 139046 242849
rect 138990 242775 139046 242784
rect 138898 238624 138954 238633
rect 138898 238559 138954 238568
rect 140292 237273 140320 263418
rect 140370 261744 140426 261753
rect 140370 261679 140426 261688
rect 140384 261442 140412 261679
rect 140372 261436 140424 261442
rect 140372 261378 140424 261384
rect 140370 260384 140426 260393
rect 140370 260319 140426 260328
rect 140384 260082 140412 260319
rect 140372 260076 140424 260082
rect 140372 260018 140424 260024
rect 140554 258888 140610 258897
rect 140554 258823 140610 258832
rect 140568 258654 140596 258823
rect 140556 258648 140608 258654
rect 140556 258590 140608 258596
rect 140554 257528 140610 257537
rect 140554 257463 140610 257472
rect 140568 257362 140596 257463
rect 140556 257356 140608 257362
rect 140556 257298 140608 257304
rect 140648 257288 140700 257294
rect 140648 257230 140700 257236
rect 140462 256168 140518 256177
rect 140462 256103 140518 256112
rect 140476 250714 140504 256103
rect 140554 254672 140610 254681
rect 140554 254607 140610 254616
rect 140568 254506 140596 254607
rect 140556 254500 140608 254506
rect 140556 254442 140608 254448
rect 140554 251952 140610 251961
rect 140554 251887 140610 251896
rect 140568 251786 140596 251887
rect 140556 251780 140608 251786
rect 140556 251722 140608 251728
rect 140476 250686 140596 250714
rect 140372 246204 140424 246210
rect 140372 246146 140424 246152
rect 140384 245569 140412 246146
rect 140568 246142 140596 250686
rect 140660 249785 140688 257230
rect 140738 250592 140794 250601
rect 140738 250527 140794 250536
rect 140646 249776 140702 249785
rect 140646 249711 140702 249720
rect 140648 247292 140700 247298
rect 140648 247234 140700 247240
rect 140660 246793 140688 247234
rect 140646 246784 140702 246793
rect 140646 246719 140702 246728
rect 140556 246136 140608 246142
rect 140556 246078 140608 246084
rect 140370 245560 140426 245569
rect 140370 245495 140426 245504
rect 140752 245410 140780 250527
rect 140384 245382 140780 245410
rect 140278 237264 140334 237273
rect 140384 237234 140412 245382
rect 140554 240664 140610 240673
rect 140554 240599 140556 240608
rect 140608 240599 140610 240608
rect 140556 240570 140608 240576
rect 140554 239304 140610 239313
rect 140554 239239 140556 239248
rect 140608 239239 140610 239248
rect 140556 239210 140608 239216
rect 140278 237199 140334 237208
rect 140372 237228 140424 237234
rect 140372 237170 140424 237176
rect 148742 236040 148798 236049
rect 167970 236040 168026 236049
rect 148798 235998 149152 236026
rect 148742 235975 148798 235984
rect 147270 235904 147326 235913
rect 142408 235862 143388 235890
rect 144308 235862 144644 235890
rect 145228 235862 145288 235890
rect 138164 233760 138216 233766
rect 138164 233702 138216 233708
rect 137612 226144 137664 226150
rect 137612 226086 137664 226092
rect 137520 225600 137572 225606
rect 137520 225542 137572 225548
rect 137334 223256 137390 223265
rect 137334 223191 137390 223200
rect 137150 220128 137206 220137
rect 137150 220063 137206 220072
rect 137058 217000 137114 217009
rect 137058 216935 137114 216944
rect 136966 210744 137022 210753
rect 136966 210679 137022 210688
rect 136876 204792 136928 204798
rect 136874 204760 136876 204769
rect 136928 204760 136930 204769
rect 136874 204695 136930 204704
rect 137336 189628 137388 189634
rect 137336 189570 137388 189576
rect 137348 185729 137376 189570
rect 137334 185720 137390 185729
rect 137334 185655 137390 185664
rect 137150 143288 137206 143297
rect 137150 143223 137206 143232
rect 136874 141928 136930 141937
rect 136874 141863 136930 141872
rect 136888 141422 136916 141863
rect 136876 141416 136928 141422
rect 136876 141358 136928 141364
rect 136888 140146 136916 141358
rect 136888 140118 137008 140146
rect 136876 139036 136928 139042
rect 136876 138978 136928 138984
rect 136888 132961 136916 138978
rect 136874 132952 136930 132961
rect 136874 132887 136930 132896
rect 136876 132372 136928 132378
rect 136876 132314 136928 132320
rect 136888 120449 136916 132314
rect 136980 123305 137008 140118
rect 137164 137138 137192 143223
rect 137334 141112 137390 141121
rect 137334 141047 137390 141056
rect 137244 140668 137296 140674
rect 137244 140610 137296 140616
rect 137256 140305 137284 140610
rect 137348 140606 137376 141047
rect 137336 140600 137388 140606
rect 137336 140542 137388 140548
rect 137242 140296 137298 140305
rect 137242 140231 137298 140240
rect 137152 137132 137204 137138
rect 137152 137074 137204 137080
rect 137256 129833 137284 140231
rect 137348 132378 137376 140542
rect 137428 137132 137480 137138
rect 137428 137074 137480 137080
rect 137336 132372 137388 132378
rect 137336 132314 137388 132320
rect 137242 129824 137298 129833
rect 137242 129759 137298 129768
rect 137440 127550 137468 137074
rect 137060 127544 137112 127550
rect 137060 127486 137112 127492
rect 137428 127544 137480 127550
rect 137428 127486 137480 127492
rect 137072 126025 137100 127486
rect 137058 126016 137114 126025
rect 137058 125951 137114 125960
rect 136966 123296 137022 123305
rect 136966 123231 137022 123240
rect 136874 120440 136930 120449
rect 136874 120375 136930 120384
rect 136874 113232 136930 113241
rect 136874 113167 136930 113176
rect 136888 112998 136916 113167
rect 136876 112992 136928 112998
rect 136876 112934 136928 112940
rect 136876 110952 136928 110958
rect 136876 110894 136928 110900
rect 136888 110793 136916 110894
rect 136874 110784 136930 110793
rect 136874 110719 136930 110728
rect 137532 98553 137560 225542
rect 137612 225328 137664 225334
rect 137612 225270 137664 225276
rect 137624 191985 137652 225270
rect 137704 215876 137756 215882
rect 137704 215818 137756 215824
rect 137610 191976 137666 191985
rect 137610 191911 137666 191920
rect 137716 189634 137744 215818
rect 138176 208305 138204 233702
rect 138162 208296 138218 208305
rect 138162 208231 138218 208240
rect 137796 202072 137848 202078
rect 137796 202014 137848 202020
rect 137704 189628 137756 189634
rect 137704 189570 137756 189576
rect 137808 188698 137836 202014
rect 137624 188670 137836 188698
rect 137624 182601 137652 188670
rect 137794 188576 137850 188585
rect 137794 188511 137850 188520
rect 137808 188342 137836 188511
rect 142408 188342 142436 235862
rect 144616 233154 144644 235862
rect 145154 235360 145210 235369
rect 145154 235295 145156 235304
rect 145208 235295 145210 235304
rect 145156 235266 145208 235272
rect 144604 233148 144656 233154
rect 144604 233090 144656 233096
rect 145260 233086 145288 235862
rect 146226 235670 146254 235876
rect 146824 235862 147270 235890
rect 145340 235664 145392 235670
rect 145340 235606 145392 235612
rect 146214 235664 146266 235670
rect 146214 235606 146266 235612
rect 145248 233080 145300 233086
rect 145248 233022 145300 233028
rect 145154 216184 145210 216193
rect 145154 216119 145210 216128
rect 145168 215882 145196 216119
rect 145156 215876 145208 215882
rect 145156 215818 145208 215824
rect 145352 204798 145380 235606
rect 146824 233766 146852 235862
rect 148172 235862 148232 235890
rect 147270 235839 147326 235848
rect 148204 234961 148232 235862
rect 149124 235194 149152 235998
rect 167970 235975 168026 235984
rect 150104 235862 150440 235890
rect 150412 235262 150440 235862
rect 150688 235862 151024 235890
rect 150400 235256 150452 235262
rect 150400 235198 150452 235204
rect 149112 235188 149164 235194
rect 149112 235130 149164 235136
rect 148190 234952 148246 234961
rect 148190 234887 148246 234896
rect 146812 233760 146864 233766
rect 146812 233702 146864 233708
rect 149296 233760 149348 233766
rect 150688 233737 150716 235862
rect 152022 235641 152050 235876
rect 152620 235862 152956 235890
rect 153968 235862 154304 235890
rect 154888 235862 155224 235890
rect 155900 235862 156144 235890
rect 156820 235862 157156 235890
rect 157832 235862 158168 235890
rect 158752 235862 158904 235890
rect 159764 235862 160100 235890
rect 160684 235862 161020 235890
rect 161696 235862 162032 235890
rect 152008 235632 152064 235641
rect 152008 235567 152064 235576
rect 152620 235330 152648 235862
rect 152608 235324 152660 235330
rect 152608 235266 152660 235272
rect 149296 233702 149348 233708
rect 150674 233728 150730 233737
rect 149308 222820 149336 233702
rect 150674 233663 150730 233672
rect 150688 233222 150716 233663
rect 153344 233556 153396 233562
rect 153344 233498 153396 233504
rect 151964 233420 152016 233426
rect 151964 233362 152016 233368
rect 150676 233216 150728 233222
rect 150676 233158 150728 233164
rect 151044 233216 151096 233222
rect 151044 233158 151096 233164
rect 150584 232876 150636 232882
rect 150584 232818 150636 232824
rect 150596 222698 150624 232818
rect 151056 222820 151084 233158
rect 151976 222820 152004 233362
rect 150150 222670 150624 222698
rect 153356 222562 153384 233498
rect 153712 233284 153764 233290
rect 153712 233226 153764 233232
rect 153724 222820 153752 233226
rect 154276 232474 154304 235862
rect 154724 233692 154776 233698
rect 154724 233634 154776 233640
rect 154264 232468 154316 232474
rect 154264 232410 154316 232416
rect 154736 222698 154764 233634
rect 155196 232610 155224 235862
rect 155460 232944 155512 232950
rect 155460 232886 155512 232892
rect 155184 232604 155236 232610
rect 155184 232546 155236 232552
rect 155472 222820 155500 232886
rect 156116 232678 156144 235862
rect 156380 233012 156432 233018
rect 156380 232954 156432 232960
rect 156104 232672 156156 232678
rect 156104 232614 156156 232620
rect 156392 222820 156420 232954
rect 157128 232542 157156 235862
rect 158140 232678 158168 235862
rect 158876 232746 158904 235862
rect 158864 232740 158916 232746
rect 158864 232682 158916 232688
rect 158036 232672 158088 232678
rect 158036 232614 158088 232620
rect 158128 232672 158180 232678
rect 158128 232614 158180 232620
rect 157576 232604 157628 232610
rect 157576 232546 157628 232552
rect 157116 232536 157168 232542
rect 157116 232478 157168 232484
rect 156748 232468 156800 232474
rect 156748 232410 156800 232416
rect 154658 222670 154764 222698
rect 156760 222698 156788 232410
rect 157588 222698 157616 232546
rect 158048 225470 158076 232614
rect 160072 232542 160100 235862
rect 160336 232672 160388 232678
rect 160336 232614 160388 232620
rect 159140 232536 159192 232542
rect 159140 232478 159192 232484
rect 160060 232536 160112 232542
rect 160060 232478 160112 232484
rect 158036 225464 158088 225470
rect 158036 225406 158088 225412
rect 159048 225464 159100 225470
rect 159048 225406 159100 225412
rect 159060 222820 159088 225406
rect 159152 222698 159180 232478
rect 160348 222834 160376 232614
rect 160992 232474 161020 235862
rect 161808 232740 161860 232746
rect 161808 232682 161860 232688
rect 160980 232468 161032 232474
rect 160980 232410 161032 232416
rect 160348 222806 160822 222834
rect 161820 222698 161848 232682
rect 162004 225470 162032 235862
rect 162280 235862 162616 235890
rect 163292 235862 163628 235890
rect 164548 235862 164608 235890
rect 162280 233766 162308 235862
rect 162268 233760 162320 233766
rect 162268 233702 162320 233708
rect 163292 232882 163320 235862
rect 164580 233222 164608 235862
rect 165224 235862 165560 235890
rect 166144 235862 166480 235890
rect 167340 235862 167492 235890
rect 165224 233426 165252 235862
rect 166144 233562 166172 235862
rect 166132 233556 166184 233562
rect 166132 233498 166184 233504
rect 165212 233420 165264 233426
rect 165212 233362 165264 233368
rect 167340 233290 167368 235862
rect 167694 235768 167750 235777
rect 167694 235703 167750 235712
rect 167708 235262 167736 235703
rect 167696 235256 167748 235262
rect 167696 235198 167748 235204
rect 167984 235194 168012 235975
rect 168076 235862 168412 235890
rect 169088 235862 169424 235890
rect 170008 235862 170344 235890
rect 167972 235188 168024 235194
rect 167972 235130 168024 235136
rect 168076 233698 168104 235862
rect 168064 233692 168116 233698
rect 168064 233634 168116 233640
rect 167328 233284 167380 233290
rect 167328 233226 167380 233232
rect 164568 233216 164620 233222
rect 164568 233158 164620 233164
rect 165120 233148 165172 233154
rect 165120 233090 165172 233096
rect 163280 232876 163332 232882
rect 163280 232818 163332 232824
rect 162268 232536 162320 232542
rect 162268 232478 162320 232484
rect 161992 225464 162044 225470
rect 161992 225406 162044 225412
rect 162280 222834 162308 232478
rect 163188 232468 163240 232474
rect 163188 232410 163240 232416
rect 163200 222834 163228 232410
rect 164382 226656 164438 226665
rect 164382 226591 164438 226600
rect 164396 226257 164424 226591
rect 164382 226248 164438 226257
rect 164382 226183 164438 226192
rect 164384 225464 164436 225470
rect 164384 225406 164436 225412
rect 162280 222806 162662 222834
rect 163200 222806 163490 222834
rect 164396 222820 164424 225406
rect 156760 222670 157326 222698
rect 157588 222670 158154 222698
rect 159152 222670 159994 222698
rect 161742 222670 161848 222698
rect 152818 222534 153384 222562
rect 165132 219282 165160 233090
rect 169088 232950 169116 235862
rect 170008 233018 170036 235862
rect 169996 233012 170048 233018
rect 169996 232954 170048 232960
rect 169076 232944 169128 232950
rect 169076 232886 169128 232892
rect 165120 219276 165172 219282
rect 165120 219218 165172 219224
rect 145340 204792 145392 204798
rect 145340 204734 145392 204740
rect 145154 202856 145210 202865
rect 145154 202791 145210 202800
rect 145168 202078 145196 202791
rect 145156 202072 145208 202078
rect 145156 202014 145208 202020
rect 145614 189528 145670 189537
rect 145614 189463 145670 189472
rect 137796 188336 137848 188342
rect 137796 188278 137848 188284
rect 142396 188336 142448 188342
rect 142396 188278 142448 188284
rect 143040 188336 143092 188342
rect 143040 188278 143092 188284
rect 138900 188268 138952 188274
rect 138900 188210 138952 188216
rect 137610 182592 137666 182601
rect 137610 182527 137666 182536
rect 138912 179473 138940 188210
rect 138898 179464 138954 179473
rect 138898 179399 138954 179408
rect 143052 172702 143080 188278
rect 145628 188274 145656 189463
rect 145616 188268 145668 188274
rect 145616 188210 145668 188216
rect 149216 181202 149244 182836
rect 149204 181196 149256 181202
rect 149204 181138 149256 181144
rect 149768 181134 149796 182836
rect 150320 182822 150426 182850
rect 149756 181128 149808 181134
rect 149756 181070 149808 181076
rect 149204 180924 149256 180930
rect 149204 180866 149256 180872
rect 147824 180856 147876 180862
rect 147824 180798 147876 180804
rect 145064 180788 145116 180794
rect 145064 180730 145116 180736
rect 143684 180584 143736 180590
rect 143684 180526 143736 180532
rect 143040 172696 143092 172702
rect 143040 172638 143092 172644
rect 143696 169794 143724 180526
rect 145076 169794 145104 180730
rect 146444 180652 146496 180658
rect 146444 180594 146496 180600
rect 146456 169794 146484 180594
rect 147836 169794 147864 180798
rect 149216 169794 149244 180866
rect 150320 172838 150348 182822
rect 151056 181338 151084 182836
rect 151622 182822 151728 182850
rect 151044 181332 151096 181338
rect 151044 181274 151096 181280
rect 150584 181060 150636 181066
rect 150584 181002 150636 181008
rect 150308 172832 150360 172838
rect 150308 172774 150360 172780
rect 150596 169794 150624 181002
rect 151700 172566 151728 182822
rect 152252 181338 152280 182836
rect 152910 182822 153384 182850
rect 151872 181332 151924 181338
rect 151872 181274 151924 181280
rect 152240 181332 152292 181338
rect 152240 181274 152292 181280
rect 153252 181332 153304 181338
rect 153252 181274 153304 181280
rect 151884 172770 151912 181274
rect 151964 180992 152016 180998
rect 151964 180934 152016 180940
rect 151872 172764 151924 172770
rect 151872 172706 151924 172712
rect 151688 172560 151740 172566
rect 151688 172502 151740 172508
rect 151976 169794 152004 180934
rect 153160 173036 153212 173042
rect 153160 172978 153212 172984
rect 153172 172430 153200 172978
rect 153264 172634 153292 181274
rect 153356 173042 153384 182822
rect 153448 181338 153476 182836
rect 154106 182822 154672 182850
rect 153436 181332 153488 181338
rect 153436 181274 153488 181280
rect 153344 173036 153396 173042
rect 153344 172978 153396 172984
rect 154540 172968 154592 172974
rect 154540 172910 154592 172916
rect 153344 172900 153396 172906
rect 153344 172842 153396 172848
rect 153252 172628 153304 172634
rect 153252 172570 153304 172576
rect 153160 172424 153212 172430
rect 153160 172366 153212 172372
rect 153356 169794 153384 172842
rect 143572 169766 143724 169794
rect 144952 169766 145104 169794
rect 146332 169766 146484 169794
rect 147712 169766 147864 169794
rect 149092 169766 149244 169794
rect 150564 169766 150624 169794
rect 151944 169766 152004 169794
rect 153324 169766 153384 169794
rect 154552 169794 154580 172910
rect 154644 172362 154672 182822
rect 154736 182057 154764 182836
rect 154722 182048 154778 182057
rect 154722 181983 154778 181992
rect 154724 181332 154776 181338
rect 154724 181274 154776 181280
rect 154736 172498 154764 181274
rect 155288 181241 155316 182836
rect 155274 181232 155330 181241
rect 155274 181167 155330 181176
rect 155932 180561 155960 182836
rect 156576 180561 156604 182836
rect 157220 180833 157248 182836
rect 157206 180824 157262 180833
rect 157206 180759 157262 180768
rect 157772 180697 157800 182836
rect 158220 181196 158272 181202
rect 158220 181138 158272 181144
rect 157758 180688 157814 180697
rect 157758 180623 157814 180632
rect 155918 180552 155974 180561
rect 155918 180487 155974 180496
rect 156562 180552 156618 180561
rect 156562 180487 156618 180496
rect 158232 173042 158260 181138
rect 158416 180969 158444 182836
rect 159060 181105 159088 182836
rect 159046 181096 159102 181105
rect 159046 181031 159102 181040
rect 158402 180960 158458 180969
rect 158402 180895 158458 180904
rect 159612 180590 159640 182836
rect 160256 180794 160284 182836
rect 160336 181128 160388 181134
rect 160336 181070 160388 181076
rect 160244 180788 160296 180794
rect 160244 180730 160296 180736
rect 159600 180584 159652 180590
rect 159600 180526 159652 180532
rect 158220 173036 158272 173042
rect 158220 172978 158272 172984
rect 158956 173036 159008 173042
rect 158956 172978 159008 172984
rect 155736 172696 155788 172702
rect 155736 172638 155788 172644
rect 157852 172696 157904 172702
rect 157852 172638 157904 172644
rect 154724 172492 154776 172498
rect 154724 172434 154776 172440
rect 154632 172356 154684 172362
rect 154632 172298 154684 172304
rect 155748 169794 155776 172638
rect 157864 169794 157892 172638
rect 158968 169794 158996 172978
rect 160348 169794 160376 181070
rect 160900 180658 160928 182836
rect 161452 180862 161480 182836
rect 162096 180930 162124 182836
rect 162740 181066 162768 182836
rect 162728 181060 162780 181066
rect 162728 181002 162780 181008
rect 163292 180998 163320 182836
rect 163280 180992 163332 180998
rect 163280 180934 163332 180940
rect 162084 180924 162136 180930
rect 162084 180866 162136 180872
rect 161440 180856 161492 180862
rect 161440 180798 161492 180804
rect 160888 180652 160940 180658
rect 160888 180594 160940 180600
rect 163936 172906 163964 182836
rect 164594 182822 164700 182850
rect 164672 172974 164700 182822
rect 164660 172968 164712 172974
rect 164660 172910 164712 172916
rect 163924 172900 163976 172906
rect 163924 172842 163976 172848
rect 161716 172832 161768 172838
rect 161716 172774 161768 172780
rect 161728 169794 161756 172774
rect 163096 172764 163148 172770
rect 163096 172706 163148 172712
rect 163108 169794 163136 172706
rect 165132 172702 165160 219218
rect 167878 212784 167934 212793
rect 167878 212719 167934 212728
rect 167892 203370 167920 212719
rect 167880 203364 167932 203370
rect 167880 203306 167932 203312
rect 167970 192792 168026 192801
rect 167970 192727 168026 192736
rect 167984 192626 168012 192727
rect 167972 192620 168024 192626
rect 167972 192562 168024 192568
rect 170652 175762 170680 268926
rect 173490 263104 173546 263113
rect 173490 263039 173546 263048
rect 173398 261744 173454 261753
rect 173398 261679 173454 261688
rect 173124 257288 173176 257294
rect 173124 257230 173176 257236
rect 173136 254386 173164 257230
rect 173306 256168 173362 256177
rect 173306 256103 173362 256112
rect 173320 255934 173348 256103
rect 173308 255928 173360 255934
rect 173308 255870 173360 255876
rect 173306 254672 173362 254681
rect 173306 254607 173362 254616
rect 173320 254506 173348 254607
rect 173308 254500 173360 254506
rect 173308 254442 173360 254448
rect 173136 254358 173348 254386
rect 173320 249105 173348 254358
rect 173306 249096 173362 249105
rect 173306 249031 173362 249040
rect 173412 248930 173440 261679
rect 173504 250290 173532 263039
rect 173766 260384 173822 260393
rect 173766 260319 173822 260328
rect 173674 257528 173730 257537
rect 173674 257463 173730 257472
rect 173584 255588 173636 255594
rect 173584 255530 173636 255536
rect 173596 250601 173624 255530
rect 173582 250592 173638 250601
rect 173582 250527 173638 250536
rect 173584 250352 173636 250358
rect 173584 250294 173636 250300
rect 173492 250284 173544 250290
rect 173492 250226 173544 250232
rect 173400 248924 173452 248930
rect 173400 248866 173452 248872
rect 173492 248720 173544 248726
rect 173492 248662 173544 248668
rect 173504 247745 173532 248662
rect 173490 247736 173546 247745
rect 173490 247671 173546 247680
rect 173308 246544 173360 246550
rect 173308 246486 173360 246492
rect 173320 246385 173348 246486
rect 173306 246376 173362 246385
rect 173306 246311 173362 246320
rect 172756 246204 172808 246210
rect 172756 246146 172808 246152
rect 172768 244889 172796 246146
rect 172754 244880 172810 244889
rect 172754 244815 172810 244824
rect 173124 244028 173176 244034
rect 173124 243970 173176 243976
rect 173136 243529 173164 243970
rect 173122 243520 173178 243529
rect 173122 243455 173178 243464
rect 173596 240786 173624 250294
rect 173688 246074 173716 257463
rect 173780 248862 173808 260319
rect 189328 260082 189356 268994
rect 189420 268990 189448 269470
rect 196688 268990 196716 269538
rect 203772 269058 203800 271916
rect 203760 269052 203812 269058
rect 203760 268994 203812 269000
rect 189408 268984 189460 268990
rect 189408 268926 189460 268932
rect 196676 268984 196728 268990
rect 196676 268926 196728 268932
rect 210948 268922 210976 271916
rect 210016 268916 210068 268922
rect 210016 268858 210068 268864
rect 210936 268916 210988 268922
rect 210936 268858 210988 268864
rect 210028 268394 210056 268858
rect 218032 268417 218060 271916
rect 209936 268366 210056 268394
rect 218018 268408 218074 268417
rect 209936 261306 209964 268366
rect 218018 268343 218074 268352
rect 203852 261300 203904 261306
rect 203852 261242 203904 261248
rect 209924 261300 209976 261306
rect 209924 261242 209976 261248
rect 189316 260076 189368 260082
rect 189316 260018 189368 260024
rect 190512 260076 190564 260082
rect 190512 260018 190564 260024
rect 173858 258888 173914 258897
rect 173858 258823 173914 258832
rect 173768 248856 173820 248862
rect 173768 248798 173820 248804
rect 173872 247570 173900 258823
rect 190524 257772 190552 260018
rect 203864 257772 203892 261242
rect 225208 260694 225236 271916
rect 225840 262932 225892 262938
rect 225840 262874 225892 262880
rect 225748 261436 225800 261442
rect 225748 261378 225800 261384
rect 217192 260688 217244 260694
rect 217192 260630 217244 260636
rect 225196 260688 225248 260694
rect 225196 260630 225248 260636
rect 217204 257772 217232 260630
rect 181034 257392 181090 257401
rect 181034 257327 181090 257336
rect 181048 257294 181076 257327
rect 181036 257288 181088 257294
rect 181036 257230 181088 257236
rect 181034 256440 181090 256449
rect 181034 256375 181090 256384
rect 181048 255934 181076 256375
rect 176160 255928 176212 255934
rect 176160 255870 176212 255876
rect 178276 255928 178328 255934
rect 178276 255870 178328 255876
rect 181036 255928 181088 255934
rect 181036 255870 181088 255876
rect 173950 253312 174006 253321
rect 173950 253247 174006 253256
rect 173860 247564 173912 247570
rect 173860 247506 173912 247512
rect 173676 246068 173728 246074
rect 173676 246010 173728 246016
rect 173964 243422 173992 253247
rect 174042 251952 174098 251961
rect 174042 251887 174044 251896
rect 174096 251887 174098 251896
rect 174044 251858 174096 251864
rect 174044 251780 174096 251786
rect 174044 251722 174096 251728
rect 173952 243416 174004 243422
rect 173952 243358 174004 243364
rect 174056 242169 174084 251722
rect 176172 246142 176200 255870
rect 176344 254568 176396 254574
rect 176344 254510 176396 254516
rect 176252 254500 176304 254506
rect 176252 254442 176304 254448
rect 176160 246136 176212 246142
rect 176160 246078 176212 246084
rect 176264 244782 176292 254442
rect 176356 246210 176384 254510
rect 178288 248726 178316 255870
rect 181586 255624 181642 255633
rect 181586 255559 181642 255568
rect 222712 255588 222764 255594
rect 181034 254672 181090 254681
rect 181034 254607 181090 254616
rect 181048 254574 181076 254607
rect 181036 254568 181088 254574
rect 181036 254510 181088 254516
rect 181600 254506 181628 255559
rect 222712 255530 222764 255536
rect 179196 254500 179248 254506
rect 179196 254442 179248 254448
rect 181588 254500 181640 254506
rect 181588 254442 181640 254448
rect 179012 253480 179064 253486
rect 179012 253422 179064 253428
rect 178920 251916 178972 251922
rect 178920 251858 178972 251864
rect 178276 248720 178328 248726
rect 178276 248662 178328 248668
rect 176344 246204 176396 246210
rect 176344 246146 176396 246152
rect 176252 244776 176304 244782
rect 176252 244718 176304 244724
rect 178932 243014 178960 251858
rect 179024 244034 179052 253422
rect 179208 246550 179236 254442
rect 181034 253856 181090 253865
rect 181034 253791 181090 253800
rect 181048 253486 181076 253791
rect 181036 253480 181088 253486
rect 181036 253422 181088 253428
rect 222724 253026 222752 255530
rect 225760 255066 225788 261378
rect 225852 255186 225880 262874
rect 226208 260076 226260 260082
rect 226208 260018 226260 260024
rect 226116 257288 226168 257294
rect 226116 257230 226168 257236
rect 225930 255624 225986 255633
rect 225930 255559 225986 255568
rect 225944 255186 225972 255559
rect 225840 255180 225892 255186
rect 225840 255122 225892 255128
rect 225932 255180 225984 255186
rect 225932 255122 225984 255128
rect 225760 255038 225972 255066
rect 225840 254976 225892 254982
rect 225840 254918 225892 254924
rect 225746 253856 225802 253865
rect 225746 253791 225802 253800
rect 225760 253418 225788 253791
rect 225748 253412 225800 253418
rect 225748 253354 225800 253360
rect 222632 252998 222752 253026
rect 181586 252904 181642 252913
rect 181586 252839 181642 252848
rect 181600 251786 181628 252839
rect 181678 252088 181734 252097
rect 181678 252023 181734 252032
rect 181588 251780 181640 251786
rect 181588 251722 181640 251728
rect 181496 250284 181548 250290
rect 181496 250226 181548 250232
rect 181508 249785 181536 250226
rect 181494 249776 181550 249785
rect 181494 249711 181550 249720
rect 179196 246544 179248 246550
rect 179196 246486 179248 246492
rect 181588 246136 181640 246142
rect 181588 246078 181640 246084
rect 181600 245433 181628 246078
rect 181586 245424 181642 245433
rect 181586 245359 181642 245368
rect 179012 244028 179064 244034
rect 179012 243970 179064 243976
rect 181692 243506 181720 252023
rect 182322 251136 182378 251145
rect 182322 251071 182378 251080
rect 222632 251122 222660 252998
rect 222632 251094 222844 251122
rect 182336 250358 182364 251071
rect 182324 250352 182376 250358
rect 181770 250320 181826 250329
rect 182324 250294 182376 250300
rect 181770 250255 181826 250264
rect 181600 243478 181720 243506
rect 181784 243506 181812 250255
rect 181956 248924 182008 248930
rect 181956 248866 182008 248872
rect 181864 248856 181916 248862
rect 181864 248798 181916 248804
rect 181876 248289 181904 248798
rect 181968 248697 181996 248866
rect 181954 248688 182010 248697
rect 181954 248623 182010 248632
rect 181862 248280 181918 248289
rect 181862 248215 181918 248224
rect 182324 247564 182376 247570
rect 182324 247506 182376 247512
rect 182336 247201 182364 247506
rect 182322 247192 182378 247201
rect 182322 247127 182378 247136
rect 182324 246204 182376 246210
rect 182324 246146 182376 246152
rect 182336 245841 182364 246146
rect 182322 245832 182378 245841
rect 182322 245767 182378 245776
rect 182324 244776 182376 244782
rect 182324 244718 182376 244724
rect 182336 244617 182364 244718
rect 182322 244608 182378 244617
rect 182322 244543 182378 244552
rect 222632 243506 222660 251094
rect 222816 251038 222844 251094
rect 222804 251032 222856 251038
rect 222804 250974 222856 250980
rect 225852 250442 225880 254918
rect 225760 250414 225880 250442
rect 225760 249377 225788 250414
rect 225838 250320 225894 250329
rect 225838 250255 225894 250264
rect 225746 249368 225802 249377
rect 225746 249303 225802 249312
rect 225852 248998 225880 250255
rect 225840 248992 225892 248998
rect 225840 248934 225892 248940
rect 225944 248425 225972 255038
rect 226022 251136 226078 251145
rect 226022 251071 226078 251080
rect 225930 248416 225986 248425
rect 225930 248351 225986 248360
rect 225564 245252 225616 245258
rect 225564 245194 225616 245200
rect 225576 244889 225604 245194
rect 225562 244880 225618 244889
rect 225562 244815 225618 244824
rect 225564 244776 225616 244782
rect 225564 244718 225616 244724
rect 225576 244073 225604 244718
rect 225562 244064 225618 244073
rect 225562 243999 225618 244008
rect 181784 243478 181996 243506
rect 181036 243416 181088 243422
rect 181034 243384 181036 243393
rect 181088 243384 181090 243393
rect 181034 243319 181090 243328
rect 178920 243008 178972 243014
rect 178920 242950 178972 242956
rect 181220 243008 181272 243014
rect 181220 242950 181272 242956
rect 181232 242849 181260 242950
rect 181218 242840 181274 242849
rect 181218 242775 181274 242784
rect 174042 242160 174098 242169
rect 174042 242095 174098 242104
rect 173320 240758 173624 240786
rect 173320 239313 173348 240758
rect 173582 240664 173638 240673
rect 181600 240634 181628 243478
rect 173582 240599 173584 240608
rect 173636 240599 173638 240608
rect 181588 240628 181640 240634
rect 173584 240570 173636 240576
rect 181588 240570 181640 240576
rect 173306 239304 173362 239313
rect 181968 239274 181996 243478
rect 222448 243478 222660 243506
rect 222002 241982 222200 242010
rect 185648 239342 185676 241860
rect 189236 239721 189264 241860
rect 189222 239712 189278 239721
rect 189222 239647 189278 239656
rect 192916 239449 192944 241860
rect 196504 240401 196532 241860
rect 196490 240392 196546 240401
rect 196490 240327 196546 240336
rect 192902 239440 192958 239449
rect 192902 239375 192958 239384
rect 185636 239336 185688 239342
rect 185636 239278 185688 239284
rect 186464 239336 186516 239342
rect 186464 239278 186516 239284
rect 173306 239239 173362 239248
rect 173400 239268 173452 239274
rect 173400 239210 173452 239216
rect 181956 239268 182008 239274
rect 181956 239210 182008 239216
rect 173412 237953 173440 239210
rect 173398 237944 173454 237953
rect 173398 237879 173454 237888
rect 172940 237228 172992 237234
rect 172940 237170 172992 237176
rect 172952 236593 172980 237170
rect 172938 236584 172994 236593
rect 172938 236519 172994 236528
rect 185084 230292 185136 230298
rect 185084 230234 185136 230240
rect 185096 227716 185124 230234
rect 186476 227578 186504 239278
rect 200184 238594 200212 241860
rect 203772 241738 203800 241860
rect 207452 241738 207480 241860
rect 211040 241738 211068 241860
rect 214720 241738 214748 241860
rect 203128 241710 203800 241738
rect 207268 241710 207480 241738
rect 210028 241710 211068 241738
rect 214168 241710 214748 241738
rect 200172 238588 200224 238594
rect 200172 238530 200224 238536
rect 200184 238497 200212 238530
rect 200170 238488 200226 238497
rect 200170 238423 200226 238432
rect 203128 236321 203156 241710
rect 203114 236312 203170 236321
rect 203114 236247 203170 236256
rect 203128 235874 203156 236247
rect 203116 235868 203168 235874
rect 203116 235810 203168 235816
rect 207268 234417 207296 241710
rect 210028 234553 210056 241710
rect 210014 234544 210070 234553
rect 210014 234479 210070 234488
rect 207254 234408 207310 234417
rect 207254 234343 207310 234352
rect 210016 230428 210068 230434
rect 210016 230370 210068 230376
rect 197504 230360 197556 230366
rect 197504 230302 197556 230308
rect 197516 227716 197544 230302
rect 210028 227716 210056 230370
rect 214168 230298 214196 241710
rect 218308 230366 218336 241860
rect 222172 237846 222200 241982
rect 222448 240673 222476 243478
rect 225748 242940 225800 242946
rect 225748 242882 225800 242888
rect 225760 242305 225788 242882
rect 225746 242296 225802 242305
rect 225746 242231 225802 242240
rect 222434 240664 222490 240673
rect 222434 240599 222490 240608
rect 222802 240664 222858 240673
rect 222802 240599 222858 240608
rect 221056 237840 221108 237846
rect 219766 237808 219822 237817
rect 221056 237782 221108 237788
rect 222160 237840 222212 237846
rect 222160 237782 222212 237788
rect 219766 237743 219822 237752
rect 219780 237234 219808 237743
rect 219768 237228 219820 237234
rect 219768 237170 219820 237176
rect 221068 230434 221096 237782
rect 222816 231046 222844 240599
rect 226036 239274 226064 251071
rect 226128 245841 226156 257230
rect 226220 247609 226248 260018
rect 226300 258648 226352 258654
rect 226300 258590 226352 258596
rect 226206 247600 226262 247609
rect 226206 247535 226262 247544
rect 226312 246657 226340 258590
rect 226482 257392 226538 257401
rect 226482 257327 226484 257336
rect 226536 257327 226538 257336
rect 226484 257298 226536 257304
rect 226482 256440 226538 256449
rect 226538 256398 226616 256426
rect 226482 256375 226538 256384
rect 226390 254672 226446 254681
rect 226390 254607 226446 254616
rect 226298 246648 226354 246657
rect 226298 246583 226354 246592
rect 226404 246210 226432 254607
rect 226482 252904 226538 252913
rect 226482 252839 226538 252848
rect 226392 246204 226444 246210
rect 226392 246146 226444 246152
rect 226114 245832 226170 245841
rect 226114 245767 226170 245776
rect 226496 243286 226524 252839
rect 226588 248930 226616 256398
rect 227218 252088 227274 252097
rect 227218 252023 227274 252032
rect 226576 248924 226628 248930
rect 226576 248866 226628 248872
rect 226484 243280 226536 243286
rect 226484 243222 226536 243228
rect 226484 243144 226536 243150
rect 226482 243112 226484 243121
rect 226536 243112 226538 243121
rect 226482 243047 226538 243056
rect 227232 240634 227260 252023
rect 227220 240628 227272 240634
rect 227220 240570 227272 240576
rect 226024 239268 226076 239274
rect 226024 239210 226076 239216
rect 222620 231040 222672 231046
rect 222620 230982 222672 230988
rect 222804 231040 222856 231046
rect 222804 230982 222856 230988
rect 221056 230428 221108 230434
rect 221056 230370 221108 230376
rect 218296 230360 218348 230366
rect 218296 230302 218348 230308
rect 214156 230292 214208 230298
rect 214156 230234 214208 230240
rect 222632 227646 222660 230982
rect 222436 227640 222488 227646
rect 222620 227640 222672 227646
rect 222488 227588 222554 227594
rect 222436 227582 222554 227588
rect 222620 227582 222672 227588
rect 186464 227572 186516 227578
rect 222448 227566 222554 227582
rect 186464 227514 186516 227520
rect 172020 225668 172072 225674
rect 172020 225610 172072 225616
rect 170640 175756 170692 175762
rect 170640 175698 170692 175704
rect 165120 172696 165172 172702
rect 165120 172638 165172 172644
rect 165856 172628 165908 172634
rect 165856 172570 165908 172576
rect 164476 172560 164528 172566
rect 164476 172502 164528 172508
rect 164488 169930 164516 172502
rect 165868 169930 165896 172570
rect 168616 172492 168668 172498
rect 168616 172434 168668 172440
rect 167236 172424 167288 172430
rect 167236 172366 167288 172372
rect 167248 169930 167276 172366
rect 168628 169930 168656 172434
rect 169996 172356 170048 172362
rect 169996 172298 170048 172304
rect 170008 169930 170036 172298
rect 164488 169902 164562 169930
rect 165868 169902 165942 169930
rect 167248 169902 167322 169930
rect 168628 169902 168702 169930
rect 170008 169902 170082 169930
rect 154552 169766 154704 169794
rect 155748 169766 156084 169794
rect 157556 169766 157892 169794
rect 158936 169766 158996 169794
rect 160316 169766 160376 169794
rect 161696 169766 161756 169794
rect 163076 169766 163136 169794
rect 164534 169780 164562 169902
rect 165914 169780 165942 169902
rect 167294 169780 167322 169902
rect 168674 169780 168702 169902
rect 170054 169780 170082 169902
rect 140280 169568 140332 169574
rect 140280 169510 140332 169516
rect 139634 164912 139690 164921
rect 139634 164847 139690 164856
rect 139648 164814 139676 164847
rect 139636 164808 139688 164814
rect 139636 164750 139688 164756
rect 139634 163552 139690 163561
rect 139634 163487 139636 163496
rect 139688 163487 139690 163496
rect 139636 163458 139688 163464
rect 139634 162192 139690 162201
rect 138164 162156 138216 162162
rect 139634 162127 139690 162136
rect 138164 162098 138216 162104
rect 137612 159300 137664 159306
rect 137612 159242 137664 159248
rect 137624 149514 137652 159242
rect 138176 155090 138204 162098
rect 139648 162094 139676 162127
rect 139636 162088 139688 162094
rect 139636 162030 139688 162036
rect 139634 160696 139690 160705
rect 139634 160631 139636 160640
rect 139688 160631 139690 160640
rect 139636 160602 139688 160608
rect 139634 159336 139690 159345
rect 139634 159271 139636 159280
rect 139688 159271 139690 159280
rect 139636 159242 139688 159248
rect 138900 158008 138952 158014
rect 138900 157950 138952 157956
rect 139634 157976 139690 157985
rect 138164 155084 138216 155090
rect 138164 155026 138216 155032
rect 137612 149508 137664 149514
rect 137612 149450 137664 149456
rect 138912 148193 138940 157950
rect 139634 157911 139636 157920
rect 139688 157911 139690 157920
rect 139636 157882 139688 157888
rect 139728 155084 139780 155090
rect 139728 155026 139780 155032
rect 139740 153769 139768 155026
rect 139726 153760 139782 153769
rect 139636 153724 139688 153730
rect 139726 153695 139782 153704
rect 139636 153666 139688 153672
rect 139648 152409 139676 153666
rect 139634 152400 139690 152409
rect 139634 152335 139690 152344
rect 139636 149576 139688 149582
rect 139634 149544 139636 149553
rect 139688 149544 139690 149553
rect 139634 149479 139690 149488
rect 138898 148184 138954 148193
rect 138898 148119 138954 148128
rect 140292 142617 140320 169510
rect 140554 169128 140610 169137
rect 140554 169063 140610 169072
rect 140568 168962 140596 169063
rect 140556 168956 140608 168962
rect 140556 168898 140608 168904
rect 140554 167768 140610 167777
rect 140554 167703 140610 167712
rect 140568 167602 140596 167703
rect 140556 167596 140608 167602
rect 140556 167538 140608 167544
rect 140554 166408 140610 166417
rect 140554 166343 140610 166352
rect 140568 166242 140596 166343
rect 140556 166236 140608 166242
rect 140556 166178 140608 166184
rect 140556 163448 140608 163454
rect 140556 163390 140608 163396
rect 140464 160728 140516 160734
rect 140464 160670 140516 160676
rect 140370 156616 140426 156625
rect 140370 156551 140426 156560
rect 140278 142608 140334 142617
rect 140278 142543 140334 142552
rect 140384 142034 140412 156551
rect 140476 150913 140504 160670
rect 140568 155129 140596 163390
rect 140554 155120 140610 155129
rect 140554 155055 140610 155064
rect 140462 150904 140518 150913
rect 140462 150839 140518 150848
rect 140556 146788 140608 146794
rect 140556 146730 140608 146736
rect 140568 146697 140596 146730
rect 140554 146688 140610 146697
rect 140554 146623 140610 146632
rect 140556 145428 140608 145434
rect 140556 145370 140608 145376
rect 140568 145337 140596 145370
rect 140554 145328 140610 145337
rect 140554 145263 140610 145272
rect 140556 144068 140608 144074
rect 140556 144010 140608 144016
rect 140568 143977 140596 144010
rect 140554 143968 140610 143977
rect 140554 143903 140610 143912
rect 167972 142232 168024 142238
rect 147914 142200 147970 142209
rect 147914 142135 147970 142144
rect 150674 142200 150730 142209
rect 167970 142200 167972 142209
rect 168524 142232 168576 142238
rect 168024 142200 168026 142209
rect 150730 142158 151024 142186
rect 150674 142135 150730 142144
rect 168524 142174 168576 142180
rect 167970 142135 168026 142144
rect 146810 142064 146866 142073
rect 140372 142028 140424 142034
rect 146866 142022 147496 142050
rect 146810 141999 146866 142008
rect 140372 141970 140424 141976
rect 142408 141886 143388 141914
rect 144308 141886 144644 141914
rect 145228 141886 145288 141914
rect 137612 122036 137664 122042
rect 137612 121978 137664 121984
rect 137518 98544 137574 98553
rect 137518 98479 137574 98488
rect 137624 92297 137652 121978
rect 137704 108232 137756 108238
rect 137704 108174 137756 108180
rect 137610 92288 137666 92297
rect 137610 92223 137666 92232
rect 137716 88761 137744 108174
rect 138162 94600 138218 94609
rect 138162 94535 138218 94544
rect 138176 94434 138204 94535
rect 142408 94434 142436 141886
rect 144616 139246 144644 141886
rect 144604 139240 144656 139246
rect 144604 139182 144656 139188
rect 145260 138770 145288 141886
rect 145352 141886 146240 141914
rect 145248 138764 145300 138770
rect 145248 138706 145300 138712
rect 144234 122344 144290 122353
rect 144234 122279 144290 122288
rect 144248 122042 144276 122279
rect 144236 122036 144288 122042
rect 144236 121978 144288 121984
rect 145352 110958 145380 141886
rect 147468 141354 147496 142022
rect 147928 141914 147956 142135
rect 147928 141886 148232 141914
rect 149092 141886 149152 141914
rect 150104 141886 150440 141914
rect 152036 141886 152096 141914
rect 147456 141348 147508 141354
rect 147456 141290 147508 141296
rect 147468 139897 147496 141290
rect 148204 139897 148232 141886
rect 149124 141121 149152 141886
rect 150412 141422 150440 141886
rect 150400 141416 150452 141422
rect 150400 141358 150452 141364
rect 149110 141112 149166 141121
rect 149110 141047 149166 141056
rect 152068 140441 152096 141886
rect 152712 141886 152956 141914
rect 153968 141886 154304 141914
rect 154888 141886 155224 141914
rect 155900 141886 156144 141914
rect 156820 141886 157156 141914
rect 157832 141886 158168 141914
rect 158752 141886 158904 141914
rect 159764 141886 160100 141914
rect 160684 141886 160928 141914
rect 161696 141886 162032 141914
rect 152054 140432 152110 140441
rect 152054 140367 152110 140376
rect 152712 139897 152740 141886
rect 147454 139888 147510 139897
rect 147454 139823 147510 139832
rect 148190 139888 148246 139897
rect 152698 139888 152754 139897
rect 148190 139823 148246 139832
rect 150584 139852 150636 139858
rect 152698 139823 152754 139832
rect 150584 139794 150636 139800
rect 150492 139376 150544 139382
rect 150492 139318 150544 139324
rect 149296 130332 149348 130338
rect 149296 130274 149348 130280
rect 149308 128708 149336 130274
rect 150504 128722 150532 139318
rect 150596 130338 150624 139794
rect 151780 139716 151832 139722
rect 151780 139658 151832 139664
rect 151792 130338 151820 139658
rect 151872 139444 151924 139450
rect 151872 139386 151924 139392
rect 150584 130332 150636 130338
rect 150584 130274 150636 130280
rect 151044 130332 151096 130338
rect 151044 130274 151096 130280
rect 151780 130332 151832 130338
rect 151780 130274 151832 130280
rect 150150 128694 150532 128722
rect 151056 128708 151084 130274
rect 151884 128722 151912 139386
rect 152712 139178 152740 139823
rect 154276 139586 154304 141886
rect 154264 139580 154316 139586
rect 154264 139522 154316 139528
rect 154724 139512 154776 139518
rect 154724 139454 154776 139460
rect 154632 139308 154684 139314
rect 154632 139250 154684 139256
rect 152700 139172 152752 139178
rect 152700 139114 152752 139120
rect 153344 139172 153396 139178
rect 153344 139114 153396 139120
rect 153356 130082 153384 139114
rect 153712 130332 153764 130338
rect 153712 130274 153764 130280
rect 153172 130054 153384 130082
rect 153172 128722 153200 130054
rect 151884 128694 151990 128722
rect 152818 128694 153200 128722
rect 153724 128708 153752 130274
rect 154644 128708 154672 139250
rect 154736 130338 154764 139454
rect 155196 138634 155224 141886
rect 156116 139790 156144 141886
rect 156104 139784 156156 139790
rect 156104 139726 156156 139732
rect 156104 139648 156156 139654
rect 156104 139590 156156 139596
rect 155184 138628 155236 138634
rect 155184 138570 155236 138576
rect 156116 131630 156144 139590
rect 157128 138906 157156 141886
rect 157576 139784 157628 139790
rect 157576 139726 157628 139732
rect 157484 139716 157536 139722
rect 157484 139658 157536 139664
rect 157300 139580 157352 139586
rect 157300 139522 157352 139528
rect 157116 138900 157168 138906
rect 157116 138842 157168 138848
rect 155460 131624 155512 131630
rect 155460 131566 155512 131572
rect 156104 131624 156156 131630
rect 156104 131566 156156 131572
rect 154724 130332 154776 130338
rect 154724 130274 154776 130280
rect 155472 128708 155500 131566
rect 156380 130332 156432 130338
rect 156380 130274 156432 130280
rect 156392 128708 156420 130274
rect 157312 128708 157340 139522
rect 157496 130338 157524 139658
rect 157588 138974 157616 139726
rect 158140 139450 158168 141886
rect 158876 139586 158904 141886
rect 160072 139722 160100 141886
rect 160060 139716 160112 139722
rect 160060 139658 160112 139664
rect 158864 139580 158916 139586
rect 158864 139522 158916 139528
rect 160900 139450 160928 141886
rect 162004 139586 162032 141886
rect 162280 141886 162616 141914
rect 163292 141886 163628 141914
rect 164548 141886 164608 141914
rect 162280 139858 162308 141886
rect 162268 139852 162320 139858
rect 162268 139794 162320 139800
rect 162636 139716 162688 139722
rect 162636 139658 162688 139664
rect 160980 139580 161032 139586
rect 160980 139522 161032 139528
rect 161992 139580 162044 139586
rect 161992 139522 162044 139528
rect 158128 139444 158180 139450
rect 158128 139386 158180 139392
rect 160796 139444 160848 139450
rect 160796 139386 160848 139392
rect 160888 139444 160940 139450
rect 160888 139386 160940 139392
rect 157576 138968 157628 138974
rect 157576 138910 157628 138916
rect 158220 138968 158272 138974
rect 158220 138910 158272 138916
rect 158036 138628 158088 138634
rect 158036 138570 158088 138576
rect 157484 130332 157536 130338
rect 157484 130274 157536 130280
rect 158048 128586 158076 138570
rect 158232 130338 158260 138910
rect 159968 138900 160020 138906
rect 159968 138842 160020 138848
rect 158220 130332 158272 130338
rect 158220 130274 158272 130280
rect 159048 130332 159100 130338
rect 159048 130274 159100 130280
rect 159060 128708 159088 130274
rect 159980 128708 160008 138842
rect 160808 128708 160836 139386
rect 160992 131494 161020 139522
rect 160980 131488 161032 131494
rect 160980 131430 161032 131436
rect 161716 131488 161768 131494
rect 161716 131430 161768 131436
rect 161728 128708 161756 131430
rect 162648 128708 162676 139658
rect 163004 139580 163056 139586
rect 163004 139522 163056 139528
rect 163016 130338 163044 139522
rect 163292 139382 163320 141886
rect 164580 139926 164608 141886
rect 165224 141886 165560 141914
rect 166144 141886 166480 141914
rect 167340 141886 167492 141914
rect 164568 139920 164620 139926
rect 164568 139862 164620 139868
rect 163464 139444 163516 139450
rect 163464 139386 163516 139392
rect 163280 139376 163332 139382
rect 163280 139318 163332 139324
rect 163004 130332 163056 130338
rect 163004 130274 163056 130280
rect 163476 128708 163504 139386
rect 165224 139178 165252 141886
rect 165212 139172 165264 139178
rect 165212 139114 165264 139120
rect 166144 139042 166172 141886
rect 167340 139518 167368 141886
rect 167984 141422 168012 142135
rect 168076 141886 168412 141914
rect 167972 141416 168024 141422
rect 167972 141358 168024 141364
rect 167328 139512 167380 139518
rect 167328 139454 167380 139460
rect 168076 139314 168104 141886
rect 168536 141801 168564 142174
rect 169088 141886 169424 141914
rect 170008 141886 170344 141914
rect 168522 141792 168578 141801
rect 168522 141727 168578 141736
rect 169088 139722 169116 141886
rect 170008 139790 170036 141886
rect 169996 139784 170048 139790
rect 169996 139726 170048 139732
rect 169076 139716 169128 139722
rect 169076 139658 169128 139664
rect 168064 139308 168116 139314
rect 168064 139250 168116 139256
rect 166132 139036 166184 139042
rect 166132 138978 166184 138984
rect 164384 130332 164436 130338
rect 164384 130274 164436 130280
rect 164396 128708 164424 130274
rect 158048 128558 158154 128586
rect 169996 125436 170048 125442
rect 169996 125378 170048 125384
rect 167878 118808 167934 118817
rect 167878 118743 167934 118752
rect 167892 117894 167920 118743
rect 167880 117888 167932 117894
rect 167880 117830 167932 117836
rect 146626 113232 146682 113241
rect 146626 113167 146682 113176
rect 146640 112998 146668 113167
rect 146628 112992 146680 112998
rect 146628 112934 146680 112940
rect 145340 110952 145392 110958
rect 145340 110894 145392 110900
rect 143958 108880 144014 108889
rect 143958 108815 144014 108824
rect 143972 108238 144000 108815
rect 143960 108232 144012 108238
rect 143960 108174 144012 108180
rect 164934 100040 164990 100049
rect 164934 99975 164990 99984
rect 164948 98689 164976 99975
rect 167878 98816 167934 98825
rect 167878 98751 167934 98760
rect 164934 98680 164990 98689
rect 164934 98615 164990 98624
rect 167892 98582 167920 98751
rect 167880 98576 167932 98582
rect 167880 98518 167932 98524
rect 138164 94428 138216 94434
rect 138164 94370 138216 94376
rect 142396 94428 142448 94434
rect 142396 94370 142448 94376
rect 137702 88752 137758 88761
rect 137702 88687 137758 88696
rect 137888 86064 137940 86070
rect 137888 86006 137940 86012
rect 137900 85769 137928 86006
rect 137886 85760 137942 85769
rect 137886 85695 137942 85704
rect 139636 76408 139688 76414
rect 139636 76350 139688 76356
rect 139648 75297 139676 76350
rect 142408 75682 142436 94370
rect 145798 90112 145854 90121
rect 145798 90047 145854 90056
rect 145064 86812 145116 86818
rect 145064 86754 145116 86760
rect 145076 75818 145104 86754
rect 145812 86070 145840 90047
rect 155458 88888 155514 88897
rect 149216 87158 149244 88860
rect 149768 87362 149796 88860
rect 150412 87498 150440 88860
rect 150400 87492 150452 87498
rect 150400 87434 150452 87440
rect 149756 87356 149808 87362
rect 149756 87298 149808 87304
rect 151056 87294 151084 88860
rect 151622 88846 152004 88874
rect 151044 87288 151096 87294
rect 151044 87230 151096 87236
rect 149204 87152 149256 87158
rect 149204 87094 149256 87100
rect 150584 87084 150636 87090
rect 150584 87026 150636 87032
rect 149204 87016 149256 87022
rect 149204 86958 149256 86964
rect 146444 86948 146496 86954
rect 146444 86890 146496 86896
rect 145800 86064 145852 86070
rect 145800 86006 145852 86012
rect 146456 75818 146484 86890
rect 147824 86880 147876 86886
rect 147824 86822 147876 86828
rect 147836 75818 147864 86822
rect 149216 75818 149244 86958
rect 150596 75818 150624 87026
rect 151976 78998 152004 88846
rect 152252 86138 152280 88860
rect 152910 88846 153384 88874
rect 152240 86132 152292 86138
rect 152240 86074 152292 86080
rect 153252 86132 153304 86138
rect 153252 86074 153304 86080
rect 151964 78992 152016 78998
rect 151964 78934 152016 78940
rect 151964 78856 152016 78862
rect 151964 78798 152016 78804
rect 151976 75818 152004 78798
rect 153264 78726 153292 86074
rect 153356 79082 153384 88846
rect 153448 86138 153476 88860
rect 154106 88846 154672 88874
rect 155302 88860 155458 88874
rect 154080 87492 154132 87498
rect 154080 87434 154132 87440
rect 153436 86132 153488 86138
rect 153436 86074 153488 86080
rect 153356 79054 153476 79082
rect 153344 78924 153396 78930
rect 153344 78866 153396 78872
rect 153252 78720 153304 78726
rect 153252 78662 153304 78668
rect 153356 75818 153384 78866
rect 153448 78658 153476 79054
rect 154092 78998 154120 87434
rect 154172 87356 154224 87362
rect 154172 87298 154224 87304
rect 154184 79134 154212 87298
rect 154644 81122 154672 88846
rect 154736 87498 154764 88860
rect 155288 88846 155458 88860
rect 154724 87492 154776 87498
rect 154724 87434 154776 87440
rect 155288 87401 155316 88846
rect 155458 88823 155514 88832
rect 155734 88888 155790 88897
rect 155790 88846 156144 88874
rect 155734 88823 155790 88832
rect 156116 87537 156144 88846
rect 156102 87528 156158 87537
rect 156102 87463 156158 87472
rect 155274 87392 155330 87401
rect 155274 87327 155330 87336
rect 155460 87288 155512 87294
rect 155460 87230 155512 87236
rect 154724 86132 154776 86138
rect 154724 86074 154776 86080
rect 154460 81094 154672 81122
rect 154172 79128 154224 79134
rect 154172 79070 154224 79076
rect 154080 78992 154132 78998
rect 154080 78934 154132 78940
rect 153436 78652 153488 78658
rect 153436 78594 153488 78600
rect 154460 78522 154488 81094
rect 154736 80986 154764 86074
rect 154644 80958 154764 80986
rect 154644 78590 154672 80958
rect 155472 79202 155500 87230
rect 156576 86857 156604 88860
rect 156562 86848 156618 86857
rect 156562 86783 156618 86792
rect 157220 86721 157248 88860
rect 157772 87265 157800 88860
rect 157758 87256 157814 87265
rect 157758 87191 157814 87200
rect 157576 87152 157628 87158
rect 157576 87094 157628 87100
rect 157206 86712 157262 86721
rect 157206 86647 157262 86656
rect 155460 79196 155512 79202
rect 155460 79138 155512 79144
rect 154724 79060 154776 79066
rect 154724 79002 154776 79008
rect 154632 78584 154684 78590
rect 154632 78526 154684 78532
rect 154448 78516 154500 78522
rect 154448 78458 154500 78464
rect 154736 75818 154764 79002
rect 156104 78380 156156 78386
rect 156104 78322 156156 78328
rect 156116 75818 156144 78322
rect 157588 75818 157616 87094
rect 158416 86993 158444 88860
rect 159060 87129 159088 88860
rect 159046 87120 159102 87129
rect 159046 87055 159102 87064
rect 158402 86984 158458 86993
rect 158402 86919 158458 86928
rect 159612 86818 159640 88860
rect 160256 86954 160284 88860
rect 160244 86948 160296 86954
rect 160244 86890 160296 86896
rect 160900 86886 160928 88860
rect 160980 87424 161032 87430
rect 160980 87366 161032 87372
rect 160888 86880 160940 86886
rect 160888 86822 160940 86828
rect 159600 86812 159652 86818
rect 159600 86754 159652 86760
rect 158956 79128 159008 79134
rect 158956 79070 159008 79076
rect 158968 75818 158996 79070
rect 160992 79066 161020 87366
rect 161452 87022 161480 88860
rect 162096 87090 162124 88860
rect 162464 88846 162754 88874
rect 162084 87084 162136 87090
rect 162084 87026 162136 87032
rect 161440 87016 161492 87022
rect 161440 86958 161492 86964
rect 162464 86290 162492 88846
rect 161820 86262 162492 86290
rect 161716 79196 161768 79202
rect 161716 79138 161768 79144
rect 160980 79060 161032 79066
rect 160980 79002 161032 79008
rect 160336 78992 160388 78998
rect 160336 78934 160388 78940
rect 160348 75818 160376 78934
rect 161728 75818 161756 79138
rect 161820 78862 161848 86262
rect 162360 86200 162412 86206
rect 162360 86142 162412 86148
rect 161808 78856 161860 78862
rect 161808 78798 161860 78804
rect 162372 78386 162400 86142
rect 163292 86138 163320 88860
rect 163936 87430 163964 88860
rect 163924 87424 163976 87430
rect 163924 87366 163976 87372
rect 164580 86206 164608 88860
rect 164568 86200 164620 86206
rect 164568 86142 164620 86148
rect 162452 86132 162504 86138
rect 162452 86074 162504 86080
rect 163280 86132 163332 86138
rect 163280 86074 163332 86080
rect 162464 78930 162492 86074
rect 162452 78924 162504 78930
rect 162452 78866 162504 78872
rect 163096 78788 163148 78794
rect 163096 78730 163148 78736
rect 162360 78380 162412 78386
rect 162360 78322 162412 78328
rect 163108 75818 163136 78730
rect 164568 78720 164620 78726
rect 164568 78662 164620 78668
rect 164580 75818 164608 78662
rect 165948 78652 166000 78658
rect 165948 78594 166000 78600
rect 165960 75818 165988 78594
rect 167328 78584 167380 78590
rect 167328 78526 167380 78532
rect 167340 75818 167368 78526
rect 168708 78516 168760 78522
rect 168708 78458 168760 78464
rect 168720 75818 168748 78458
rect 170008 76090 170036 125378
rect 170652 81922 170680 175698
rect 171284 144816 171336 144822
rect 171284 144758 171336 144764
rect 171296 141354 171324 144758
rect 171284 141348 171336 141354
rect 171284 141290 171336 141296
rect 170732 139240 170784 139246
rect 170732 139182 170784 139188
rect 170744 125442 170772 139182
rect 170732 125436 170784 125442
rect 170732 125378 170784 125384
rect 172032 87498 172060 225610
rect 178918 219584 178974 219593
rect 178918 219519 178974 219528
rect 178932 219282 178960 219519
rect 178920 219276 178972 219282
rect 178920 219218 178972 219224
rect 178920 203364 178972 203370
rect 178920 203306 178972 203312
rect 178932 202865 178960 203306
rect 178918 202856 178974 202865
rect 178918 202791 178974 202800
rect 173400 192620 173452 192626
rect 173400 192562 173452 192568
rect 173412 191674 173440 192562
rect 173400 191668 173452 191674
rect 173400 191610 173452 191616
rect 178920 191668 178972 191674
rect 178920 191610 178972 191616
rect 178932 186273 178960 191610
rect 178918 186264 178974 186273
rect 178918 186199 178974 186208
rect 178274 178240 178330 178249
rect 178274 178175 178330 178184
rect 182138 178240 182194 178249
rect 182194 178212 182442 178226
rect 182194 178198 182456 178212
rect 182138 178175 182194 178184
rect 178288 175830 178316 178175
rect 182428 175830 182456 178198
rect 178276 175824 178328 175830
rect 178276 175766 178328 175772
rect 182416 175824 182468 175830
rect 182876 175824 182928 175830
rect 182416 175766 182468 175772
rect 182874 175792 182876 175801
rect 182928 175792 182930 175801
rect 189512 175762 189540 177940
rect 182874 175727 182930 175736
rect 189500 175756 189552 175762
rect 189500 175698 189552 175704
rect 196688 175694 196716 177940
rect 196676 175688 196728 175694
rect 196676 175630 196728 175636
rect 190604 175212 190656 175218
rect 190604 175154 190656 175160
rect 176160 175144 176212 175150
rect 176160 175086 176212 175092
rect 173582 169128 173638 169137
rect 173582 169063 173638 169072
rect 173398 167768 173454 167777
rect 173398 167703 173454 167712
rect 173306 164912 173362 164921
rect 173306 164847 173362 164856
rect 172848 161544 172900 161550
rect 172848 161486 172900 161492
rect 172860 156625 172888 161486
rect 172846 156616 172902 156625
rect 172846 156551 172902 156560
rect 172940 153928 172992 153934
rect 172940 153870 172992 153876
rect 172952 153769 172980 153870
rect 172938 153760 172994 153769
rect 173320 153730 173348 164847
rect 173412 155022 173440 167703
rect 173490 166408 173546 166417
rect 173490 166343 173546 166352
rect 173400 155016 173452 155022
rect 173400 154958 173452 154964
rect 172938 153695 172994 153704
rect 173308 153724 173360 153730
rect 173308 153666 173360 153672
rect 173504 153662 173532 166343
rect 173596 156450 173624 169063
rect 174042 163552 174098 163561
rect 174042 163487 174098 163496
rect 173674 162192 173730 162201
rect 173674 162127 173730 162136
rect 173584 156444 173636 156450
rect 173584 156386 173636 156392
rect 173492 153656 173544 153662
rect 173492 153598 173544 153604
rect 173216 153180 173268 153186
rect 173216 153122 173268 153128
rect 173228 152409 173256 153122
rect 173214 152400 173270 152409
rect 173214 152335 173270 152344
rect 173688 150942 173716 162127
rect 173950 160696 174006 160705
rect 173950 160631 173952 160640
rect 174004 160631 174006 160640
rect 173952 160602 174004 160608
rect 173952 159368 174004 159374
rect 173950 159336 173952 159345
rect 174004 159336 174006 159345
rect 173950 159271 174006 159280
rect 173860 158008 173912 158014
rect 173766 157976 173822 157985
rect 173860 157950 173912 157956
rect 173766 157911 173768 157920
rect 173820 157911 173822 157920
rect 173768 157882 173820 157888
rect 173768 156512 173820 156518
rect 173768 156454 173820 156460
rect 173676 150936 173728 150942
rect 173676 150878 173728 150884
rect 173780 145337 173808 156454
rect 173872 146697 173900 157950
rect 174056 155242 174084 163487
rect 174056 155214 174176 155242
rect 173952 155152 174004 155158
rect 173952 155094 174004 155100
rect 174042 155120 174098 155129
rect 173858 146688 173914 146697
rect 173858 146623 173914 146632
rect 173766 145328 173822 145337
rect 173766 145263 173822 145272
rect 173964 143977 173992 155094
rect 174042 155055 174044 155064
rect 174096 155055 174098 155064
rect 174044 155026 174096 155032
rect 174148 154970 174176 155214
rect 174056 154942 174176 154970
rect 174056 152370 174084 154942
rect 174044 152364 174096 152370
rect 174044 152306 174096 152312
rect 174042 150904 174098 150913
rect 174042 150839 174098 150848
rect 174056 150806 174084 150839
rect 174044 150800 174096 150806
rect 174044 150742 174096 150748
rect 174042 149544 174098 149553
rect 174042 149479 174044 149488
rect 174096 149479 174098 149488
rect 174044 149450 174096 149456
rect 174044 148216 174096 148222
rect 174042 148184 174044 148193
rect 174096 148184 174098 148193
rect 174042 148119 174098 148128
rect 173950 143968 174006 143977
rect 173950 143903 174006 143912
rect 173582 142608 173638 142617
rect 173582 142543 173638 142552
rect 173596 142034 173624 142543
rect 173584 142028 173636 142034
rect 173584 141970 173636 141976
rect 175514 125472 175570 125481
rect 175514 125407 175516 125416
rect 175568 125407 175570 125416
rect 175516 125378 175568 125384
rect 173400 98576 173452 98582
rect 173400 98518 173452 98524
rect 173412 92598 173440 98518
rect 173400 92592 173452 92598
rect 173400 92534 173452 92540
rect 175516 92592 175568 92598
rect 175516 92534 175568 92540
rect 175528 92297 175556 92534
rect 175514 92288 175570 92297
rect 175514 92223 175570 92232
rect 172020 87492 172072 87498
rect 172020 87434 172072 87440
rect 170640 81916 170692 81922
rect 170640 81858 170692 81864
rect 176172 81854 176200 175086
rect 190616 163946 190644 175154
rect 196688 175150 196716 175630
rect 203772 175218 203800 177940
rect 203760 175212 203812 175218
rect 203760 175154 203812 175160
rect 196676 175144 196728 175150
rect 196676 175086 196728 175092
rect 210948 166990 210976 177940
rect 218032 175529 218060 177940
rect 218018 175520 218074 175529
rect 218018 175455 218074 175464
rect 222160 168616 222212 168622
rect 222160 168558 222212 168564
rect 203852 166984 203904 166990
rect 203852 166926 203904 166932
rect 210936 166984 210988 166990
rect 210936 166926 210988 166932
rect 190616 163918 190736 163946
rect 190708 163674 190736 163918
rect 203864 163796 203892 166926
rect 217192 166848 217244 166854
rect 217192 166790 217244 166796
rect 217204 163796 217232 166790
rect 190538 163646 190736 163674
rect 179012 163448 179064 163454
rect 182324 163448 182376 163454
rect 179012 163390 179064 163396
rect 182322 163416 182324 163425
rect 182376 163416 182378 163425
rect 178828 162088 178880 162094
rect 178828 162030 178880 162036
rect 177540 160660 177592 160666
rect 177540 160602 177592 160608
rect 176252 157940 176304 157946
rect 176252 157882 176304 157888
rect 176264 149582 176292 157882
rect 177552 150874 177580 160602
rect 178840 153934 178868 162030
rect 178920 159300 178972 159306
rect 178920 159242 178972 159248
rect 178828 153928 178880 153934
rect 178828 153870 178880 153876
rect 177540 150868 177592 150874
rect 177540 150810 177592 150816
rect 176252 149576 176304 149582
rect 176252 149518 176304 149524
rect 178932 149514 178960 159242
rect 179024 155090 179052 163390
rect 182322 163351 182378 163360
rect 181770 162464 181826 162473
rect 181770 162399 181826 162408
rect 181784 162094 181812 162399
rect 181772 162088 181824 162094
rect 181772 162030 181824 162036
rect 182322 161648 182378 161657
rect 182322 161583 182378 161592
rect 181678 160696 181734 160705
rect 179104 160660 179156 160666
rect 182336 160666 182364 161583
rect 181678 160631 181734 160640
rect 182324 160660 182376 160666
rect 179104 160602 179156 160608
rect 179012 155084 179064 155090
rect 179012 155026 179064 155032
rect 179116 153186 179144 160602
rect 180392 159368 180444 159374
rect 180392 159310 180444 159316
rect 180298 158384 180354 158393
rect 180298 158319 180354 158328
rect 179104 153180 179156 153186
rect 179104 153122 179156 153128
rect 178920 149508 178972 149514
rect 178920 149450 178972 149456
rect 180312 148222 180340 158319
rect 180404 148601 180432 159310
rect 181128 155084 181180 155090
rect 181128 155026 181180 155032
rect 181140 154721 181168 155026
rect 181126 154712 181182 154721
rect 181126 154647 181182 154656
rect 181404 153724 181456 153730
rect 181404 153666 181456 153672
rect 181416 153225 181444 153666
rect 181402 153216 181458 153225
rect 181402 153151 181458 153160
rect 181036 150800 181088 150806
rect 181036 150742 181088 150748
rect 181048 150670 181076 150742
rect 181692 150670 181720 160631
rect 182324 160602 182376 160608
rect 182322 159880 182378 159889
rect 182322 159815 182378 159824
rect 182336 159306 182364 159815
rect 182324 159300 182376 159306
rect 182324 159242 182376 159248
rect 182322 158112 182378 158121
rect 182322 158047 182378 158056
rect 182336 157946 182364 158047
rect 182324 157940 182376 157946
rect 182324 157882 182376 157888
rect 181770 157160 181826 157169
rect 181770 157095 181826 157104
rect 181784 156518 181812 157095
rect 181772 156512 181824 156518
rect 181772 156454 181824 156460
rect 182324 156444 182376 156450
rect 182324 156386 182376 156392
rect 182230 156344 182286 156353
rect 182230 156279 182286 156288
rect 182244 155158 182272 156279
rect 182336 156081 182364 156386
rect 182322 156072 182378 156081
rect 182322 156007 182378 156016
rect 182232 155152 182284 155158
rect 182232 155094 182284 155100
rect 181956 153656 182008 153662
rect 181954 153624 181956 153633
rect 182008 153624 182010 153633
rect 181954 153559 182010 153568
rect 182324 152364 182376 152370
rect 182324 152306 182376 152312
rect 182336 152137 182364 152306
rect 182322 152128 182378 152137
rect 182322 152063 182378 152072
rect 182324 150936 182376 150942
rect 182322 150904 182324 150913
rect 182376 150904 182378 150913
rect 182232 150868 182284 150874
rect 182322 150839 182378 150848
rect 182232 150810 182284 150816
rect 181036 150664 181088 150670
rect 181036 150606 181088 150612
rect 181680 150664 181732 150670
rect 182244 150641 182272 150810
rect 181680 150606 181732 150612
rect 182230 150632 182286 150641
rect 182230 150567 182286 150576
rect 182324 149576 182376 149582
rect 182324 149518 182376 149524
rect 180390 148592 180446 148601
rect 180390 148527 180446 148536
rect 182336 148329 182364 149518
rect 182322 148320 182378 148329
rect 182322 148255 182378 148264
rect 180300 148216 180352 148222
rect 180300 148158 180352 148164
rect 185648 145434 185676 147884
rect 185636 145428 185688 145434
rect 185636 145370 185688 145376
rect 189236 144822 189264 147884
rect 189224 144816 189276 144822
rect 189224 144758 189276 144764
rect 185084 144748 185136 144754
rect 185084 144690 185136 144696
rect 185096 133740 185124 144690
rect 192916 144657 192944 147884
rect 192902 144648 192958 144657
rect 192902 144583 192958 144592
rect 196504 144113 196532 147884
rect 197504 144816 197556 144822
rect 197504 144758 197556 144764
rect 196490 144104 196546 144113
rect 196490 144039 196546 144048
rect 196858 144104 196914 144113
rect 196858 144039 196914 144048
rect 196872 142238 196900 144039
rect 196860 142232 196912 142238
rect 196860 142174 196912 142180
rect 197516 133740 197544 144758
rect 197686 143968 197742 143977
rect 197686 143903 197742 143912
rect 197700 135137 197728 143903
rect 200184 142306 200212 147884
rect 203772 144521 203800 147884
rect 207452 147762 207480 147884
rect 207268 147734 207480 147762
rect 203758 144512 203814 144521
rect 203758 144447 203814 144456
rect 203772 143394 203800 144447
rect 203760 143388 203812 143394
rect 203760 143330 203812 143336
rect 200172 142300 200224 142306
rect 200172 142242 200224 142248
rect 200184 141937 200212 142242
rect 200170 141928 200226 141937
rect 200170 141863 200226 141872
rect 207268 141121 207296 147734
rect 211040 143462 211068 147884
rect 214720 144754 214748 147884
rect 218308 144822 218336 147884
rect 218296 144816 218348 144822
rect 218296 144758 218348 144764
rect 221988 144754 222016 147884
rect 222172 145434 222200 168558
rect 225208 166854 225236 177940
rect 225840 168956 225892 168962
rect 225840 168898 225892 168904
rect 225196 166848 225248 166854
rect 225196 166790 225248 166796
rect 225748 164808 225800 164814
rect 225748 164750 225800 164756
rect 222436 161612 222488 161618
rect 222436 161554 222488 161560
rect 222448 157146 222476 161554
rect 225654 160696 225710 160705
rect 225654 160631 225710 160640
rect 225564 159980 225616 159986
rect 225564 159922 225616 159928
rect 222804 157192 222856 157198
rect 222448 157140 222804 157146
rect 222448 157134 222856 157140
rect 222448 157118 222844 157134
rect 222160 145428 222212 145434
rect 222160 145370 222212 145376
rect 214708 144748 214760 144754
rect 214708 144690 214760 144696
rect 218940 144748 218992 144754
rect 218940 144690 218992 144696
rect 221976 144748 222028 144754
rect 221976 144690 222028 144696
rect 211028 143456 211080 143462
rect 211028 143398 211080 143404
rect 211040 143161 211068 143398
rect 211026 143152 211082 143161
rect 211026 143087 211082 143096
rect 207254 141112 207310 141121
rect 207254 141047 207310 141056
rect 207268 140606 207296 141047
rect 207256 140600 207308 140606
rect 207256 140542 207308 140548
rect 218952 136730 218980 144690
rect 219674 142064 219730 142073
rect 219674 141999 219676 142008
rect 219728 141999 219730 142008
rect 219676 141970 219728 141976
rect 210016 136724 210068 136730
rect 210016 136666 210068 136672
rect 218940 136724 218992 136730
rect 218940 136666 218992 136672
rect 197686 135128 197742 135137
rect 197686 135063 197742 135072
rect 210028 133740 210056 136666
rect 222448 133754 222476 157118
rect 225576 151010 225604 159922
rect 225564 151004 225616 151010
rect 225564 150946 225616 150952
rect 225668 150942 225696 160631
rect 225760 152681 225788 164750
rect 225852 155401 225880 168898
rect 226024 167596 226076 167602
rect 226024 167538 226076 167544
rect 225932 166236 225984 166242
rect 225932 166178 225984 166184
rect 225838 155392 225894 155401
rect 225838 155327 225894 155336
rect 225944 153633 225972 166178
rect 226036 154449 226064 167538
rect 226300 163516 226352 163522
rect 226300 163458 226352 163464
rect 226116 163448 226168 163454
rect 226312 163425 226340 163458
rect 226116 163390 226168 163396
rect 226298 163416 226354 163425
rect 226022 154440 226078 154449
rect 226022 154375 226078 154384
rect 225930 153624 225986 153633
rect 225930 153559 225986 153568
rect 225746 152672 225802 152681
rect 225746 152607 225802 152616
rect 226128 151865 226156 163390
rect 226298 163351 226354 163360
rect 226298 162464 226354 162473
rect 226298 162399 226300 162408
rect 226352 162399 226354 162408
rect 226300 162370 226352 162376
rect 226300 162088 226352 162094
rect 226300 162030 226352 162036
rect 226312 159986 226340 162030
rect 226390 161648 226446 161657
rect 226390 161583 226446 161592
rect 226404 160666 226432 161583
rect 226392 160660 226444 160666
rect 226392 160602 226444 160608
rect 226300 159980 226352 159986
rect 226300 159922 226352 159928
rect 226298 159880 226354 159889
rect 226298 159815 226354 159824
rect 226312 159374 226340 159815
rect 226300 159368 226352 159374
rect 226300 159310 226352 159316
rect 227220 159300 227272 159306
rect 227220 159242 227272 159248
rect 226390 158928 226446 158937
rect 226390 158863 226446 158872
rect 226298 158112 226354 158121
rect 226298 158047 226354 158056
rect 226114 151856 226170 151865
rect 226114 151791 226170 151800
rect 226208 151004 226260 151010
rect 226208 150946 226260 150952
rect 225656 150936 225708 150942
rect 226220 150913 226248 150946
rect 225656 150878 225708 150884
rect 226206 150904 226262 150913
rect 225564 150868 225616 150874
rect 226206 150839 226262 150848
rect 225564 150810 225616 150816
rect 225576 150097 225604 150810
rect 225562 150088 225618 150097
rect 225562 150023 225618 150032
rect 225288 149440 225340 149446
rect 225288 149382 225340 149388
rect 225300 149145 225328 149382
rect 225286 149136 225342 149145
rect 225286 149071 225342 149080
rect 225196 148692 225248 148698
rect 225196 148634 225248 148640
rect 225208 148329 225236 148634
rect 225194 148320 225250 148329
rect 225194 148255 225250 148264
rect 226312 146794 226340 158047
rect 226404 158014 226432 158863
rect 226392 158008 226444 158014
rect 226392 157950 226444 157956
rect 226390 157160 226446 157169
rect 226390 157095 226446 157104
rect 226300 146788 226352 146794
rect 226300 146730 226352 146736
rect 226404 145434 226432 157095
rect 226482 156344 226538 156353
rect 226482 156279 226538 156288
rect 226392 145428 226444 145434
rect 226392 145370 226444 145376
rect 226496 144074 226524 156279
rect 227232 149446 227260 159242
rect 227312 157940 227364 157946
rect 227312 157882 227364 157888
rect 227220 149440 227272 149446
rect 227220 149382 227272 149388
rect 227324 148698 227352 157882
rect 227312 148692 227364 148698
rect 227312 148634 227364 148640
rect 226484 144068 226536 144074
rect 226484 144010 226536 144016
rect 222448 133726 222554 133754
rect 176252 117888 176304 117894
rect 176252 117830 176304 117836
rect 176264 108889 176292 117830
rect 176250 108880 176306 108889
rect 176250 108815 176306 108824
rect 178734 84264 178790 84273
rect 178734 84199 178790 84208
rect 182322 84264 182378 84273
rect 182378 84236 182442 84250
rect 182378 84222 182456 84236
rect 182322 84199 182378 84208
rect 178748 81990 178776 84199
rect 182428 81990 182456 84222
rect 178736 81984 178788 81990
rect 178736 81926 178788 81932
rect 182416 81984 182468 81990
rect 182416 81926 182468 81932
rect 189512 81922 189540 83828
rect 189500 81916 189552 81922
rect 189500 81858 189552 81864
rect 196688 81854 196716 83828
rect 176160 81848 176212 81854
rect 176160 81790 176212 81796
rect 196676 81848 196728 81854
rect 196676 81790 196728 81796
rect 203772 81310 203800 83828
rect 190604 81304 190656 81310
rect 190604 81246 190656 81252
rect 203760 81304 203812 81310
rect 203760 81246 203812 81252
rect 173860 76408 173912 76414
rect 173860 76350 173912 76356
rect 170008 76062 170082 76090
rect 144952 75790 145104 75818
rect 146332 75790 146484 75818
rect 147712 75790 147864 75818
rect 149092 75790 149244 75818
rect 150564 75790 150624 75818
rect 151944 75790 152004 75818
rect 153324 75790 153384 75818
rect 154704 75790 154764 75818
rect 156084 75790 156144 75818
rect 157556 75790 157616 75818
rect 158936 75790 158996 75818
rect 160316 75790 160376 75818
rect 161696 75790 161756 75818
rect 163076 75790 163136 75818
rect 164548 75790 164608 75818
rect 165928 75790 165988 75818
rect 167308 75790 167368 75818
rect 168688 75790 168748 75818
rect 170054 75804 170082 76062
rect 142408 75654 143572 75682
rect 173872 75297 173900 76350
rect 139634 75288 139690 75297
rect 139634 75223 139690 75232
rect 173858 75288 173914 75297
rect 173858 75223 173914 75232
rect 174042 74200 174098 74209
rect 174042 74135 174098 74144
rect 139726 73792 139782 73801
rect 174056 73762 174084 74135
rect 139726 73727 139782 73736
rect 174044 73756 174096 73762
rect 139542 72568 139598 72577
rect 139542 72503 139598 72512
rect 139556 69478 139584 72503
rect 139634 71072 139690 71081
rect 139634 71007 139690 71016
rect 139648 70974 139676 71007
rect 139636 70968 139688 70974
rect 139636 70910 139688 70916
rect 139740 69546 139768 73727
rect 174044 73698 174096 73704
rect 181036 73756 181088 73762
rect 181036 73698 181088 73704
rect 172938 73248 172994 73257
rect 172938 73183 172994 73192
rect 172952 72402 172980 73183
rect 172940 72396 172992 72402
rect 172940 72338 172992 72344
rect 180944 72396 180996 72402
rect 180944 72338 180996 72344
rect 173306 72160 173362 72169
rect 173306 72095 173362 72104
rect 139910 71480 139966 71489
rect 139910 71415 139966 71424
rect 139818 69576 139874 69585
rect 139728 69540 139780 69546
rect 139818 69511 139874 69520
rect 139728 69482 139780 69488
rect 139544 69472 139596 69478
rect 139544 69414 139596 69420
rect 139634 68352 139690 68361
rect 139634 68287 139690 68296
rect 139648 68254 139676 68287
rect 136784 68248 136836 68254
rect 136784 68190 136836 68196
rect 139636 68248 139688 68254
rect 139636 68190 139688 68196
rect 135956 66888 136008 66894
rect 135956 66830 136008 66836
rect 135968 65330 135996 66830
rect 136140 66820 136192 66826
rect 136140 66762 136192 66768
rect 135956 65324 136008 65330
rect 135956 65266 136008 65272
rect 136152 64038 136180 66762
rect 136796 65398 136824 68190
rect 139726 67400 139782 67409
rect 139726 67335 139782 67344
rect 139634 67128 139690 67137
rect 139634 67063 139690 67072
rect 139648 66826 139676 67063
rect 139740 66894 139768 67335
rect 139728 66888 139780 66894
rect 139728 66830 139780 66836
rect 139636 66820 139688 66826
rect 139636 66762 139688 66768
rect 139832 66758 139860 69511
rect 139924 68186 139952 71415
rect 173320 70974 173348 72095
rect 174042 71072 174098 71081
rect 174042 71007 174044 71016
rect 174096 71007 174098 71016
rect 178460 71036 178512 71042
rect 174044 70978 174096 70984
rect 178460 70978 178512 70984
rect 173308 70968 173360 70974
rect 173308 70910 173360 70916
rect 178276 70968 178328 70974
rect 178276 70910 178328 70916
rect 174042 70120 174098 70129
rect 174042 70055 174098 70064
rect 174056 69954 174084 70055
rect 174044 69948 174096 69954
rect 174044 69890 174096 69896
rect 172938 69032 172994 69041
rect 172938 68967 172994 68976
rect 172952 68254 172980 68967
rect 172940 68248 172992 68254
rect 172940 68190 172992 68196
rect 178288 68186 178316 70910
rect 178368 69948 178420 69954
rect 178368 69890 178420 69896
rect 139912 68180 139964 68186
rect 139912 68122 139964 68128
rect 178276 68180 178328 68186
rect 178276 68122 178328 68128
rect 173858 67944 173914 67953
rect 173858 67879 173914 67888
rect 173400 67568 173452 67574
rect 173400 67510 173452 67516
rect 139820 66752 139872 66758
rect 139820 66694 139872 66700
rect 139910 65496 139966 65505
rect 139910 65431 139966 65440
rect 136784 65392 136836 65398
rect 136784 65334 136836 65340
rect 139634 64272 139690 64281
rect 139634 64207 139690 64216
rect 136140 64032 136192 64038
rect 136140 63974 136192 63980
rect 139648 62610 139676 64207
rect 139726 63184 139782 63193
rect 139726 63119 139782 63128
rect 139636 62604 139688 62610
rect 139636 62546 139688 62552
rect 139634 61416 139690 61425
rect 139634 61351 139690 61360
rect 139648 59822 139676 61351
rect 139740 61250 139768 63119
rect 139818 62776 139874 62785
rect 139818 62711 139874 62720
rect 139728 61244 139780 61250
rect 139728 61186 139780 61192
rect 139726 60056 139782 60065
rect 139726 59991 139782 60000
rect 139636 59816 139688 59822
rect 139636 59758 139688 59764
rect 139740 58530 139768 59991
rect 139832 59890 139860 62711
rect 139924 62542 139952 65431
rect 139912 62536 139964 62542
rect 139912 62478 139964 62484
rect 173122 61824 173178 61833
rect 173122 61759 173178 61768
rect 173136 61658 173164 61759
rect 173124 61652 173176 61658
rect 173124 61594 173176 61600
rect 173122 60736 173178 60745
rect 173122 60671 173178 60680
rect 173136 60570 173164 60671
rect 173124 60564 173176 60570
rect 173124 60506 173176 60512
rect 139820 59884 139872 59890
rect 139820 59826 139872 59832
rect 173030 59648 173086 59657
rect 173030 59583 173086 59592
rect 140462 58968 140518 58977
rect 140462 58903 140518 58912
rect 140370 58696 140426 58705
rect 140370 58631 140426 58640
rect 139728 58524 139780 58530
rect 139728 58466 139780 58472
rect 140278 57200 140334 57209
rect 140278 57135 140334 57144
rect 136508 55804 136560 55810
rect 136508 55746 136560 55752
rect 136520 54382 136548 55746
rect 140292 55742 140320 57135
rect 140384 57102 140412 58631
rect 140372 57096 140424 57102
rect 140372 57038 140424 57044
rect 140476 57034 140504 58903
rect 173044 58802 173072 59583
rect 173032 58796 173084 58802
rect 173032 58738 173084 58744
rect 173306 57608 173362 57617
rect 173306 57543 173362 57552
rect 173320 57170 173348 57543
rect 173308 57164 173360 57170
rect 173308 57106 173360 57112
rect 140464 57028 140516 57034
rect 140464 56970 140516 56976
rect 140462 56248 140518 56257
rect 140462 56183 140518 56192
rect 140476 55810 140504 56183
rect 140464 55804 140516 55810
rect 140464 55746 140516 55752
rect 140280 55736 140332 55742
rect 140280 55678 140332 55684
rect 173412 55577 173440 67510
rect 173872 66826 173900 67879
rect 174042 66992 174098 67001
rect 174042 66927 174044 66936
rect 174096 66927 174098 66936
rect 174044 66898 174096 66904
rect 173860 66820 173912 66826
rect 173860 66762 173912 66768
rect 178380 66486 178408 69890
rect 178368 66480 178420 66486
rect 178368 66422 178420 66428
rect 178472 66214 178500 70978
rect 180956 68497 180984 72338
rect 181048 69449 181076 73698
rect 190616 69834 190644 81246
rect 210948 73014 210976 83828
rect 218032 76414 218060 83828
rect 225208 80630 225236 83828
rect 224460 80624 224512 80630
rect 224460 80566 224512 80572
rect 225196 80624 225248 80630
rect 225196 80566 225248 80572
rect 218020 76408 218072 76414
rect 218020 76350 218072 76356
rect 224472 73014 224500 80566
rect 226576 73756 226628 73762
rect 226576 73698 226628 73704
rect 204128 73008 204180 73014
rect 204128 72950 204180 72956
rect 210936 73008 210988 73014
rect 210936 72950 210988 72956
rect 217560 73008 217612 73014
rect 217560 72950 217612 72956
rect 224460 73008 224512 73014
rect 224460 72950 224512 72956
rect 204140 69834 204168 72950
rect 217572 69834 217600 72950
rect 190538 69806 190644 69834
rect 203878 69806 204168 69834
rect 217218 69806 217600 69834
rect 225932 69540 225984 69546
rect 225932 69482 225984 69488
rect 181034 69440 181090 69449
rect 181034 69375 181090 69384
rect 225944 68497 225972 69482
rect 226482 69440 226538 69449
rect 226588 69426 226616 73698
rect 226538 69398 226616 69426
rect 226482 69375 226538 69384
rect 180942 68488 180998 68497
rect 180942 68423 180998 68432
rect 225930 68488 225986 68497
rect 225930 68423 225986 68432
rect 180944 68248 180996 68254
rect 180944 68190 180996 68196
rect 179104 66956 179156 66962
rect 179104 66898 179156 66904
rect 178460 66208 178512 66214
rect 178460 66150 178512 66156
rect 173858 65904 173914 65913
rect 173858 65839 173914 65848
rect 173872 65738 173900 65839
rect 173860 65732 173912 65738
rect 173860 65674 173912 65680
rect 178828 65732 178880 65738
rect 178828 65674 178880 65680
rect 173490 64952 173546 64961
rect 173490 64887 173492 64896
rect 173544 64887 173546 64896
rect 175884 64916 175936 64922
rect 173492 64858 173544 64864
rect 175884 64858 175936 64864
rect 173490 63864 173546 63873
rect 173490 63799 173546 63808
rect 173504 62678 173532 63799
rect 174042 62776 174098 62785
rect 174042 62711 174044 62720
rect 174096 62711 174098 62720
rect 174044 62682 174096 62688
rect 173492 62672 173544 62678
rect 173492 62614 173544 62620
rect 175608 62672 175660 62678
rect 175608 62614 175660 62620
rect 175516 61652 175568 61658
rect 175516 61594 175568 61600
rect 175528 59890 175556 61594
rect 175620 61250 175648 62614
rect 175896 62610 175924 64858
rect 178276 62740 178328 62746
rect 178276 62682 178328 62688
rect 175884 62604 175936 62610
rect 175884 62546 175936 62552
rect 175608 61244 175660 61250
rect 175608 61186 175660 61192
rect 175792 60564 175844 60570
rect 175792 60506 175844 60512
rect 175516 59884 175568 59890
rect 175516 59826 175568 59832
rect 175700 58796 175752 58802
rect 175700 58738 175752 58744
rect 173582 58696 173638 58705
rect 173582 58631 173584 58640
rect 173636 58631 173638 58640
rect 175608 58660 175660 58666
rect 173584 58602 173636 58608
rect 175608 58602 175660 58608
rect 175516 57164 175568 57170
rect 175516 57106 175568 57112
rect 173490 56656 173546 56665
rect 173490 56591 173546 56600
rect 173504 56082 173532 56591
rect 173492 56076 173544 56082
rect 173492 56018 173544 56024
rect 175528 55742 175556 57106
rect 175620 56626 175648 58602
rect 175608 56620 175660 56626
rect 175608 56562 175660 56568
rect 175712 56558 175740 58738
rect 175804 58530 175832 60506
rect 178288 59754 178316 62682
rect 178840 62542 178868 65674
rect 179116 64038 179144 66898
rect 180956 64417 180984 68190
rect 181404 68180 181456 68186
rect 181404 68122 181456 68128
rect 226300 68180 226352 68186
rect 226300 68122 226352 68128
rect 181416 67681 181444 68122
rect 226312 67681 226340 68122
rect 181402 67672 181458 67681
rect 181402 67607 181458 67616
rect 226298 67672 226354 67681
rect 226298 67607 226354 67616
rect 223448 67568 223500 67574
rect 223448 67510 223500 67516
rect 181772 66820 181824 66826
rect 181772 66762 181824 66768
rect 180942 64408 180998 64417
rect 180942 64343 180998 64352
rect 181784 64145 181812 66762
rect 182140 66480 182192 66486
rect 181954 66448 182010 66457
rect 182140 66422 182192 66428
rect 181954 66383 182010 66392
rect 181968 66214 181996 66383
rect 181956 66208 182008 66214
rect 181956 66150 182008 66156
rect 182152 65913 182180 66422
rect 182138 65904 182194 65913
rect 182138 65839 182194 65848
rect 181770 64136 181826 64145
rect 181770 64071 181826 64080
rect 179104 64032 179156 64038
rect 179104 63974 179156 63980
rect 182324 64032 182376 64038
rect 182324 63974 182376 63980
rect 182336 63193 182364 63974
rect 182322 63184 182378 63193
rect 182322 63119 182378 63128
rect 181588 62604 181640 62610
rect 181588 62546 181640 62552
rect 178828 62536 178880 62542
rect 178828 62478 178880 62484
rect 181600 61425 181628 62546
rect 182324 62536 182376 62542
rect 182324 62478 182376 62484
rect 182336 62377 182364 62478
rect 182322 62368 182378 62377
rect 182322 62303 182378 62312
rect 181586 61416 181642 61425
rect 181586 61351 181642 61360
rect 181220 61244 181272 61250
rect 181220 61186 181272 61192
rect 181232 60473 181260 61186
rect 181218 60464 181274 60473
rect 181218 60399 181274 60408
rect 181128 59884 181180 59890
rect 181128 59826 181180 59832
rect 178276 59748 178328 59754
rect 178276 59690 178328 59696
rect 181036 59748 181088 59754
rect 181036 59690 181088 59696
rect 181048 59657 181076 59690
rect 181034 59648 181090 59657
rect 181034 59583 181090 59592
rect 181140 58705 181168 59826
rect 181126 58696 181182 58705
rect 181126 58631 181182 58640
rect 175792 58524 175844 58530
rect 175792 58466 175844 58472
rect 181036 58524 181088 58530
rect 181036 58466 181088 58472
rect 181048 57889 181076 58466
rect 181034 57880 181090 57889
rect 181034 57815 181090 57824
rect 181034 56656 181090 56665
rect 181034 56591 181090 56600
rect 181128 56620 181180 56626
rect 181048 56558 181076 56591
rect 181128 56562 181180 56568
rect 175700 56552 175752 56558
rect 175700 56494 175752 56500
rect 181036 56552 181088 56558
rect 181036 56494 181088 56500
rect 181140 56121 181168 56562
rect 181126 56112 181182 56121
rect 175608 56076 175660 56082
rect 181126 56047 181182 56056
rect 175608 56018 175660 56024
rect 175516 55736 175568 55742
rect 175516 55678 175568 55684
rect 173398 55568 173454 55577
rect 173398 55503 173454 55512
rect 140646 55296 140702 55305
rect 140646 55231 140702 55240
rect 140660 55062 140688 55231
rect 140648 55056 140700 55062
rect 140648 54998 140700 55004
rect 140370 54480 140426 54489
rect 140370 54415 140372 54424
rect 140424 54415 140426 54424
rect 173582 54480 173638 54489
rect 173582 54415 173584 54424
rect 140372 54386 140424 54392
rect 173636 54415 173638 54424
rect 173584 54386 173636 54392
rect 136508 54376 136560 54382
rect 136508 54318 136560 54324
rect 175620 54246 175648 56018
rect 181036 55736 181088 55742
rect 181036 55678 181088 55684
rect 181048 55169 181076 55678
rect 181034 55160 181090 55169
rect 181034 55095 181090 55104
rect 223460 55062 223488 67510
rect 226392 66752 226444 66758
rect 226298 66720 226354 66729
rect 226392 66694 226444 66700
rect 226298 66655 226300 66664
rect 226352 66655 226354 66664
rect 226300 66626 226352 66632
rect 226404 65913 226432 66694
rect 226390 65904 226446 65913
rect 226390 65839 226446 65848
rect 225932 65392 225984 65398
rect 225932 65334 225984 65340
rect 225944 64145 225972 65334
rect 226208 65324 226260 65330
rect 226208 65266 226260 65272
rect 226220 64961 226248 65266
rect 226206 64952 226262 64961
rect 226206 64887 226262 64896
rect 225930 64136 225986 64145
rect 225930 64071 225986 64080
rect 225748 64032 225800 64038
rect 225748 63974 225800 63980
rect 225760 63193 225788 63974
rect 225746 63184 225802 63193
rect 225746 63119 225802 63128
rect 226300 62604 226352 62610
rect 226300 62546 226352 62552
rect 226312 62377 226340 62546
rect 226298 62368 226354 62377
rect 226298 62303 226354 62312
rect 226300 61448 226352 61454
rect 226298 61416 226300 61425
rect 226352 61416 226354 61425
rect 226298 61351 226354 61360
rect 225748 61244 225800 61250
rect 225748 61186 225800 61192
rect 225760 60473 225788 61186
rect 225746 60464 225802 60473
rect 225746 60399 225802 60408
rect 226300 59884 226352 59890
rect 226300 59826 226352 59832
rect 226312 59657 226340 59826
rect 226298 59648 226354 59657
rect 226298 59583 226354 59592
rect 225748 59476 225800 59482
rect 225748 59418 225800 59424
rect 225760 58705 225788 59418
rect 225746 58696 225802 58705
rect 225746 58631 225802 58640
rect 225564 58524 225616 58530
rect 225564 58466 225616 58472
rect 225576 57889 225604 58466
rect 225562 57880 225618 57889
rect 225562 57815 225618 57824
rect 226300 57096 226352 57102
rect 226300 57038 226352 57044
rect 225656 57028 225708 57034
rect 225656 56970 225708 56976
rect 225668 56121 225696 56970
rect 226312 56937 226340 57038
rect 226298 56928 226354 56937
rect 226298 56863 226354 56872
rect 225654 56112 225710 56121
rect 225654 56047 225710 56056
rect 226484 55804 226536 55810
rect 226484 55746 226536 55752
rect 226392 55736 226444 55742
rect 226392 55678 226444 55684
rect 226404 55169 226432 55678
rect 226390 55160 226446 55169
rect 226390 55095 226446 55104
rect 223448 55056 223500 55062
rect 223448 54998 223500 55004
rect 181034 54344 181090 54353
rect 181034 54279 181090 54288
rect 181048 54246 181076 54279
rect 175608 54240 175660 54246
rect 175608 54182 175660 54188
rect 181036 54240 181088 54246
rect 181036 54182 181088 54188
rect 217560 54172 217612 54178
rect 217560 54114 217612 54120
rect 140556 53696 140608 53702
rect 140556 53638 140608 53644
rect 173584 53696 173636 53702
rect 173584 53638 173636 53644
rect 140568 53537 140596 53638
rect 173596 53537 173624 53638
rect 140554 53528 140610 53537
rect 140554 53463 140610 53472
rect 173582 53528 173638 53537
rect 173582 53463 173638 53472
rect 140004 53016 140056 53022
rect 140004 52958 140056 52964
rect 171836 53016 171888 53022
rect 171836 52958 171888 52964
rect 140016 52449 140044 52958
rect 171848 52449 171876 52958
rect 140002 52440 140058 52449
rect 140002 52375 140058 52384
rect 171834 52440 171890 52449
rect 171834 52375 171890 52384
rect 134760 51588 134812 51594
rect 134760 51530 134812 51536
rect 185004 51526 185032 53908
rect 187304 51594 187332 53908
rect 187292 51588 187344 51594
rect 187292 51530 187344 51536
rect 184992 51520 185044 51526
rect 184992 51462 185044 51468
rect 173306 51352 173362 51361
rect 173306 51287 173362 51296
rect 142854 51080 142910 51089
rect 142854 51015 142910 51024
rect 140646 50808 140702 50817
rect 140646 50743 140702 50752
rect 140370 50400 140426 50409
rect 140660 50370 140688 50743
rect 140370 50335 140426 50344
rect 140648 50364 140700 50370
rect 140384 50302 140412 50335
rect 140648 50306 140700 50312
rect 140372 50296 140424 50302
rect 140372 50238 140424 50244
rect 140554 49040 140610 49049
rect 140554 48975 140610 48984
rect 140568 48942 140596 48975
rect 140556 48936 140608 48942
rect 140556 48878 140608 48884
rect 140002 48088 140058 48097
rect 140002 48023 140058 48032
rect 140016 47718 140044 48023
rect 140004 47712 140056 47718
rect 140004 47654 140056 47660
rect 142868 47582 142896 51015
rect 170456 50976 170508 50982
rect 170456 50918 170508 50924
rect 170468 50658 170496 50918
rect 170546 50672 170602 50681
rect 170192 50630 170546 50658
rect 147730 48088 147786 48097
rect 147436 48046 147730 48074
rect 153986 48088 154042 48097
rect 150564 48046 150624 48074
rect 147730 48023 147786 48032
rect 144400 47910 144736 47938
rect 142856 47576 142908 47582
rect 142856 47518 142908 47524
rect 144708 46018 144736 47910
rect 144696 46012 144748 46018
rect 144696 45954 144748 45960
rect 150596 45882 150624 48046
rect 153448 48046 153986 48074
rect 153448 45950 153476 48046
rect 153986 48023 154042 48032
rect 165960 48046 166448 48074
rect 160058 47952 160114 47961
rect 156820 47910 156880 47938
rect 156852 47514 156880 47910
rect 159520 47910 160058 47938
rect 159520 47582 159548 47910
rect 162984 47910 163044 47938
rect 160058 47887 160114 47896
rect 159508 47576 159560 47582
rect 159508 47518 159560 47524
rect 156840 47508 156892 47514
rect 156840 47450 156892 47456
rect 163016 46601 163044 47910
rect 163002 46592 163058 46601
rect 163002 46527 163058 46536
rect 153436 45944 153488 45950
rect 153436 45886 153488 45892
rect 150584 45876 150636 45882
rect 150584 45818 150636 45824
rect 163016 45785 163044 46527
rect 165960 45921 165988 48046
rect 166420 47825 166448 48046
rect 168890 47952 168946 47961
rect 168946 47910 169576 47938
rect 168890 47887 168946 47896
rect 166406 47816 166462 47825
rect 166406 47751 166462 47760
rect 167234 47816 167290 47825
rect 167234 47751 167290 47760
rect 167248 46086 167276 47751
rect 167694 47544 167750 47553
rect 167694 47479 167696 47488
rect 167748 47479 167750 47488
rect 167696 47450 167748 47456
rect 167236 46080 167288 46086
rect 169548 46057 169576 47910
rect 169720 46080 169772 46086
rect 167236 46022 167288 46028
rect 169534 46048 169590 46057
rect 169534 45983 169590 45992
rect 169718 46048 169720 46057
rect 169772 46048 169774 46057
rect 169718 45983 169774 45992
rect 165946 45912 166002 45921
rect 165946 45847 166002 45856
rect 163002 45776 163058 45785
rect 163002 45711 163058 45720
rect 169548 45406 169576 45983
rect 169536 45400 169588 45406
rect 169536 45342 169588 45348
rect 169732 44794 169760 45983
rect 170192 45882 170220 50630
rect 170546 50607 170602 50616
rect 173320 50370 173348 51287
rect 185084 50908 185136 50914
rect 185084 50850 185136 50856
rect 173582 50400 173638 50409
rect 173308 50364 173360 50370
rect 173582 50335 173638 50344
rect 173308 50306 173360 50312
rect 173596 50302 173624 50335
rect 173584 50296 173636 50302
rect 173584 50238 173636 50244
rect 182140 49548 182192 49554
rect 182140 49490 182192 49496
rect 182152 49321 182180 49490
rect 172938 49312 172994 49321
rect 182138 49312 182194 49321
rect 172938 49247 172994 49256
rect 181968 49270 182138 49298
rect 172952 48942 172980 49247
rect 172940 48936 172992 48942
rect 172940 48878 172992 48884
rect 173306 48360 173362 48369
rect 173306 48295 173362 48304
rect 173320 47514 173348 48295
rect 181864 48188 181916 48194
rect 181864 48130 181916 48136
rect 181876 47961 181904 48130
rect 181862 47952 181918 47961
rect 181862 47887 181918 47896
rect 173308 47508 173360 47514
rect 173308 47450 173360 47456
rect 181968 46442 181996 49270
rect 182138 49247 182194 49256
rect 182232 48188 182284 48194
rect 182232 48130 182284 48136
rect 182138 46728 182194 46737
rect 182138 46663 182194 46672
rect 181876 46414 181996 46442
rect 170180 45876 170232 45882
rect 170180 45818 170232 45824
rect 169720 44788 169772 44794
rect 169720 44730 169772 44736
rect 129160 40702 129464 40730
rect 126388 36628 126440 36634
rect 126388 36570 126440 36576
rect 127124 36628 127176 36634
rect 127124 36570 127176 36576
rect 126400 34746 126428 36570
rect 91132 34718 91284 34746
rect 93616 34718 93676 34746
rect 96100 34718 96436 34746
rect 98584 34718 98644 34746
rect 101068 34718 101404 34746
rect 103552 34718 103612 34746
rect 106128 34718 106464 34746
rect 108612 34718 108672 34746
rect 111096 34718 111432 34746
rect 113580 34718 113640 34746
rect 116064 34718 116124 34746
rect 118640 34718 118700 34746
rect 121124 34718 121460 34746
rect 123608 34718 123852 34746
rect 126092 34718 126428 34746
rect 129160 34610 129188 40702
rect 128576 34582 129188 34610
rect 88484 32956 88536 32962
rect 88484 32898 88536 32904
rect 88390 26056 88446 26065
rect 88390 25991 88446 26000
rect 88022 23336 88078 23345
rect 88022 23271 88078 23280
rect 88496 20761 88524 32898
rect 181876 23345 181904 46414
rect 181956 45400 182008 45406
rect 181954 45368 181956 45377
rect 182048 45400 182100 45406
rect 182008 45368 182010 45377
rect 182048 45342 182100 45348
rect 181954 45303 182010 45312
rect 181968 33681 181996 45303
rect 182060 44794 182088 45342
rect 182048 44788 182100 44794
rect 182048 44730 182100 44736
rect 181954 33672 182010 33681
rect 181954 33607 182010 33616
rect 182060 30825 182088 44730
rect 182046 30816 182102 30825
rect 182046 30751 182102 30760
rect 182152 28105 182180 46663
rect 182138 28096 182194 28105
rect 182138 28031 182194 28040
rect 182244 26065 182272 48130
rect 185096 34732 185124 50850
rect 187304 50681 187332 51530
rect 189696 50982 189724 53908
rect 191996 51633 192024 53908
rect 191982 51624 192038 51633
rect 191982 51559 192038 51568
rect 189684 50976 189736 50982
rect 189684 50918 189736 50924
rect 190604 50976 190656 50982
rect 190604 50918 190656 50924
rect 187290 50672 187346 50681
rect 187290 50607 187346 50616
rect 187568 47508 187620 47514
rect 187568 47450 187620 47456
rect 187580 34732 187608 47450
rect 190616 34610 190644 50918
rect 194388 49554 194416 53908
rect 196124 51044 196176 51050
rect 196124 50986 196176 50992
rect 194376 49548 194428 49554
rect 194376 49490 194428 49496
rect 192536 48936 192588 48942
rect 192536 48878 192588 48884
rect 192548 34732 192576 48878
rect 196136 37450 196164 50986
rect 196688 48194 196716 53908
rect 197504 50296 197556 50302
rect 197504 50238 197556 50244
rect 196676 48188 196728 48194
rect 196676 48130 196728 48136
rect 195020 37444 195072 37450
rect 195020 37386 195072 37392
rect 196124 37444 196176 37450
rect 196124 37386 196176 37392
rect 195032 34732 195060 37386
rect 197516 34732 197544 50238
rect 199080 46737 199108 53908
rect 200264 51112 200316 51118
rect 200264 51054 200316 51060
rect 199066 46728 199122 46737
rect 199066 46663 199122 46672
rect 200276 34746 200304 51054
rect 201472 45406 201500 53908
rect 203772 51633 203800 53908
rect 203758 51624 203814 51633
rect 203758 51559 203814 51568
rect 205784 51180 205836 51186
rect 205784 51122 205836 51128
rect 202564 50364 202616 50370
rect 202564 50306 202616 50312
rect 201460 45400 201512 45406
rect 201460 45342 201512 45348
rect 200106 34718 200304 34746
rect 202576 34732 202604 50306
rect 205796 44674 205824 51122
rect 206164 50914 206192 53908
rect 207900 53288 207952 53294
rect 207900 53230 207952 53236
rect 207912 51361 207940 53230
rect 207898 51352 207954 51361
rect 207898 51287 207954 51296
rect 208464 50982 208492 53908
rect 210856 51050 210884 53908
rect 212500 53696 212552 53702
rect 212500 53638 212552 53644
rect 212512 53129 212540 53638
rect 212498 53120 212554 53129
rect 212498 53055 212554 53064
rect 213248 51118 213276 53908
rect 215548 51186 215576 53908
rect 215536 51180 215588 51186
rect 215536 51122 215588 51128
rect 213236 51112 213288 51118
rect 213236 51054 213288 51060
rect 210844 51044 210896 51050
rect 210844 50986 210896 50992
rect 208452 50976 208504 50982
rect 208452 50918 208504 50924
rect 206152 50908 206204 50914
rect 206152 50850 206204 50856
rect 211304 50432 211356 50438
rect 211304 50374 211356 50380
rect 205612 44646 205824 44674
rect 205612 35154 205640 44646
rect 211316 37790 211344 50374
rect 212590 47408 212646 47417
rect 212590 47343 212646 47352
rect 210016 37784 210068 37790
rect 207530 37752 207586 37761
rect 210016 37726 210068 37732
rect 211304 37784 211356 37790
rect 211304 37726 211356 37732
rect 207530 37687 207586 37696
rect 205520 35126 205640 35154
rect 205520 34746 205548 35126
rect 205074 34718 205548 34746
rect 207544 34732 207572 37687
rect 210028 34732 210056 37726
rect 212604 34732 212632 47343
rect 215076 37784 215128 37790
rect 215076 37726 215128 37732
rect 215088 34732 215116 37726
rect 217572 34732 217600 54114
rect 217940 50438 217968 53908
rect 220240 50982 220268 53908
rect 222632 51458 222660 53908
rect 220964 51452 221016 51458
rect 220964 51394 221016 51400
rect 222620 51452 222672 51458
rect 222620 51394 222672 51400
rect 218940 50976 218992 50982
rect 218940 50918 218992 50924
rect 220228 50976 220280 50982
rect 220228 50918 220280 50924
rect 217928 50432 217980 50438
rect 217928 50374 217980 50380
rect 218952 37790 218980 50918
rect 220976 37790 221004 51394
rect 223460 44674 223488 54998
rect 226496 54353 226524 55746
rect 226482 54344 226538 54353
rect 226482 54279 226538 54288
rect 223092 44646 223488 44674
rect 218940 37784 218992 37790
rect 218940 37726 218992 37732
rect 220044 37784 220096 37790
rect 220044 37726 220096 37732
rect 220964 37784 221016 37790
rect 220964 37726 221016 37732
rect 220056 34732 220084 37726
rect 223092 35154 223120 44646
rect 223000 35126 223120 35154
rect 223000 34746 223028 35126
rect 222554 34718 223028 34746
rect 190078 34582 190644 34610
rect 182324 33024 182376 33030
rect 182324 32966 182376 32972
rect 182230 26056 182286 26065
rect 182230 25991 182286 26000
rect 181862 23336 181918 23345
rect 181862 23271 181918 23280
rect 182336 20761 182364 32966
rect 88482 20752 88538 20761
rect 88482 20687 88538 20696
rect 182322 20752 182378 20761
rect 182322 20687 182378 20696
rect 92420 18942 92664 18970
rect 92636 16846 92664 18942
rect 96868 18942 97388 18970
rect 102356 18942 102416 18970
rect 92624 16840 92676 16846
rect 92624 16782 92676 16788
rect 80756 16772 80808 16778
rect 80756 16714 80808 16720
rect 67876 16704 67928 16710
rect 67876 16646 67928 16652
rect 54996 16636 55048 16642
rect 54996 16578 55048 16584
rect 29236 16568 29288 16574
rect 29236 16510 29288 16516
rect 16356 16432 16408 16438
rect 16356 16374 16408 16380
rect 13044 15616 13096 15622
rect 13042 15584 13044 15593
rect 16080 15616 16132 15622
rect 13096 15584 13098 15593
rect 16080 15558 16132 15564
rect 13042 15519 13098 15528
rect 16368 9304 16396 16374
rect 29248 9304 29276 16510
rect 42116 16500 42168 16506
rect 42116 16442 42168 16448
rect 42128 9304 42156 16442
rect 55008 9304 55036 16578
rect 67888 9304 67916 16646
rect 80768 9304 80796 16714
rect 96868 12290 96896 18942
rect 102388 16778 102416 18942
rect 107080 18942 107416 18970
rect 112048 18942 112384 18970
rect 117016 18942 117352 18970
rect 122076 18942 122412 18970
rect 127228 18942 127380 18970
rect 105136 16840 105188 16846
rect 105136 16782 105188 16788
rect 102376 16772 102428 16778
rect 102376 16714 102428 16720
rect 105148 12358 105176 16782
rect 107080 16710 107108 18942
rect 107068 16704 107120 16710
rect 107068 16646 107120 16652
rect 112048 16642 112076 18942
rect 112036 16636 112088 16642
rect 112036 16578 112088 16584
rect 117016 16506 117044 18942
rect 122076 16574 122104 18942
rect 122064 16568 122116 16574
rect 122064 16510 122116 16516
rect 117004 16500 117056 16506
rect 117004 16442 117056 16448
rect 119396 16500 119448 16506
rect 119396 16442 119448 16448
rect 105136 12352 105188 12358
rect 105136 12294 105188 12300
rect 106516 12352 106568 12358
rect 106516 12294 106568 12300
rect 93636 12284 93688 12290
rect 93636 12226 93688 12232
rect 96856 12284 96908 12290
rect 96856 12226 96908 12232
rect 93648 9304 93676 12226
rect 106528 9304 106556 12294
rect 119408 9304 119436 16442
rect 127228 16438 127256 18942
rect 186384 17118 186412 18956
rect 191352 17118 191380 18956
rect 196320 17118 196348 18956
rect 185176 17112 185228 17118
rect 185176 17054 185228 17060
rect 186372 17112 186424 17118
rect 186372 17054 186424 17060
rect 191340 17112 191392 17118
rect 191340 17054 191392 17060
rect 192076 17112 192128 17118
rect 192076 17054 192128 17060
rect 196124 17112 196176 17118
rect 196124 17054 196176 17060
rect 196308 17112 196360 17118
rect 196308 17054 196360 17060
rect 170916 16704 170968 16710
rect 170916 16646 170968 16652
rect 158036 16636 158088 16642
rect 158036 16578 158088 16584
rect 145156 16568 145208 16574
rect 145156 16510 145208 16516
rect 127216 16432 127268 16438
rect 127216 16374 127268 16380
rect 132276 16432 132328 16438
rect 132276 16374 132328 16380
rect 132288 9304 132316 16374
rect 145168 9304 145196 16510
rect 158048 9304 158076 16578
rect 170928 9304 170956 16646
rect 183796 12352 183848 12358
rect 183796 12294 183848 12300
rect 183808 9304 183836 12294
rect 185188 12290 185216 17054
rect 185176 12284 185228 12290
rect 185176 12226 185228 12232
rect 192088 12154 192116 17054
rect 196136 12358 196164 17054
rect 201380 16710 201408 18956
rect 201368 16704 201420 16710
rect 201368 16646 201420 16652
rect 206348 16642 206376 18956
rect 206336 16636 206388 16642
rect 206336 16578 206388 16584
rect 211316 16574 211344 18956
rect 211304 16568 211356 16574
rect 211304 16510 211356 16516
rect 216376 16438 216404 18956
rect 221344 16506 221372 18956
rect 221332 16500 221384 16506
rect 221332 16442 221384 16448
rect 216364 16432 216416 16438
rect 216364 16374 216416 16380
rect 222436 16432 222488 16438
rect 222436 16374 222488 16380
rect 196124 12352 196176 12358
rect 196124 12294 196176 12300
rect 209556 12284 209608 12290
rect 209556 12226 209608 12232
rect 192076 12148 192128 12154
rect 192076 12090 192128 12096
rect 196676 12148 196728 12154
rect 196676 12090 196728 12096
rect 196688 9304 196716 12090
rect 209568 9304 209596 12226
rect 222448 9304 222476 16374
rect 228612 12290 228640 388538
rect 231004 388346 231032 396206
rect 249036 395198 249064 396206
rect 266608 396206 266728 396234
rect 249024 395192 249076 395198
rect 249024 395134 249076 395140
rect 266608 392426 266636 396206
rect 284364 393809 284392 396344
rect 284350 393800 284406 393809
rect 284350 393735 284406 393744
rect 299440 393288 299492 393294
rect 299440 393230 299492 393236
rect 266608 392398 266728 392426
rect 265860 388528 265912 388534
rect 265860 388470 265912 388476
rect 230912 388318 231032 388346
rect 230912 382822 230940 388318
rect 249116 385604 249168 385610
rect 249116 385546 249168 385552
rect 230900 382816 230952 382822
rect 230900 382758 230952 382764
rect 249128 378826 249156 385546
rect 249036 378798 249156 378826
rect 249036 375954 249064 378798
rect 248932 375948 248984 375954
rect 248932 375890 248984 375896
rect 249024 375948 249076 375954
rect 249024 375890 249076 375896
rect 248944 375206 248972 375890
rect 228784 375200 228836 375206
rect 228784 375142 228836 375148
rect 248932 375200 248984 375206
rect 248932 375142 248984 375148
rect 228692 333788 228744 333794
rect 228692 333730 228744 333736
rect 228704 262666 228732 333730
rect 228796 332978 228824 375142
rect 229980 371800 230032 371806
rect 229980 371742 230032 371748
rect 228784 332972 228836 332978
rect 228784 332914 228836 332920
rect 228692 262660 228744 262666
rect 228692 262602 228744 262608
rect 228692 255928 228744 255934
rect 228692 255870 228744 255876
rect 228704 245258 228732 255870
rect 228692 245252 228744 245258
rect 228692 245194 228744 245200
rect 229992 232338 230020 371742
rect 233476 357928 233528 357934
rect 233476 357870 233528 357876
rect 233488 357769 233516 357870
rect 233474 357760 233530 357769
rect 233474 357695 233530 357704
rect 233476 356568 233528 356574
rect 233474 356536 233476 356545
rect 233528 356536 233530 356545
rect 233474 356471 233530 356480
rect 233476 355208 233528 355214
rect 233474 355176 233476 355185
rect 233528 355176 233530 355185
rect 233474 355111 233530 355120
rect 233568 355140 233620 355146
rect 233568 355082 233620 355088
rect 233580 354641 233608 355082
rect 233566 354632 233622 354641
rect 233566 354567 233622 354576
rect 233476 353848 233528 353854
rect 233476 353790 233528 353796
rect 233488 353553 233516 353790
rect 233474 353544 233530 353553
rect 233474 353479 233530 353488
rect 233476 352420 233528 352426
rect 233476 352362 233528 352368
rect 233488 352329 233516 352362
rect 233474 352320 233530 352329
rect 233474 352255 233530 352264
rect 231636 351332 231688 351338
rect 231636 351274 231688 351280
rect 231176 349768 231228 349774
rect 231176 349710 231228 349716
rect 231188 348278 231216 349710
rect 231648 349706 231676 351274
rect 233568 351060 233620 351066
rect 233568 351002 233620 351008
rect 233476 350992 233528 350998
rect 233474 350960 233476 350969
rect 233528 350960 233530 350969
rect 233474 350895 233530 350904
rect 233580 350425 233608 351002
rect 233566 350416 233622 350425
rect 233566 350351 233622 350360
rect 231636 349700 231688 349706
rect 231636 349642 231688 349648
rect 233476 349700 233528 349706
rect 233476 349642 233528 349648
rect 233488 349609 233516 349642
rect 233474 349600 233530 349609
rect 233474 349535 233530 349544
rect 233292 348408 233344 348414
rect 233292 348350 233344 348356
rect 231176 348272 231228 348278
rect 231176 348214 231228 348220
rect 233304 346481 233332 348350
rect 233384 348340 233436 348346
rect 233384 348282 233436 348288
rect 233396 346889 233424 348282
rect 233476 348272 233528 348278
rect 233474 348240 233476 348249
rect 233528 348240 233530 348249
rect 233474 348175 233530 348184
rect 233382 346880 233438 346889
rect 233382 346815 233438 346824
rect 233290 346472 233346 346481
rect 233290 346407 233346 346416
rect 234580 345620 234632 345626
rect 234580 345562 234632 345568
rect 233476 345552 233528 345558
rect 233476 345494 233528 345500
rect 233488 345257 233516 345494
rect 233474 345248 233530 345257
rect 233474 345183 233530 345192
rect 234488 344260 234540 344266
rect 234488 344202 234540 344208
rect 234396 344192 234448 344198
rect 234396 344134 234448 344140
rect 233476 344124 233528 344130
rect 233476 344066 233528 344072
rect 233488 344033 233516 344066
rect 233474 344024 233530 344033
rect 233474 343959 233530 343968
rect 230532 342832 230584 342838
rect 230532 342774 230584 342780
rect 230544 340050 230572 342774
rect 232004 341540 232056 341546
rect 232004 341482 232056 341488
rect 231820 341472 231872 341478
rect 231820 341414 231872 341420
rect 230532 340044 230584 340050
rect 230532 339986 230584 339992
rect 231832 338554 231860 341414
rect 231912 338752 231964 338758
rect 231912 338694 231964 338700
rect 231820 338548 231872 338554
rect 231820 338490 231872 338496
rect 231544 337664 231596 337670
rect 231544 337606 231596 337612
rect 230716 335964 230768 335970
rect 230716 335906 230768 335912
rect 230728 333114 230756 335906
rect 231556 334134 231584 337606
rect 231924 335902 231952 338694
rect 232016 338622 232044 341482
rect 234408 341313 234436 344134
rect 234500 342265 234528 344202
rect 234592 342673 234620 345562
rect 234578 342664 234634 342673
rect 234578 342599 234634 342608
rect 234486 342256 234542 342265
rect 234486 342191 234542 342200
rect 234394 341304 234450 341313
rect 234394 341239 234450 341248
rect 233568 340112 233620 340118
rect 233568 340054 233620 340060
rect 233476 340044 233528 340050
rect 233476 339986 233528 339992
rect 233488 339953 233516 339986
rect 233474 339944 233530 339953
rect 233474 339879 233530 339888
rect 232004 338616 232056 338622
rect 233476 338616 233528 338622
rect 232004 338558 232056 338564
rect 233474 338584 233476 338593
rect 233528 338584 233530 338593
rect 233474 338519 233530 338528
rect 233580 337097 233608 340054
rect 234120 338684 234172 338690
rect 234120 338626 234172 338632
rect 233660 338548 233712 338554
rect 233660 338490 233712 338496
rect 233672 338185 233700 338490
rect 233658 338176 233714 338185
rect 233658 338111 233714 338120
rect 233566 337088 233622 337097
rect 233566 337023 233622 337032
rect 231912 335896 231964 335902
rect 233476 335896 233528 335902
rect 231912 335838 231964 335844
rect 233474 335864 233476 335873
rect 233528 335864 233530 335873
rect 233474 335799 233530 335808
rect 234132 334377 234160 338626
rect 234118 334368 234174 334377
rect 234118 334303 234174 334312
rect 231544 334128 231596 334134
rect 231544 334070 231596 334076
rect 234304 334128 234356 334134
rect 234304 334070 234356 334076
rect 234316 333969 234344 334070
rect 234302 333960 234358 333969
rect 234302 333895 234358 333904
rect 230992 333584 231044 333590
rect 231820 333584 231872 333590
rect 230992 333526 231044 333532
rect 231818 333552 231820 333561
rect 231872 333552 231874 333561
rect 230716 333108 230768 333114
rect 230716 333050 230768 333056
rect 230898 332192 230954 332201
rect 230898 332127 230954 332136
rect 230806 331512 230862 331521
rect 230806 331447 230862 331456
rect 230716 326988 230768 326994
rect 230716 326930 230768 326936
rect 230728 298473 230756 326930
rect 230820 307857 230848 331447
rect 230912 310985 230940 332127
rect 231004 320369 231032 333526
rect 231818 333487 231874 333496
rect 231360 333176 231412 333182
rect 231360 333118 231412 333124
rect 231372 332201 231400 333118
rect 233936 333108 233988 333114
rect 233936 333050 233988 333056
rect 233948 333017 233976 333050
rect 233934 333008 233990 333017
rect 231452 332972 231504 332978
rect 233934 332943 233990 332952
rect 231452 332914 231504 332920
rect 231358 332192 231414 332201
rect 231358 332127 231414 332136
rect 231464 331521 231492 332914
rect 233476 331748 233528 331754
rect 233476 331690 233528 331696
rect 233488 331521 233516 331690
rect 231450 331512 231506 331521
rect 231450 331447 231506 331456
rect 233474 331512 233530 331521
rect 233474 331447 233530 331456
rect 231728 330660 231780 330666
rect 231728 330602 231780 330608
rect 231740 329034 231768 330602
rect 233474 330288 233530 330297
rect 233474 330223 233530 330232
rect 233488 329238 233516 330223
rect 252610 330152 252666 330161
rect 252666 330110 252776 330138
rect 252610 330087 252666 330096
rect 251966 330016 252022 330025
rect 251856 329974 251966 330002
rect 251966 329951 252022 329960
rect 236248 329838 237412 329866
rect 238332 329838 238668 329866
rect 239252 329838 239588 329866
rect 233476 329232 233528 329238
rect 233476 329174 233528 329180
rect 231360 329028 231412 329034
rect 231360 328970 231412 328976
rect 231728 329028 231780 329034
rect 231728 328970 231780 328976
rect 230990 320360 231046 320369
rect 230990 320295 231046 320304
rect 231372 314113 231400 328970
rect 231452 328960 231504 328966
rect 231452 328902 231504 328908
rect 231464 327606 231492 328902
rect 231452 327600 231504 327606
rect 231452 327542 231504 327548
rect 231464 317241 231492 327542
rect 232004 327464 232056 327470
rect 232004 327406 232056 327412
rect 232016 326994 232044 327406
rect 232096 327124 232148 327130
rect 232096 327066 232148 327072
rect 232004 326988 232056 326994
rect 232004 326930 232056 326936
rect 231450 317232 231506 317241
rect 231450 317167 231506 317176
rect 231358 314104 231414 314113
rect 231358 314039 231414 314048
rect 230898 310976 230954 310985
rect 230898 310911 230954 310920
rect 231452 309716 231504 309722
rect 231452 309658 231504 309664
rect 230806 307848 230862 307857
rect 230806 307783 230862 307792
rect 230714 298464 230770 298473
rect 230714 298399 230770 298408
rect 230806 294656 230862 294665
rect 230806 294591 230862 294600
rect 230072 253208 230124 253214
rect 230072 253150 230124 253156
rect 230084 243150 230112 253150
rect 230164 251780 230216 251786
rect 230164 251722 230216 251728
rect 230072 243144 230124 243150
rect 230072 243086 230124 243092
rect 230176 242946 230204 251722
rect 230164 242940 230216 242946
rect 230164 242882 230216 242888
rect 230714 234408 230770 234417
rect 230714 234343 230770 234352
rect 230728 234145 230756 234343
rect 230714 234136 230770 234145
rect 230714 234071 230770 234080
rect 229980 232332 230032 232338
rect 229980 232274 230032 232280
rect 228692 225396 228744 225402
rect 228692 225338 228744 225344
rect 228704 51526 228732 225338
rect 230728 223265 230756 234071
rect 230714 223256 230770 223265
rect 230714 223191 230770 223200
rect 230820 200689 230848 294591
rect 231082 289080 231138 289089
rect 231082 289015 231138 289024
rect 230900 238588 230952 238594
rect 230900 238530 230952 238536
rect 230912 237953 230940 238530
rect 230898 237944 230954 237953
rect 230898 237879 230954 237888
rect 230912 217009 230940 237879
rect 230992 235868 231044 235874
rect 230992 235810 231044 235816
rect 231004 235194 231032 235810
rect 230992 235188 231044 235194
rect 230992 235130 231044 235136
rect 231004 220137 231032 235130
rect 230990 220128 231046 220137
rect 230990 220063 231046 220072
rect 230898 217000 230954 217009
rect 230898 216935 230954 216944
rect 230806 200680 230862 200689
rect 230806 200615 230862 200624
rect 230714 197552 230770 197561
rect 230714 197487 230770 197496
rect 228784 158008 228836 158014
rect 228784 157950 228836 157956
rect 228796 148222 228824 157950
rect 228784 148216 228836 148222
rect 228784 148158 228836 148164
rect 230728 104401 230756 197487
rect 230820 107937 230848 200615
rect 231096 194977 231124 289015
rect 231358 285272 231414 285281
rect 231358 285207 231414 285216
rect 231174 234952 231230 234961
rect 231174 234887 231230 234896
rect 231188 234553 231216 234887
rect 231174 234544 231230 234553
rect 231174 234479 231230 234488
rect 231188 226393 231216 234479
rect 231174 226384 231230 226393
rect 231174 226319 231230 226328
rect 231372 226218 231400 285207
rect 231464 279705 231492 309658
rect 232002 304720 232058 304729
rect 232108 304706 232136 327066
rect 233476 327056 233528 327062
rect 233476 326998 233528 327004
rect 232058 304678 232136 304706
rect 232002 304655 232058 304664
rect 232108 304214 232136 304678
rect 232096 304208 232148 304214
rect 232096 304150 232148 304156
rect 232740 304208 232792 304214
rect 232740 304150 232792 304156
rect 232002 301592 232058 301601
rect 232002 301527 232058 301536
rect 232016 301426 232044 301527
rect 232004 301420 232056 301426
rect 232004 301362 232056 301368
rect 231544 295912 231596 295918
rect 231544 295854 231596 295860
rect 231450 279696 231506 279705
rect 231450 279631 231506 279640
rect 231556 276577 231584 295854
rect 231820 283536 231872 283542
rect 231820 283478 231872 283484
rect 231634 282824 231690 282833
rect 231634 282759 231636 282768
rect 231688 282759 231690 282768
rect 231636 282730 231688 282736
rect 231832 282674 231860 283478
rect 231648 282646 231860 282674
rect 231542 276568 231598 276577
rect 231542 276503 231598 276512
rect 231648 273449 231676 282646
rect 232752 274401 232780 304150
rect 233488 301426 233516 326998
rect 233476 301420 233528 301426
rect 233476 301362 233528 301368
rect 234120 301420 234172 301426
rect 234120 301362 234172 301368
rect 234132 275110 234160 301362
rect 236248 283066 236276 329838
rect 238640 327198 238668 329838
rect 239560 327538 239588 329838
rect 239928 329838 240264 329866
rect 241184 329838 241520 329866
rect 242196 329838 242532 329866
rect 239548 327532 239600 327538
rect 239548 327474 239600 327480
rect 238628 327192 238680 327198
rect 238628 327134 238680 327140
rect 239928 326858 239956 329838
rect 238996 326852 239048 326858
rect 238996 326794 239048 326800
rect 239916 326852 239968 326858
rect 239916 326794 239968 326800
rect 239008 319990 239036 326794
rect 241492 326654 241520 329838
rect 241756 327396 241808 327402
rect 241756 327338 241808 327344
rect 241480 326648 241532 326654
rect 241480 326590 241532 326596
rect 241768 320058 241796 327338
rect 242504 326518 242532 329838
rect 242780 329838 243116 329866
rect 244128 329838 244372 329866
rect 245048 329838 245384 329866
rect 246060 329838 246396 329866
rect 246980 329838 247224 329866
rect 247992 329838 248328 329866
rect 248912 329838 249156 329866
rect 242780 327402 242808 329838
rect 242768 327396 242820 327402
rect 242768 327338 242820 327344
rect 244240 327124 244292 327130
rect 244240 327066 244292 327072
rect 242492 326512 242544 326518
rect 242492 326454 242544 326460
rect 244252 326314 244280 327066
rect 244344 326450 244372 329838
rect 244424 327192 244476 327198
rect 244424 327134 244476 327140
rect 244332 326444 244384 326450
rect 244332 326386 244384 326392
rect 243228 326308 243280 326314
rect 243228 326250 243280 326256
rect 244240 326308 244292 326314
rect 244240 326250 244292 326256
rect 243240 320670 243268 326250
rect 243228 320664 243280 320670
rect 243228 320606 243280 320612
rect 243780 320664 243832 320670
rect 243780 320606 243832 320612
rect 243596 320528 243648 320534
rect 243596 320470 243648 320476
rect 241756 320052 241808 320058
rect 241756 319994 241808 320000
rect 238996 319984 239048 319990
rect 238996 319926 239048 319932
rect 243608 316810 243636 320470
rect 243300 316782 243636 316810
rect 243792 316810 243820 320606
rect 244436 320602 244464 327134
rect 244516 326376 244568 326382
rect 244516 326318 244568 326324
rect 244424 320596 244476 320602
rect 244424 320538 244476 320544
rect 244528 316810 244556 326318
rect 245356 326314 245384 329838
rect 245896 326852 245948 326858
rect 245896 326794 245948 326800
rect 245344 326308 245396 326314
rect 245344 326250 245396 326256
rect 245908 320670 245936 326794
rect 246368 326586 246396 329838
rect 247196 327198 247224 329838
rect 247184 327192 247236 327198
rect 247184 327134 247236 327140
rect 248300 326994 248328 329838
rect 248840 327532 248892 327538
rect 248840 327474 248892 327480
rect 248288 326988 248340 326994
rect 248288 326930 248340 326936
rect 247276 326784 247328 326790
rect 247276 326726 247328 326732
rect 246356 326580 246408 326586
rect 246356 326522 246408 326528
rect 245896 320664 245948 320670
rect 245896 320606 245948 320612
rect 246448 320664 246500 320670
rect 246448 320606 246500 320612
rect 246264 320188 246316 320194
rect 246264 320130 246316 320136
rect 246276 316810 246304 320130
rect 243792 316782 244128 316810
rect 244528 316782 245048 316810
rect 245968 316782 246304 316810
rect 246460 316810 246488 320606
rect 247288 316810 247316 326726
rect 248656 326716 248708 326722
rect 248656 326658 248708 326664
rect 248668 320534 248696 326658
rect 248748 326308 248800 326314
rect 248748 326250 248800 326256
rect 248656 320528 248708 320534
rect 248656 320470 248708 320476
rect 248760 320330 248788 326250
rect 248748 320324 248800 320330
rect 248748 320266 248800 320272
rect 248852 319718 248880 327474
rect 249128 327470 249156 329838
rect 249588 329838 249924 329866
rect 250508 329838 250844 329866
rect 253728 329838 253788 329866
rect 254372 329838 254708 329866
rect 255720 329838 256056 329866
rect 249588 327538 249616 329838
rect 250508 327538 250536 329838
rect 253728 329034 253756 329838
rect 253716 329028 253768 329034
rect 253716 328970 253768 328976
rect 254372 327606 254400 329838
rect 254360 327600 254412 327606
rect 256028 327577 256056 329838
rect 256304 329838 256640 329866
rect 257316 329838 257652 329866
rect 258420 329838 258572 329866
rect 259248 329838 259584 329866
rect 260168 329838 260504 329866
rect 261180 329838 261516 329866
rect 262100 329838 262436 329866
rect 263112 329838 263448 329866
rect 264124 329838 264368 329866
rect 254360 327542 254412 327548
rect 256014 327568 256070 327577
rect 249576 327532 249628 327538
rect 249576 327474 249628 327480
rect 250496 327532 250548 327538
rect 256014 327503 256070 327512
rect 250496 327474 250548 327480
rect 249116 327464 249168 327470
rect 249116 327406 249168 327412
rect 248932 327396 248984 327402
rect 248932 327338 248984 327344
rect 248944 320602 248972 327338
rect 249588 327062 249616 327474
rect 250508 327266 250536 327474
rect 256304 327402 256332 329838
rect 256292 327396 256344 327402
rect 256292 327338 256344 327344
rect 250496 327260 250548 327266
rect 250496 327202 250548 327208
rect 257316 327130 257344 329838
rect 258420 327266 258448 329838
rect 258408 327260 258460 327266
rect 258408 327202 258460 327208
rect 258960 327192 259012 327198
rect 258960 327134 259012 327140
rect 257304 327124 257356 327130
rect 257304 327066 257356 327072
rect 249576 327056 249628 327062
rect 249576 326998 249628 327004
rect 250036 327056 250088 327062
rect 250036 326998 250088 327004
rect 248932 320596 248984 320602
rect 248932 320538 248984 320544
rect 249116 320528 249168 320534
rect 249116 320470 249168 320476
rect 248932 320120 248984 320126
rect 248932 320062 248984 320068
rect 248840 319712 248892 319718
rect 248840 319654 248892 319660
rect 248944 316810 248972 320062
rect 246460 316782 246796 316810
rect 247288 316782 247716 316810
rect 248636 316782 248972 316810
rect 249128 316810 249156 320470
rect 250048 316810 250076 326998
rect 252888 326648 252940 326654
rect 252888 326590 252940 326596
rect 250956 320664 251008 320670
rect 250956 320606 251008 320612
rect 250968 316810 250996 320606
rect 252796 319984 252848 319990
rect 252796 319926 252848 319932
rect 251784 319712 251836 319718
rect 251784 319654 251836 319660
rect 251796 316810 251824 319654
rect 252808 316810 252836 319926
rect 252900 316946 252928 326590
rect 258316 326580 258368 326586
rect 258316 326522 258368 326528
rect 254084 326512 254136 326518
rect 254084 326454 254136 326460
rect 253532 326444 253584 326450
rect 253532 326386 253584 326392
rect 253544 319582 253572 326386
rect 253532 319576 253584 319582
rect 253532 319518 253584 319524
rect 254096 319394 254124 326454
rect 254544 326308 254596 326314
rect 254544 326250 254596 326256
rect 254556 320194 254584 326250
rect 257120 320324 257172 320330
rect 257120 320266 257172 320272
rect 254544 320188 254596 320194
rect 254544 320130 254596 320136
rect 255556 320052 255608 320058
rect 255556 319994 255608 320000
rect 254096 319366 254400 319394
rect 252900 316918 253296 316946
rect 253268 316810 253296 316918
rect 254372 316810 254400 319366
rect 255568 316810 255596 319994
rect 256292 319576 256344 319582
rect 256292 319518 256344 319524
rect 256304 316810 256332 319518
rect 257132 316810 257160 320266
rect 258328 317082 258356 326522
rect 258328 317054 258402 317082
rect 249128 316782 249464 316810
rect 250048 316782 250384 316810
rect 250968 316782 251304 316810
rect 251796 316782 252132 316810
rect 252808 316782 253052 316810
rect 253268 316782 253972 316810
rect 254372 316782 254800 316810
rect 255568 316782 255720 316810
rect 256304 316782 256640 316810
rect 257132 316782 257468 316810
rect 258374 316796 258402 317054
rect 258972 313122 259000 327134
rect 259248 326314 259276 329838
rect 260168 326858 260196 329838
rect 260156 326852 260208 326858
rect 260156 326794 260208 326800
rect 261180 326790 261208 329838
rect 261168 326784 261220 326790
rect 261168 326726 261220 326732
rect 262100 326654 262128 329838
rect 263112 326722 263140 329838
rect 264124 327062 264152 329838
rect 264112 327056 264164 327062
rect 264112 326998 264164 327004
rect 263100 326716 263152 326722
rect 263100 326658 263152 326664
rect 259696 326648 259748 326654
rect 259696 326590 259748 326596
rect 262088 326648 262140 326654
rect 262088 326590 262140 326596
rect 259236 326308 259288 326314
rect 259236 326250 259288 326256
rect 259708 320126 259736 326590
rect 259696 320120 259748 320126
rect 259696 320062 259748 320068
rect 258960 313116 259012 313122
rect 258960 313058 259012 313064
rect 240650 310160 240706 310169
rect 240650 310095 240706 310104
rect 240664 309722 240692 310095
rect 240652 309716 240704 309722
rect 240652 309658 240704 309664
rect 240926 296832 240982 296841
rect 240926 296767 240982 296776
rect 240940 295918 240968 296767
rect 240928 295912 240980 295918
rect 240928 295854 240980 295860
rect 240376 283536 240428 283542
rect 240374 283504 240376 283513
rect 240428 283504 240430 283513
rect 240374 283439 240430 283448
rect 236236 283060 236288 283066
rect 236236 283002 236288 283008
rect 236880 283060 236932 283066
rect 236880 283002 236932 283008
rect 236248 282794 236276 283002
rect 236236 282788 236288 282794
rect 236236 282730 236288 282736
rect 234120 275104 234172 275110
rect 234120 275046 234172 275052
rect 232738 274392 232794 274401
rect 232738 274327 232794 274336
rect 234132 273886 234160 275046
rect 234120 273880 234172 273886
rect 234120 273822 234172 273828
rect 234764 273880 234816 273886
rect 234764 273822 234816 273828
rect 231634 273440 231690 273449
rect 231634 273375 231690 273384
rect 233474 263104 233530 263113
rect 233474 263039 233530 263048
rect 233488 262938 233516 263039
rect 233476 262932 233528 262938
rect 233476 262874 233528 262880
rect 233474 261744 233530 261753
rect 233474 261679 233530 261688
rect 233488 261442 233516 261679
rect 233476 261436 233528 261442
rect 233476 261378 233528 261384
rect 233474 260384 233530 260393
rect 233474 260319 233530 260328
rect 233488 260082 233516 260319
rect 233476 260076 233528 260082
rect 233476 260018 233528 260024
rect 233474 258888 233530 258897
rect 233474 258823 233530 258832
rect 233488 258654 233516 258823
rect 233476 258648 233528 258654
rect 233476 258590 233528 258596
rect 233474 257528 233530 257537
rect 233474 257463 233530 257472
rect 232832 257356 232884 257362
rect 232832 257298 232884 257304
rect 232738 254672 232794 254681
rect 232738 254607 232794 254616
rect 232752 244782 232780 254607
rect 232844 249785 232872 257298
rect 233488 257294 233516 257463
rect 233476 257288 233528 257294
rect 233476 257230 233528 257236
rect 233474 256168 233530 256177
rect 233474 256103 233530 256112
rect 233488 255934 233516 256103
rect 233476 255928 233528 255934
rect 233476 255870 233528 255876
rect 234580 255180 234632 255186
rect 234580 255122 234632 255128
rect 234212 253412 234264 253418
rect 234212 253354 234264 253360
rect 233474 253312 233530 253321
rect 233474 253247 233530 253256
rect 233488 253214 233516 253247
rect 233476 253208 233528 253214
rect 233476 253150 233528 253156
rect 233566 251952 233622 251961
rect 233566 251887 233622 251896
rect 233580 251786 233608 251887
rect 233568 251780 233620 251786
rect 233568 251722 233620 251728
rect 233476 251032 233528 251038
rect 233474 251000 233476 251009
rect 233528 251000 233530 251009
rect 233474 250935 233530 250944
rect 232830 249776 232886 249785
rect 232830 249711 232886 249720
rect 234120 248992 234172 248998
rect 234120 248934 234172 248940
rect 233476 248924 233528 248930
rect 233476 248866 233528 248872
rect 233488 248425 233516 248866
rect 233474 248416 233530 248425
rect 233474 248351 233530 248360
rect 233476 246204 233528 246210
rect 233476 246146 233528 246152
rect 233488 245569 233516 246146
rect 233474 245560 233530 245569
rect 233474 245495 233530 245504
rect 232740 244776 232792 244782
rect 232740 244718 232792 244724
rect 233476 243280 233528 243286
rect 233476 243222 233528 243228
rect 233488 242849 233516 243222
rect 233474 242840 233530 242849
rect 233474 242775 233530 242784
rect 233474 240664 233530 240673
rect 233474 240599 233476 240608
rect 233528 240599 233530 240608
rect 233476 240570 233528 240576
rect 233474 239304 233530 239313
rect 233474 239239 233476 239248
rect 233528 239239 233530 239248
rect 233476 239210 233528 239216
rect 234132 238633 234160 248934
rect 234224 244209 234252 253354
rect 234592 246929 234620 255122
rect 234578 246920 234634 246929
rect 234578 246855 234634 246864
rect 234210 244200 234266 244209
rect 234210 244135 234266 244144
rect 234118 238624 234174 238633
rect 234118 238559 234174 238568
rect 233476 237228 233528 237234
rect 233476 237170 233528 237176
rect 233488 237137 233516 237170
rect 233474 237128 233530 237137
rect 233474 237063 233530 237072
rect 234776 233766 234804 273822
rect 236892 266406 236920 283002
rect 243208 276934 243544 276962
rect 243760 276934 244096 276962
rect 244404 276934 244464 276962
rect 245048 276934 245384 276962
rect 245600 276934 245752 276962
rect 246244 276934 246580 276962
rect 246888 276934 247132 276962
rect 247440 276934 247776 276962
rect 248084 276934 248604 276962
rect 248728 276934 249064 276962
rect 243516 274906 243544 276934
rect 243504 274900 243556 274906
rect 243504 274842 243556 274848
rect 244068 274838 244096 276934
rect 244056 274832 244108 274838
rect 244056 274774 244108 274780
rect 243044 274764 243096 274770
rect 243044 274706 243096 274712
rect 241664 274696 241716 274702
rect 241664 274638 241716 274644
rect 240284 274628 240336 274634
rect 240284 274570 240336 274576
rect 238904 274560 238956 274566
rect 238904 274502 238956 274508
rect 237524 274492 237576 274498
rect 237524 274434 237576 274440
rect 236880 266400 236932 266406
rect 236880 266342 236932 266348
rect 237536 263770 237564 274434
rect 238916 263770 238944 274502
rect 240296 263770 240324 274570
rect 241676 263770 241704 274638
rect 243056 263770 243084 274706
rect 244436 266610 244464 276934
rect 245356 273818 245384 276934
rect 245344 273812 245396 273818
rect 245344 273754 245396 273760
rect 244884 266740 244936 266746
rect 244884 266682 244936 266688
rect 244424 266604 244476 266610
rect 244424 266546 244476 266552
rect 244896 263770 244924 266682
rect 245724 266474 245752 276934
rect 246552 274294 246580 276934
rect 246540 274288 246592 274294
rect 246540 274230 246592 274236
rect 245804 273812 245856 273818
rect 245804 273754 245856 273760
rect 245816 266678 245844 273754
rect 246264 266808 246316 266814
rect 246264 266750 246316 266756
rect 245804 266672 245856 266678
rect 245804 266614 245856 266620
rect 245712 266468 245764 266474
rect 245712 266410 245764 266416
rect 246276 263770 246304 266750
rect 247104 266270 247132 276934
rect 247274 274392 247330 274401
rect 247274 274327 247330 274336
rect 247184 274288 247236 274294
rect 247184 274230 247236 274236
rect 247196 266542 247224 274230
rect 247288 274022 247316 274327
rect 247276 274016 247328 274022
rect 247276 273958 247328 273964
rect 247748 273818 247776 276934
rect 247828 274016 247880 274022
rect 247826 273984 247828 273993
rect 247880 273984 247882 273993
rect 247826 273919 247882 273928
rect 247736 273812 247788 273818
rect 247736 273754 247788 273760
rect 248472 273812 248524 273818
rect 248472 273754 248524 273760
rect 247644 266876 247696 266882
rect 247644 266818 247696 266824
rect 247184 266536 247236 266542
rect 247184 266478 247236 266484
rect 247092 266264 247144 266270
rect 247092 266206 247144 266212
rect 247656 263770 247684 266818
rect 248484 266338 248512 273754
rect 248472 266332 248524 266338
rect 248472 266274 248524 266280
rect 248576 266202 248604 276934
rect 249036 273818 249064 276934
rect 249128 276934 249280 276962
rect 249588 276934 249924 276962
rect 250568 276934 250904 276962
rect 249128 275110 249156 276934
rect 249116 275104 249168 275110
rect 249116 275046 249168 275052
rect 249588 274022 249616 276934
rect 250876 274401 250904 276934
rect 250968 276934 251212 276962
rect 251764 276934 252100 276962
rect 252408 276934 252744 276962
rect 253052 276934 253204 276962
rect 250862 274392 250918 274401
rect 250862 274327 250918 274336
rect 249576 274016 249628 274022
rect 249576 273958 249628 273964
rect 250968 273857 250996 276934
rect 252072 274537 252100 276934
rect 252716 274673 252744 276934
rect 252980 274900 253032 274906
rect 252980 274842 253032 274848
rect 252702 274664 252758 274673
rect 252702 274599 252758 274608
rect 252058 274528 252114 274537
rect 252058 274463 252114 274472
rect 250954 273848 251010 273857
rect 249024 273812 249076 273818
rect 249024 273754 249076 273760
rect 249944 273812 249996 273818
rect 250954 273783 251010 273792
rect 249944 273754 249996 273760
rect 248564 266196 248616 266202
rect 248564 266138 248616 266144
rect 249024 265584 249076 265590
rect 249024 265526 249076 265532
rect 249036 263770 249064 265526
rect 237536 263742 237596 263770
rect 238916 263742 238976 263770
rect 240296 263742 240356 263770
rect 241676 263742 241736 263770
rect 243056 263742 243116 263770
rect 244588 263742 244924 263770
rect 245968 263742 246304 263770
rect 247348 263742 247684 263770
rect 248728 263742 249064 263770
rect 249956 263482 249984 273754
rect 250036 266400 250088 266406
rect 250036 266342 250088 266348
rect 250048 263770 250076 266342
rect 251876 265720 251928 265726
rect 251876 265662 251928 265668
rect 251888 263770 251916 265662
rect 252992 264042 253020 274842
rect 253176 274809 253204 276934
rect 253268 276934 253604 276962
rect 253162 274800 253218 274809
rect 253162 274735 253218 274744
rect 253268 274498 253296 276934
rect 254234 276690 254262 276948
rect 254188 276662 254262 276690
rect 254556 276934 254892 276962
rect 255108 276934 255444 276962
rect 255752 276934 256088 276962
rect 256212 276934 256732 276962
rect 256948 276934 257284 276962
rect 257592 276934 257928 276962
rect 258328 276934 258572 276962
rect 254188 274566 254216 276662
rect 254452 274832 254504 274838
rect 254452 274774 254504 274780
rect 254176 274560 254228 274566
rect 254176 274502 254228 274508
rect 253256 274492 253308 274498
rect 253256 274434 253308 274440
rect 250048 263742 250108 263770
rect 251580 263742 251916 263770
rect 252946 264014 253020 264042
rect 252946 263756 252974 264014
rect 254464 263770 254492 274774
rect 254556 274634 254584 276934
rect 255108 274702 255136 276934
rect 255752 274770 255780 276934
rect 255740 274764 255792 274770
rect 255740 274706 255792 274712
rect 255096 274696 255148 274702
rect 255096 274638 255148 274644
rect 254544 274628 254596 274634
rect 254544 274570 254596 274576
rect 256212 273970 256240 276934
rect 254820 273948 254872 273954
rect 254820 273890 254872 273896
rect 255660 273942 256240 273970
rect 254832 266882 254860 273890
rect 254820 266876 254872 266882
rect 254820 266818 254872 266824
rect 255660 266746 255688 273942
rect 256200 273880 256252 273886
rect 256200 273822 256252 273828
rect 255648 266740 255700 266746
rect 255648 266682 255700 266688
rect 255556 266604 255608 266610
rect 255556 266546 255608 266552
rect 254340 263742 254492 263770
rect 255568 263770 255596 266546
rect 256212 265590 256240 273822
rect 256948 273818 256976 276934
rect 257592 273954 257620 276934
rect 257580 273948 257632 273954
rect 257580 273890 257632 273896
rect 258328 273886 258356 276934
rect 258316 273880 258368 273886
rect 258316 273822 258368 273828
rect 256292 273812 256344 273818
rect 256292 273754 256344 273760
rect 256936 273812 256988 273818
rect 256936 273754 256988 273760
rect 256304 266814 256332 273754
rect 256292 266808 256344 266814
rect 256292 266750 256344 266756
rect 256936 266672 256988 266678
rect 256936 266614 256988 266620
rect 256200 265584 256252 265590
rect 256200 265526 256252 265532
rect 256948 263770 256976 266614
rect 258408 266468 258460 266474
rect 258408 266410 258460 266416
rect 258420 263770 258448 266410
rect 258972 265726 259000 313058
rect 261718 306216 261774 306225
rect 261718 306151 261774 306160
rect 261732 297210 261760 306151
rect 261720 297204 261772 297210
rect 261720 297146 261772 297152
rect 261258 286360 261314 286369
rect 261258 286295 261260 286304
rect 261312 286295 261314 286304
rect 261260 286266 261312 286272
rect 259696 266536 259748 266542
rect 259696 266478 259748 266484
rect 258960 265720 259012 265726
rect 258960 265662 259012 265668
rect 259708 263770 259736 266478
rect 262456 266332 262508 266338
rect 262456 266274 262508 266280
rect 261076 266264 261128 266270
rect 261076 266206 261128 266212
rect 261088 263770 261116 266206
rect 262468 263770 262496 266274
rect 263836 266196 263888 266202
rect 263836 266138 263888 266144
rect 263848 263770 263876 266138
rect 255568 263742 255720 263770
rect 256948 263742 257100 263770
rect 258420 263742 258572 263770
rect 259708 263742 259952 263770
rect 261088 263742 261332 263770
rect 262468 263742 262712 263770
rect 263848 263742 264092 263770
rect 249944 263476 249996 263482
rect 249944 263418 249996 263424
rect 262640 236208 262692 236214
rect 244238 236176 244294 236185
rect 244128 236134 244238 236162
rect 262640 236150 262692 236156
rect 244238 236111 244294 236120
rect 244988 235998 245048 236026
rect 242490 235904 242546 235913
rect 236248 235862 237412 235890
rect 238332 235862 238668 235890
rect 239252 235862 239588 235890
rect 234764 233760 234816 233766
rect 234764 233702 234816 233708
rect 234776 233358 234804 233702
rect 231452 233352 231504 233358
rect 231452 233294 231504 233300
rect 234764 233352 234816 233358
rect 234764 233294 234816 233300
rect 231360 226212 231412 226218
rect 231360 226154 231412 226160
rect 231360 215876 231412 215882
rect 231360 215818 231412 215824
rect 230898 194968 230954 194977
rect 230898 194903 230954 194912
rect 231082 194968 231138 194977
rect 231082 194903 231138 194912
rect 230806 107928 230862 107937
rect 230806 107863 230862 107872
rect 230714 104392 230770 104401
rect 230714 104327 230770 104336
rect 230912 100049 230940 194903
rect 231372 185729 231400 215818
rect 231464 207761 231492 233294
rect 231728 233284 231780 233290
rect 231728 233226 231780 233232
rect 231636 233216 231688 233222
rect 231636 233158 231688 233164
rect 231542 216592 231598 216601
rect 231542 216527 231598 216536
rect 231450 207752 231506 207761
rect 231450 207687 231506 207696
rect 231452 202072 231504 202078
rect 231452 202014 231504 202020
rect 231358 185720 231414 185729
rect 231358 185655 231414 185664
rect 231464 182601 231492 202014
rect 231556 191985 231584 216527
rect 231648 210753 231676 233158
rect 231740 213881 231768 233226
rect 231726 213872 231782 213881
rect 231726 213807 231782 213816
rect 231634 210744 231690 210753
rect 231634 210679 231690 210688
rect 231634 204352 231690 204361
rect 231634 204287 231690 204296
rect 231648 204118 231676 204287
rect 231636 204112 231688 204118
rect 231636 204054 231688 204060
rect 231542 191976 231598 191985
rect 231542 191911 231598 191920
rect 232002 188848 232058 188857
rect 236248 188818 236276 235862
rect 238640 233154 238668 235862
rect 238628 233148 238680 233154
rect 238628 233090 238680 233096
rect 239560 226286 239588 235862
rect 239928 235862 240264 235890
rect 241184 235862 241520 235890
rect 239928 232513 239956 235862
rect 241492 233766 241520 235862
rect 242136 235862 242490 235890
rect 241480 233760 241532 233766
rect 241480 233702 241532 233708
rect 241492 233465 241520 233702
rect 241478 233456 241534 233465
rect 241478 233391 241534 233400
rect 242136 233222 242164 235862
rect 242490 235839 242546 235848
rect 243056 235862 243116 235890
rect 243056 233737 243084 235862
rect 244988 235194 245016 235998
rect 246046 235641 246074 235876
rect 246644 235862 246980 235890
rect 247992 235862 248328 235890
rect 248912 235862 249248 235890
rect 246032 235632 246088 235641
rect 246032 235567 246088 235576
rect 244976 235188 245028 235194
rect 244976 235130 245028 235136
rect 246644 234961 246672 235862
rect 246630 234952 246686 234961
rect 246630 234887 246686 234896
rect 246264 233760 246316 233766
rect 243042 233728 243098 233737
rect 246264 233702 246316 233708
rect 243042 233663 243098 233672
rect 243056 233290 243084 233663
rect 243596 233624 243648 233630
rect 243596 233566 243648 233572
rect 243044 233284 243096 233290
rect 243044 233226 243096 233232
rect 242124 233216 242176 233222
rect 242124 233158 242176 233164
rect 239914 232504 239970 232513
rect 239914 232439 239970 232448
rect 239548 226280 239600 226286
rect 239548 226222 239600 226228
rect 243608 222834 243636 233566
rect 245344 233284 245396 233290
rect 245344 233226 245396 233232
rect 244332 233216 244384 233222
rect 244332 233158 244384 233164
rect 244344 222834 244372 233158
rect 245356 222834 245384 233226
rect 246276 222834 246304 233702
rect 246644 233329 246672 234887
rect 248012 233556 248064 233562
rect 248012 233498 248064 233504
rect 246630 233320 246686 233329
rect 246630 233255 246686 233264
rect 247092 232944 247144 232950
rect 247092 232886 247144 232892
rect 247104 222834 247132 232886
rect 248024 222834 248052 233498
rect 248300 232474 248328 235862
rect 248932 233692 248984 233698
rect 248932 233634 248984 233640
rect 248288 232468 248340 232474
rect 248288 232410 248340 232416
rect 248944 222834 248972 233634
rect 249220 225266 249248 235862
rect 249772 235862 249924 235890
rect 250844 235862 251364 235890
rect 251856 235862 252192 235890
rect 249208 225260 249260 225266
rect 249208 225202 249260 225208
rect 249772 225198 249800 235862
rect 249944 233488 249996 233494
rect 249944 233430 249996 233436
rect 249760 225192 249812 225198
rect 249760 225134 249812 225140
rect 249956 222834 249984 233430
rect 250680 233352 250732 233358
rect 250680 233294 250732 233300
rect 250692 222834 250720 233294
rect 250772 232468 250824 232474
rect 250772 232410 250824 232416
rect 243300 222806 243636 222834
rect 244128 222806 244372 222834
rect 245048 222806 245384 222834
rect 245968 222806 246304 222834
rect 246796 222806 247132 222834
rect 247716 222806 248052 222834
rect 248636 222806 248972 222834
rect 249464 222806 249984 222834
rect 250384 222806 250720 222834
rect 250784 222562 250812 232410
rect 251336 225470 251364 235862
rect 252164 232474 252192 235862
rect 252716 235862 252776 235890
rect 253788 235862 254124 235890
rect 254708 235862 255044 235890
rect 255720 235862 256056 235890
rect 252716 232610 252744 235862
rect 252704 232604 252756 232610
rect 252704 232546 252756 232552
rect 254096 232542 254124 235862
rect 254084 232536 254136 232542
rect 254084 232478 254136 232484
rect 255016 232474 255044 235862
rect 256028 232678 256056 235862
rect 256304 235862 256640 235890
rect 257316 235862 257652 235890
rect 258420 235862 258572 235890
rect 259248 235862 259584 235890
rect 260168 235862 260504 235890
rect 261180 235862 261516 235890
rect 262100 235862 262436 235890
rect 256304 233630 256332 235862
rect 256292 233624 256344 233630
rect 256292 233566 256344 233572
rect 257316 233222 257344 235862
rect 258420 233290 258448 235862
rect 259248 233766 259276 235862
rect 259236 233760 259288 233766
rect 259236 233702 259288 233708
rect 258408 233284 258460 233290
rect 258408 233226 258460 233232
rect 257304 233216 257356 233222
rect 257304 233158 257356 233164
rect 260168 232950 260196 235862
rect 261180 233562 261208 235862
rect 262100 233698 262128 235862
rect 262546 235768 262602 235777
rect 262652 235754 262680 236150
rect 262602 235726 262680 235754
rect 263112 235862 263448 235890
rect 264032 235862 264368 235890
rect 262546 235703 262602 235712
rect 262560 235194 262588 235703
rect 262548 235188 262600 235194
rect 262548 235130 262600 235136
rect 262088 233692 262140 233698
rect 262088 233634 262140 233640
rect 261168 233556 261220 233562
rect 261168 233498 261220 233504
rect 263112 233494 263140 235862
rect 263100 233488 263152 233494
rect 263100 233430 263152 233436
rect 264032 233358 264060 235862
rect 264020 233352 264072 233358
rect 264020 233294 264072 233300
rect 260156 232944 260208 232950
rect 260156 232886 260208 232892
rect 258960 232876 259012 232882
rect 258960 232818 259012 232824
rect 256016 232672 256068 232678
rect 256016 232614 256068 232620
rect 258316 232672 258368 232678
rect 258316 232614 258368 232620
rect 255556 232604 255608 232610
rect 255556 232546 255608 232552
rect 252152 232468 252204 232474
rect 252152 232410 252204 232416
rect 254176 232468 254228 232474
rect 254176 232410 254228 232416
rect 255004 232468 255056 232474
rect 255004 232410 255056 232416
rect 251324 225464 251376 225470
rect 251324 225406 251376 225412
rect 253992 225464 254044 225470
rect 253992 225406 254044 225412
rect 252152 225260 252204 225266
rect 252152 225202 252204 225208
rect 252164 222834 252192 225202
rect 253072 225192 253124 225198
rect 253072 225134 253124 225140
rect 253084 222834 253112 225134
rect 254004 222834 254032 225406
rect 252132 222806 252192 222834
rect 253052 222806 253112 222834
rect 253972 222806 254032 222834
rect 254188 222562 254216 232410
rect 255568 222698 255596 232546
rect 255648 232536 255700 232542
rect 255648 232478 255700 232484
rect 255660 222970 255688 232478
rect 256936 232468 256988 232474
rect 256936 232410 256988 232416
rect 255660 222942 256148 222970
rect 255568 222670 255720 222698
rect 256120 222562 256148 222942
rect 256948 222562 256976 232410
rect 258328 223106 258356 232614
rect 258328 223078 258402 223106
rect 258374 222820 258402 223078
rect 250784 222534 251304 222562
rect 254188 222534 254800 222562
rect 256120 222534 256640 222562
rect 256948 222534 257468 222562
rect 258972 219282 259000 232818
rect 258960 219276 259012 219282
rect 258960 219218 259012 219224
rect 240926 216184 240982 216193
rect 240926 216119 240982 216128
rect 240940 215882 240968 216119
rect 240928 215876 240980 215882
rect 240928 215818 240980 215824
rect 242214 207752 242270 207761
rect 242214 207687 242270 207696
rect 242228 204633 242256 207687
rect 242214 204624 242270 204633
rect 242214 204559 242270 204568
rect 237522 204352 237578 204361
rect 237522 204287 237578 204296
rect 237536 204118 237564 204287
rect 237524 204112 237576 204118
rect 237524 204054 237576 204060
rect 240374 202856 240430 202865
rect 240374 202791 240430 202800
rect 240388 202078 240416 202791
rect 240376 202072 240428 202078
rect 240376 202014 240428 202020
rect 242582 202040 242638 202049
rect 242582 201975 242638 201984
rect 242596 192529 242624 201975
rect 242582 192520 242638 192529
rect 242582 192455 242638 192464
rect 240374 189528 240430 189537
rect 240374 189463 240430 189472
rect 232002 188783 232004 188792
rect 232056 188783 232058 188792
rect 236236 188812 236288 188818
rect 232004 188754 232056 188760
rect 236236 188754 236288 188760
rect 236880 188812 236932 188818
rect 236880 188754 236932 188760
rect 232740 188336 232792 188342
rect 232740 188278 232792 188284
rect 231450 182592 231506 182601
rect 231450 182527 231506 182536
rect 232752 179774 232780 188278
rect 230992 179768 231044 179774
rect 230992 179710 231044 179716
rect 232740 179768 232792 179774
rect 232740 179710 232792 179716
rect 231004 179473 231032 179710
rect 230990 179464 231046 179473
rect 230990 179399 231046 179408
rect 236892 172566 236920 188754
rect 240388 188342 240416 189463
rect 240376 188336 240428 188342
rect 240376 188278 240428 188284
rect 248930 183136 248986 183145
rect 248986 183094 249280 183122
rect 248930 183071 248986 183080
rect 243208 182822 243544 182850
rect 243760 182822 244096 182850
rect 244404 182822 244464 182850
rect 245048 182822 245384 182850
rect 243516 181066 243544 182822
rect 243504 181060 243556 181066
rect 243504 181002 243556 181008
rect 244068 180998 244096 182822
rect 244056 180992 244108 180998
rect 244056 180934 244108 180940
rect 243044 180924 243096 180930
rect 243044 180866 243096 180872
rect 240284 180856 240336 180862
rect 240284 180798 240336 180804
rect 238904 180720 238956 180726
rect 238904 180662 238956 180668
rect 237524 180652 237576 180658
rect 237524 180594 237576 180600
rect 236880 172560 236932 172566
rect 236880 172502 236932 172508
rect 237536 169794 237564 180594
rect 238916 169794 238944 180662
rect 240296 169794 240324 180798
rect 241664 180788 241716 180794
rect 241664 180730 241716 180736
rect 241676 169794 241704 180730
rect 243056 169794 243084 180866
rect 244436 172770 244464 182822
rect 245356 181338 245384 182822
rect 245540 182822 245600 182850
rect 246244 182822 246580 182850
rect 245344 181332 245396 181338
rect 245344 181274 245396 181280
rect 244884 172900 244936 172906
rect 244884 172842 244936 172848
rect 244424 172764 244476 172770
rect 244424 172706 244476 172712
rect 244896 169794 244924 172842
rect 245540 172294 245568 182822
rect 245804 181332 245856 181338
rect 245804 181274 245856 181280
rect 245816 172838 245844 181274
rect 246552 180386 246580 182822
rect 246828 182822 246888 182850
rect 247440 182822 247776 182850
rect 246540 180380 246592 180386
rect 246540 180322 246592 180328
rect 246264 172968 246316 172974
rect 246264 172910 246316 172916
rect 245804 172832 245856 172838
rect 245804 172774 245856 172780
rect 245528 172288 245580 172294
rect 245528 172230 245580 172236
rect 246276 169794 246304 172910
rect 246828 172634 246856 182822
rect 247748 180522 247776 182822
rect 248024 182822 248084 182850
rect 248728 182822 249064 182850
rect 247736 180516 247788 180522
rect 247736 180458 247788 180464
rect 247184 180380 247236 180386
rect 247184 180322 247236 180328
rect 247196 172702 247224 180322
rect 247184 172696 247236 172702
rect 247184 172638 247236 172644
rect 246816 172628 246868 172634
rect 246816 172570 246868 172576
rect 247644 172492 247696 172498
rect 247644 172434 247696 172440
rect 247656 169794 247684 172434
rect 248024 172362 248052 182822
rect 249036 182193 249064 182822
rect 249588 182822 249924 182850
rect 250232 182822 250568 182850
rect 251212 182822 251364 182850
rect 249022 182184 249078 182193
rect 249022 182119 249078 182128
rect 248564 180516 248616 180522
rect 248564 180458 248616 180464
rect 248576 172430 248604 180458
rect 249588 180017 249616 182822
rect 250232 180153 250260 182822
rect 251336 180561 251364 182822
rect 251428 182822 251764 182850
rect 252408 182822 252744 182850
rect 253052 182822 253388 182850
rect 251428 180697 251456 182822
rect 252060 181332 252112 181338
rect 252060 181274 252112 181280
rect 251414 180688 251470 180697
rect 251414 180623 251470 180632
rect 251322 180552 251378 180561
rect 251322 180487 251378 180496
rect 250218 180144 250274 180153
rect 250218 180079 250274 180088
rect 249574 180008 249630 180017
rect 249574 179943 249630 179952
rect 249024 173036 249076 173042
rect 249024 172978 249076 172984
rect 248564 172424 248616 172430
rect 248564 172366 248616 172372
rect 248012 172356 248064 172362
rect 248012 172298 248064 172304
rect 249036 169794 249064 172978
rect 250036 172560 250088 172566
rect 250036 172502 250088 172508
rect 237536 169766 237596 169794
rect 238916 169766 238976 169794
rect 240296 169766 240356 169794
rect 241676 169766 241736 169794
rect 243056 169766 243116 169794
rect 244588 169766 244924 169794
rect 245968 169766 246304 169794
rect 247348 169766 247684 169794
rect 248728 169766 249064 169794
rect 250048 169794 250076 172502
rect 252072 172498 252100 181274
rect 252716 180697 252744 182822
rect 252796 181060 252848 181066
rect 252796 181002 252848 181008
rect 252702 180688 252758 180697
rect 252702 180623 252758 180632
rect 252060 172492 252112 172498
rect 252060 172434 252112 172440
rect 251876 171744 251928 171750
rect 251876 171686 251928 171692
rect 251888 169794 251916 171686
rect 250048 169766 250108 169794
rect 251580 169766 251916 169794
rect 252808 169794 252836 181002
rect 253360 180833 253388 182822
rect 253452 182822 253604 182850
rect 254248 182822 254308 182850
rect 253346 180824 253402 180833
rect 253346 180759 253402 180768
rect 253452 180658 253480 182822
rect 254176 180992 254228 180998
rect 254176 180934 254228 180940
rect 253440 180652 253492 180658
rect 253440 180594 253492 180600
rect 254188 169794 254216 180934
rect 254280 180726 254308 182822
rect 254556 182822 254892 182850
rect 255108 182822 255444 182850
rect 255752 182822 256088 182850
rect 256732 182822 256792 182850
rect 257284 182822 257344 182850
rect 254556 180862 254584 182822
rect 254544 180856 254596 180862
rect 254544 180798 254596 180804
rect 255108 180794 255136 182822
rect 255752 180930 255780 182822
rect 255740 180924 255792 180930
rect 255740 180866 255792 180872
rect 255096 180788 255148 180794
rect 255096 180730 255148 180736
rect 254268 180720 254320 180726
rect 254268 180662 254320 180668
rect 254820 179972 254872 179978
rect 254820 179914 254872 179920
rect 254832 173042 254860 179914
rect 254820 173036 254872 173042
rect 254820 172978 254872 172984
rect 256764 172906 256792 182822
rect 257316 172974 257344 182822
rect 257592 182822 257928 182850
rect 258420 182822 258572 182850
rect 257592 181338 257620 182822
rect 257580 181332 257632 181338
rect 257580 181274 257632 181280
rect 258420 179978 258448 182822
rect 258408 179972 258460 179978
rect 258408 179914 258460 179920
rect 257304 172968 257356 172974
rect 257304 172910 257356 172916
rect 256752 172900 256804 172906
rect 256752 172842 256804 172848
rect 256936 172832 256988 172838
rect 256936 172774 256988 172780
rect 255556 172764 255608 172770
rect 255556 172706 255608 172712
rect 255568 169794 255596 172706
rect 256948 169794 256976 172774
rect 258316 172628 258368 172634
rect 258316 172570 258368 172576
rect 258328 169794 258356 172570
rect 258972 171750 259000 219218
rect 261718 212784 261774 212793
rect 261718 212719 261774 212728
rect 261732 203370 261760 212719
rect 261720 203364 261772 203370
rect 261720 203306 261772 203312
rect 262362 192792 262418 192801
rect 262362 192727 262418 192736
rect 262376 192422 262404 192727
rect 262364 192416 262416 192422
rect 262364 192358 262416 192364
rect 259696 172696 259748 172702
rect 259696 172638 259748 172644
rect 258960 171744 259012 171750
rect 258960 171686 259012 171692
rect 259708 169794 259736 172638
rect 262456 172492 262508 172498
rect 262456 172434 262508 172440
rect 261168 172424 261220 172430
rect 261168 172366 261220 172372
rect 261180 169794 261208 172366
rect 262468 169794 262496 172434
rect 263836 172356 263888 172362
rect 263836 172298 263888 172304
rect 263848 169794 263876 172298
rect 252808 169766 252960 169794
rect 254188 169766 254340 169794
rect 255568 169766 255720 169794
rect 256948 169766 257100 169794
rect 258328 169766 258572 169794
rect 259708 169766 259952 169794
rect 261180 169766 261332 169794
rect 262468 169766 262712 169794
rect 263848 169766 264092 169794
rect 233474 169128 233530 169137
rect 233474 169063 233530 169072
rect 233488 168962 233516 169063
rect 233476 168956 233528 168962
rect 233476 168898 233528 168904
rect 233474 167768 233530 167777
rect 233474 167703 233530 167712
rect 233488 167602 233516 167703
rect 233476 167596 233528 167602
rect 233476 167538 233528 167544
rect 236878 167088 236934 167097
rect 236878 167023 236934 167032
rect 233474 166408 233530 166417
rect 233474 166343 233530 166352
rect 233488 166242 233516 166343
rect 233476 166236 233528 166242
rect 233476 166178 233528 166184
rect 233474 164912 233530 164921
rect 233474 164847 233530 164856
rect 233488 164814 233516 164847
rect 233476 164808 233528 164814
rect 233476 164750 233528 164756
rect 233474 163552 233530 163561
rect 232832 163516 232884 163522
rect 233474 163487 233530 163496
rect 232832 163458 232884 163464
rect 230992 162428 231044 162434
rect 230992 162370 231044 162376
rect 231004 155090 231032 162370
rect 231360 160660 231412 160666
rect 231360 160602 231412 160608
rect 230992 155084 231044 155090
rect 230992 155026 231044 155032
rect 231372 150874 231400 160602
rect 232740 159368 232792 159374
rect 232740 159310 232792 159316
rect 231360 150868 231412 150874
rect 231360 150810 231412 150816
rect 232752 149553 232780 159310
rect 232844 155129 232872 163458
rect 233488 163454 233516 163487
rect 233476 163448 233528 163454
rect 233476 163390 233528 163396
rect 233474 162192 233530 162201
rect 233474 162127 233530 162136
rect 233488 162094 233516 162127
rect 233476 162088 233528 162094
rect 233476 162030 233528 162036
rect 232924 160796 232976 160802
rect 232924 160738 232976 160744
rect 232830 155120 232886 155129
rect 232830 155055 232886 155064
rect 232936 152409 232964 160738
rect 233474 160696 233530 160705
rect 233474 160631 233476 160640
rect 233528 160631 233530 160640
rect 233476 160602 233528 160608
rect 233474 159336 233530 159345
rect 233474 159271 233476 159280
rect 233528 159271 233530 159280
rect 233476 159242 233528 159248
rect 233474 157976 233530 157985
rect 233474 157911 233476 157920
rect 233528 157911 233530 157920
rect 233476 157882 233528 157888
rect 233476 157192 233528 157198
rect 233476 157134 233528 157140
rect 233488 156625 233516 157134
rect 233474 156616 233530 156625
rect 233474 156551 233530 156560
rect 234028 155084 234080 155090
rect 234028 155026 234080 155032
rect 234040 153769 234068 155026
rect 234026 153760 234082 153769
rect 234026 153695 234082 153704
rect 232922 152400 232978 152409
rect 232922 152335 232978 152344
rect 233476 150936 233528 150942
rect 233474 150904 233476 150913
rect 233528 150904 233530 150913
rect 233474 150839 233530 150848
rect 232738 149544 232794 149553
rect 232738 149479 232794 149488
rect 233476 148216 233528 148222
rect 233474 148184 233476 148193
rect 233528 148184 233530 148193
rect 233474 148119 233530 148128
rect 233476 146788 233528 146794
rect 233476 146730 233528 146736
rect 233488 146697 233516 146730
rect 233474 146688 233530 146697
rect 233474 146623 233530 146632
rect 233476 145428 233528 145434
rect 233476 145370 233528 145376
rect 233488 145337 233516 145370
rect 233474 145328 233530 145337
rect 233474 145263 233530 145272
rect 233476 144068 233528 144074
rect 233476 144010 233528 144016
rect 233488 143977 233516 144010
rect 233474 143968 233530 143977
rect 233474 143903 233530 143912
rect 231360 143456 231412 143462
rect 231360 143398 231412 143404
rect 231176 143388 231228 143394
rect 231176 143330 231228 143336
rect 231188 141286 231216 143330
rect 231372 141354 231400 143398
rect 236892 142238 236920 167023
rect 236880 142232 236932 142238
rect 236880 142174 236932 142180
rect 238996 142232 239048 142238
rect 238996 142174 239048 142180
rect 239916 142232 239968 142238
rect 261904 142232 261956 142238
rect 242030 142200 242086 142209
rect 239968 142180 240264 142186
rect 239916 142174 240264 142180
rect 233474 142064 233530 142073
rect 233474 141999 233476 142008
rect 233528 141999 233530 142008
rect 233476 141970 233528 141976
rect 236248 141886 237412 141914
rect 238332 141886 238668 141914
rect 231360 141348 231412 141354
rect 231360 141290 231412 141296
rect 231176 141280 231228 141286
rect 231176 141222 231228 141228
rect 231084 140600 231136 140606
rect 231084 140542 231136 140548
rect 230990 140024 231046 140033
rect 230990 139959 231046 139968
rect 231004 123305 231032 139959
rect 231096 130270 231124 140542
rect 231372 132961 231400 141290
rect 231452 141280 231504 141286
rect 231452 141222 231504 141228
rect 231464 139761 231492 141222
rect 231450 139752 231506 139761
rect 231450 139687 231506 139696
rect 231358 132952 231414 132961
rect 231358 132887 231414 132896
rect 231360 131284 231412 131290
rect 231360 131226 231412 131232
rect 231084 130264 231136 130270
rect 231084 130206 231136 130212
rect 231096 129833 231124 130206
rect 231082 129824 231138 129833
rect 231082 129759 231138 129768
rect 230990 123296 231046 123305
rect 230990 123231 231046 123240
rect 230898 100040 230954 100049
rect 230898 99975 230954 99984
rect 231372 98553 231400 131226
rect 231464 126025 231492 139687
rect 231450 126016 231506 126025
rect 231450 125951 231506 125960
rect 231452 122036 231504 122042
rect 231452 121978 231504 121984
rect 231358 98544 231414 98553
rect 231358 98479 231414 98488
rect 231464 92297 231492 121978
rect 232002 109968 232058 109977
rect 232002 109903 232058 109912
rect 232016 109598 232044 109903
rect 232004 109592 232056 109598
rect 232056 109552 232136 109580
rect 232004 109534 232056 109540
rect 231544 108232 231596 108238
rect 231544 108174 231596 108180
rect 231450 92288 231506 92297
rect 231450 92223 231506 92232
rect 231556 88897 231584 108174
rect 232004 95040 232056 95046
rect 232002 95008 232004 95017
rect 232056 95008 232058 95017
rect 232002 94943 232058 94952
rect 231542 88888 231598 88897
rect 231542 88823 231598 88832
rect 231084 85792 231136 85798
rect 231082 85760 231084 85769
rect 231136 85760 231138 85769
rect 231082 85695 231138 85704
rect 230164 72396 230216 72402
rect 230164 72338 230216 72344
rect 230176 69546 230204 72338
rect 230624 70968 230676 70974
rect 230624 70910 230676 70916
rect 230164 69540 230216 69546
rect 230164 69482 230216 69488
rect 230636 66690 230664 70910
rect 230624 66684 230676 66690
rect 230624 66626 230676 66632
rect 229428 64372 229480 64378
rect 229428 64314 229480 64320
rect 229440 61454 229468 64314
rect 230440 62672 230492 62678
rect 230440 62614 230492 62620
rect 229428 61448 229480 61454
rect 229428 61390 229480 61396
rect 230452 61250 230480 62614
rect 230532 61312 230584 61318
rect 230532 61254 230584 61260
rect 230440 61244 230492 61250
rect 230440 61186 230492 61192
rect 230544 59482 230572 61254
rect 230624 59952 230676 59958
rect 230624 59894 230676 59900
rect 230532 59476 230584 59482
rect 230532 59418 230584 59424
rect 230636 58530 230664 59894
rect 230624 58524 230676 58530
rect 230624 58466 230676 58472
rect 232108 51594 232136 109552
rect 236248 95046 236276 141886
rect 238640 139246 238668 141886
rect 238628 139240 238680 139246
rect 238628 139182 238680 139188
rect 239008 109598 239036 142174
rect 239928 142158 240264 142174
rect 261902 142200 261904 142209
rect 261956 142200 261958 142209
rect 242086 142158 242532 142186
rect 242030 142135 242086 142144
rect 239252 141886 239588 141914
rect 241184 141886 241520 141914
rect 239560 139858 239588 141886
rect 239548 139852 239600 139858
rect 239548 139794 239600 139800
rect 241492 139586 241520 141886
rect 241756 139784 241808 139790
rect 241754 139752 241756 139761
rect 241808 139752 241810 139761
rect 241754 139687 241810 139696
rect 241480 139580 241532 139586
rect 241480 139522 241532 139528
rect 242504 138838 242532 142158
rect 261902 142135 261958 142144
rect 243116 141886 243268 141914
rect 243240 141801 243268 141886
rect 244068 141886 244128 141914
rect 244988 141886 245048 141914
rect 246060 141886 246396 141914
rect 243226 141792 243282 141801
rect 243226 141727 243282 141736
rect 244068 139897 244096 141886
rect 244054 139888 244110 139897
rect 244054 139823 244110 139832
rect 244988 139790 245016 141886
rect 244976 139784 245028 139790
rect 246368 139761 246396 141886
rect 246920 141886 246980 141914
rect 247992 141886 248512 141914
rect 248912 141886 249248 141914
rect 246920 141354 246948 141886
rect 246908 141348 246960 141354
rect 246908 141290 246960 141296
rect 247092 139784 247144 139790
rect 244976 139726 245028 139732
rect 246354 139752 246410 139761
rect 244332 139716 244384 139722
rect 244332 139658 244384 139664
rect 242492 138832 242544 138838
rect 242492 138774 242544 138780
rect 244344 130746 244372 139658
rect 244424 139308 244476 139314
rect 244424 139250 244476 139256
rect 243596 130740 243648 130746
rect 243596 130682 243648 130688
rect 244332 130740 244384 130746
rect 244332 130682 244384 130688
rect 242030 129552 242086 129561
rect 242030 129487 242086 129496
rect 242044 124801 242072 129487
rect 243608 128722 243636 130682
rect 244436 128722 244464 139250
rect 244988 138906 245016 139726
rect 246410 139710 246488 139738
rect 247092 139726 247144 139732
rect 246354 139687 246410 139696
rect 245804 138968 245856 138974
rect 245804 138910 245856 138916
rect 244976 138900 245028 138906
rect 244976 138842 245028 138848
rect 245816 131630 245844 138910
rect 245344 131624 245396 131630
rect 245344 131566 245396 131572
rect 245804 131624 245856 131630
rect 245804 131566 245856 131572
rect 245356 128722 245384 131566
rect 246264 130468 246316 130474
rect 246264 130410 246316 130416
rect 246276 128722 246304 130410
rect 246460 130270 246488 139710
rect 247104 130474 247132 139726
rect 247184 139036 247236 139042
rect 247184 138978 247236 138984
rect 247092 130468 247144 130474
rect 247092 130410 247144 130416
rect 246448 130264 246500 130270
rect 246446 130232 246448 130241
rect 246500 130232 246502 130241
rect 246446 130167 246502 130176
rect 247196 128722 247224 138978
rect 248012 131624 248064 131630
rect 248012 131566 248064 131572
rect 248024 128722 248052 131566
rect 248484 131222 248512 141886
rect 249220 139654 249248 141886
rect 249864 141886 249924 141914
rect 250844 141886 251180 141914
rect 251856 141886 252192 141914
rect 249208 139648 249260 139654
rect 249208 139590 249260 139596
rect 249864 139586 249892 141886
rect 251152 139926 251180 141886
rect 251140 139920 251192 139926
rect 251140 139862 251192 139868
rect 252060 139648 252112 139654
rect 252060 139590 252112 139596
rect 249668 139580 249720 139586
rect 249668 139522 249720 139528
rect 249852 139580 249904 139586
rect 249852 139522 249904 139528
rect 248564 139104 248616 139110
rect 248564 139046 248616 139052
rect 248576 131630 248604 139046
rect 249116 138832 249168 138838
rect 249116 138774 249168 138780
rect 249128 135817 249156 138774
rect 249680 138401 249708 139522
rect 251324 139444 251376 139450
rect 251324 139386 251376 139392
rect 249944 139376 249996 139382
rect 249944 139318 249996 139324
rect 249852 139172 249904 139178
rect 249852 139114 249904 139120
rect 249666 138392 249722 138401
rect 249666 138327 249722 138336
rect 249114 135808 249170 135817
rect 249114 135743 249170 135752
rect 249128 134457 249156 135743
rect 249114 134448 249170 134457
rect 249114 134383 249170 134392
rect 248564 131624 248616 131630
rect 248564 131566 248616 131572
rect 248472 131216 248524 131222
rect 248472 131158 248524 131164
rect 249864 130474 249892 139114
rect 248932 130468 248984 130474
rect 248932 130410 248984 130416
rect 249852 130468 249904 130474
rect 249852 130410 249904 130416
rect 248944 128722 248972 130410
rect 249956 128722 249984 139318
rect 250956 131216 251008 131222
rect 250956 131158 251008 131164
rect 250680 130740 250732 130746
rect 250680 130682 250732 130688
rect 250692 128722 250720 130682
rect 243300 128694 243636 128722
rect 244128 128694 244464 128722
rect 245048 128694 245384 128722
rect 245968 128694 246304 128722
rect 246796 128694 247224 128722
rect 247716 128694 248052 128722
rect 248636 128694 248972 128722
rect 249464 128694 249984 128722
rect 250384 128694 250720 128722
rect 250968 128722 250996 131158
rect 251336 130746 251364 139386
rect 251324 130740 251376 130746
rect 251324 130682 251376 130688
rect 252072 128994 252100 139590
rect 252164 138702 252192 141886
rect 252716 141886 252776 141914
rect 253788 141886 253940 141914
rect 254708 141886 255044 141914
rect 255720 141886 256056 141914
rect 252244 138900 252296 138906
rect 252244 138842 252296 138848
rect 252152 138696 252204 138702
rect 252152 138638 252204 138644
rect 252256 138537 252284 138842
rect 252716 138634 252744 141886
rect 253072 139580 253124 139586
rect 253072 139522 253124 139528
rect 252704 138628 252756 138634
rect 252704 138570 252756 138576
rect 252242 138528 252298 138537
rect 252242 138463 252298 138472
rect 252072 128966 252146 128994
rect 250968 128694 251304 128722
rect 252118 128708 252146 128966
rect 253084 128722 253112 139522
rect 253912 138838 253940 141886
rect 253992 139920 254044 139926
rect 253992 139862 254044 139868
rect 253900 138832 253952 138838
rect 253900 138774 253952 138780
rect 254004 128722 254032 139862
rect 254176 138696 254228 138702
rect 254176 138638 254228 138644
rect 253052 128694 253112 128722
rect 253972 128694 254032 128722
rect 254188 128586 254216 138638
rect 255016 138634 255044 141886
rect 256028 138702 256056 141886
rect 256304 141886 256640 141914
rect 257316 141886 257652 141914
rect 258328 141886 258572 141914
rect 259248 141886 259584 141914
rect 260168 141886 260504 141914
rect 261272 141886 261516 141914
rect 256304 139722 256332 141886
rect 256292 139716 256344 139722
rect 256292 139658 256344 139664
rect 257316 139314 257344 141886
rect 258328 139382 258356 141886
rect 259248 139790 259276 141886
rect 259236 139784 259288 139790
rect 259236 139726 259288 139732
rect 260168 139450 260196 141886
rect 261272 139518 261300 141886
rect 261916 141354 261944 142135
rect 262100 141886 262436 141914
rect 263112 141886 263448 141914
rect 264124 141886 264368 141914
rect 261904 141348 261956 141354
rect 261904 141290 261956 141296
rect 261260 139512 261312 139518
rect 261260 139454 261312 139460
rect 260156 139444 260208 139450
rect 260156 139386 260208 139392
rect 258316 139376 258368 139382
rect 258316 139318 258368 139324
rect 257304 139308 257356 139314
rect 257304 139250 257356 139256
rect 262100 139178 262128 141886
rect 263112 139586 263140 141886
rect 264124 139654 264152 141886
rect 264112 139648 264164 139654
rect 264112 139590 264164 139596
rect 263100 139580 263152 139586
rect 263100 139522 263152 139528
rect 264480 139240 264532 139246
rect 264480 139182 264532 139188
rect 262088 139172 262140 139178
rect 262088 139114 262140 139120
rect 256660 138832 256712 138838
rect 256660 138774 256712 138780
rect 256016 138696 256068 138702
rect 256016 138638 256068 138644
rect 254820 138628 254872 138634
rect 254820 138570 254872 138576
rect 255004 138628 255056 138634
rect 255004 138570 255056 138576
rect 254832 130338 254860 138570
rect 254820 130332 254872 130338
rect 254820 130274 254872 130280
rect 255556 130332 255608 130338
rect 255556 130274 255608 130280
rect 255568 128722 255596 130274
rect 256672 128722 256700 138774
rect 258684 138696 258736 138702
rect 258684 138638 258736 138644
rect 257488 138628 257540 138634
rect 257488 138570 257540 138576
rect 257500 128722 257528 138570
rect 258696 128722 258724 138638
rect 258960 132304 259012 132310
rect 258960 132246 259012 132252
rect 255568 128694 255720 128722
rect 256640 128694 256700 128722
rect 257468 128694 257528 128722
rect 258388 128694 258724 128722
rect 254188 128558 254800 128586
rect 242030 124792 242086 124801
rect 242030 124727 242086 124736
rect 240374 122208 240430 122217
rect 240374 122143 240430 122152
rect 240388 122042 240416 122143
rect 240376 122036 240428 122042
rect 240376 121978 240428 121984
rect 240098 109832 240154 109841
rect 240098 109767 240154 109776
rect 240112 109598 240140 109767
rect 238996 109592 239048 109598
rect 238996 109534 239048 109540
rect 240100 109592 240152 109598
rect 240100 109534 240152 109540
rect 240834 108880 240890 108889
rect 240834 108815 240890 108824
rect 240848 108238 240876 108815
rect 240836 108232 240888 108238
rect 240836 108174 240888 108180
rect 242030 100720 242086 100729
rect 242030 100655 242086 100664
rect 242044 95833 242072 100655
rect 242030 95824 242086 95833
rect 242030 95759 242086 95768
rect 240374 95552 240430 95561
rect 240374 95487 240430 95496
rect 236236 95040 236288 95046
rect 236236 94982 236288 94988
rect 235500 94428 235552 94434
rect 235500 94370 235552 94376
rect 235512 85798 235540 94370
rect 235500 85792 235552 85798
rect 235500 85734 235552 85740
rect 236248 79406 236276 94982
rect 240388 94434 240416 95487
rect 240376 94428 240428 94434
rect 240376 94370 240428 94376
rect 248930 89160 248986 89169
rect 248986 89118 249616 89146
rect 248930 89095 248986 89104
rect 243208 88846 243544 88874
rect 243760 88846 244096 88874
rect 244404 88846 244464 88874
rect 245048 88846 245384 88874
rect 245600 88846 245844 88874
rect 246244 88846 246580 88874
rect 246888 88846 247224 88874
rect 247440 88846 247776 88874
rect 248084 88846 248512 88874
rect 248728 88846 249064 88874
rect 243044 87152 243096 87158
rect 243044 87094 243096 87100
rect 241664 87016 241716 87022
rect 241664 86958 241716 86964
rect 240284 86880 240336 86886
rect 240284 86822 240336 86828
rect 238904 86812 238956 86818
rect 238904 86754 238956 86760
rect 236236 79400 236288 79406
rect 236236 79342 236288 79348
rect 237248 79400 237300 79406
rect 237248 79342 237300 79348
rect 233476 76408 233528 76414
rect 233476 76350 233528 76356
rect 233488 75297 233516 76350
rect 237260 75818 237288 79342
rect 238916 75818 238944 86754
rect 240296 75818 240324 86822
rect 241676 75818 241704 86958
rect 243056 75818 243084 87094
rect 243516 86138 243544 88846
rect 244068 86954 244096 88846
rect 244436 87294 244464 88846
rect 244424 87288 244476 87294
rect 244424 87230 244476 87236
rect 244056 86948 244108 86954
rect 244056 86890 244108 86896
rect 245356 86206 245384 88846
rect 245344 86200 245396 86206
rect 245344 86142 245396 86148
rect 243504 86132 243556 86138
rect 243504 86074 243556 86080
rect 245160 86132 245212 86138
rect 245160 86074 245212 86080
rect 245172 79202 245200 86074
rect 245160 79196 245212 79202
rect 245160 79138 245212 79144
rect 244884 78992 244936 78998
rect 244884 78934 244936 78940
rect 244896 75818 244924 78934
rect 245816 78794 245844 88846
rect 246552 86138 246580 88846
rect 246540 86132 246592 86138
rect 246540 86074 246592 86080
rect 247092 86132 247144 86138
rect 247092 86074 247144 86080
rect 246264 78856 246316 78862
rect 246264 78798 246316 78804
rect 245804 78788 245856 78794
rect 245804 78730 245856 78736
rect 246276 75818 246304 78798
rect 247104 78726 247132 86074
rect 247092 78720 247144 78726
rect 247092 78662 247144 78668
rect 247196 78590 247224 88846
rect 247748 86138 247776 88846
rect 247736 86132 247788 86138
rect 247736 86074 247788 86080
rect 247644 78924 247696 78930
rect 247644 78866 247696 78872
rect 247184 78584 247236 78590
rect 247184 78526 247236 78532
rect 247656 75818 247684 78866
rect 248484 78522 248512 88846
rect 249036 87430 249064 88846
rect 249024 87424 249076 87430
rect 249024 87366 249076 87372
rect 249588 86177 249616 89118
rect 250218 89024 250274 89033
rect 250274 88982 250568 89010
rect 250218 88959 250274 88968
rect 249666 88888 249722 88897
rect 249722 88846 249924 88874
rect 251212 88846 251364 88874
rect 249666 88823 249722 88832
rect 251336 86721 251364 88846
rect 251750 88625 251778 88860
rect 252072 88846 252408 88874
rect 253052 88846 253388 88874
rect 251736 88616 251792 88625
rect 251736 88551 251792 88560
rect 251322 86712 251378 86721
rect 251322 86647 251378 86656
rect 252072 86313 252100 88846
rect 252980 86948 253032 86954
rect 252980 86890 253032 86896
rect 252058 86304 252114 86313
rect 252058 86239 252114 86248
rect 252152 86268 252204 86274
rect 252152 86210 252204 86216
rect 252060 86200 252112 86206
rect 249574 86168 249630 86177
rect 248564 86132 248616 86138
rect 252060 86142 252112 86148
rect 249574 86103 249630 86112
rect 248564 86074 248616 86080
rect 248576 78658 248604 86074
rect 252072 79202 252100 86142
rect 251416 79196 251468 79202
rect 251416 79138 251468 79144
rect 252060 79196 252112 79202
rect 252060 79138 252112 79144
rect 249024 79128 249076 79134
rect 249024 79070 249076 79076
rect 248564 78652 248616 78658
rect 248564 78594 248616 78600
rect 248472 78516 248524 78522
rect 248472 78458 248524 78464
rect 249036 75818 249064 79070
rect 250404 78380 250456 78386
rect 250404 78322 250456 78328
rect 250416 75818 250444 78322
rect 237260 75790 237596 75818
rect 238916 75790 238976 75818
rect 240296 75790 240356 75818
rect 241676 75790 241736 75818
rect 243056 75790 243116 75818
rect 244588 75790 244924 75818
rect 245968 75790 246304 75818
rect 247348 75790 247684 75818
rect 248728 75790 249064 75818
rect 250108 75790 250444 75818
rect 251428 75818 251456 79138
rect 252164 78998 252192 86210
rect 252152 78992 252204 78998
rect 252152 78934 252204 78940
rect 252992 76090 253020 86890
rect 253360 86857 253388 88846
rect 253452 88846 253604 88874
rect 254248 88846 254308 88874
rect 253346 86848 253402 86857
rect 253452 86818 253480 88846
rect 254176 87288 254228 87294
rect 254176 87230 254228 87236
rect 253346 86783 253402 86792
rect 253440 86812 253492 86818
rect 253440 86754 253492 86760
rect 252946 76062 253020 76090
rect 251428 75790 251580 75818
rect 252946 75804 252974 76062
rect 254188 75818 254216 87230
rect 254280 86886 254308 88846
rect 254556 88846 254892 88874
rect 255108 88846 255444 88874
rect 255752 88846 256088 88874
rect 256212 88846 256732 88874
rect 256948 88846 257284 88874
rect 257684 88846 257928 88874
rect 258420 88846 258572 88874
rect 254556 87022 254584 88846
rect 255108 87158 255136 88846
rect 255096 87152 255148 87158
rect 255096 87094 255148 87100
rect 254544 87016 254596 87022
rect 254544 86958 254596 86964
rect 254268 86880 254320 86886
rect 254268 86822 254320 86828
rect 255752 86274 255780 88846
rect 255740 86268 255792 86274
rect 255740 86210 255792 86216
rect 256212 86154 256240 88846
rect 255660 86126 256240 86154
rect 256948 86138 256976 88846
rect 257580 86540 257632 86546
rect 257580 86482 257632 86488
rect 256292 86132 256344 86138
rect 255556 79196 255608 79202
rect 255556 79138 255608 79144
rect 255568 75818 255596 79138
rect 255660 78862 255688 86126
rect 256292 86074 256344 86080
rect 256936 86132 256988 86138
rect 256936 86074 256988 86080
rect 256200 86064 256252 86070
rect 256200 86006 256252 86012
rect 256212 79134 256240 86006
rect 256200 79128 256252 79134
rect 256200 79070 256252 79076
rect 256304 78930 256332 86074
rect 256292 78924 256344 78930
rect 256292 78866 256344 78872
rect 255648 78856 255700 78862
rect 255648 78798 255700 78804
rect 256936 78788 256988 78794
rect 256936 78730 256988 78736
rect 256948 75818 256976 78730
rect 257592 78386 257620 86482
rect 257684 86206 257712 88846
rect 258420 86546 258448 88846
rect 258972 87430 259000 132246
rect 264492 125306 264520 139182
rect 263836 125300 263888 125306
rect 263836 125242 263888 125248
rect 264480 125300 264532 125306
rect 264480 125242 264532 125248
rect 262362 118808 262418 118817
rect 262362 118743 262418 118752
rect 262376 117962 262404 118743
rect 262364 117956 262416 117962
rect 262364 117898 262416 117904
rect 261166 98816 261222 98825
rect 261166 98751 261222 98760
rect 261180 98582 261208 98751
rect 261168 98576 261220 98582
rect 261168 98518 261220 98524
rect 258960 87424 259012 87430
rect 258960 87366 259012 87372
rect 258408 86540 258460 86546
rect 258408 86482 258460 86488
rect 257672 86200 257724 86206
rect 257672 86142 257724 86148
rect 258408 78720 258460 78726
rect 258408 78662 258460 78668
rect 257580 78380 257632 78386
rect 257580 78322 257632 78328
rect 258420 75818 258448 78662
rect 261076 78652 261128 78658
rect 261076 78594 261128 78600
rect 259696 78584 259748 78590
rect 259696 78526 259748 78532
rect 259708 75818 259736 78526
rect 261088 75818 261116 78594
rect 262456 78516 262508 78522
rect 262456 78458 262508 78464
rect 262468 75818 262496 78458
rect 263848 75818 263876 125242
rect 254188 75790 254340 75818
rect 255568 75790 255720 75818
rect 256948 75790 257100 75818
rect 258420 75790 258572 75818
rect 259708 75790 259952 75818
rect 261088 75790 261332 75818
rect 262468 75790 262712 75818
rect 263848 75790 264092 75818
rect 233474 75288 233530 75297
rect 233474 75223 233530 75232
rect 233474 73792 233530 73801
rect 233474 73727 233476 73736
rect 233528 73727 233530 73736
rect 233476 73698 233528 73704
rect 233474 72568 233530 72577
rect 233474 72503 233530 72512
rect 233488 72402 233516 72503
rect 233476 72396 233528 72402
rect 233476 72338 233528 72344
rect 233474 71480 233530 71489
rect 233474 71415 233530 71424
rect 233488 68186 233516 71415
rect 233566 71072 233622 71081
rect 233566 71007 233622 71016
rect 233580 70974 233608 71007
rect 233568 70968 233620 70974
rect 233568 70910 233620 70916
rect 233566 69576 233622 69585
rect 233566 69511 233622 69520
rect 233476 68180 233528 68186
rect 233476 68122 233528 68128
rect 233474 67264 233530 67273
rect 233474 67199 233530 67208
rect 233488 65398 233516 67199
rect 233580 66758 233608 69511
rect 233658 68352 233714 68361
rect 233658 68287 233714 68296
rect 233568 66752 233620 66758
rect 233568 66694 233620 66700
rect 233476 65392 233528 65398
rect 233476 65334 233528 65340
rect 233672 65330 233700 68287
rect 234210 66992 234266 67001
rect 234210 66927 234266 66936
rect 233660 65324 233712 65330
rect 233660 65266 233712 65272
rect 233474 64544 233530 64553
rect 233474 64479 233530 64488
rect 233488 64378 233516 64479
rect 233476 64372 233528 64378
rect 233476 64314 233528 64320
rect 234224 64038 234252 66927
rect 234394 65496 234450 65505
rect 234394 65431 234450 65440
rect 234212 64032 234264 64038
rect 234212 63974 234264 63980
rect 233474 63184 233530 63193
rect 233474 63119 233530 63128
rect 233488 62678 233516 63119
rect 233566 62776 233622 62785
rect 233566 62711 233622 62720
rect 233476 62672 233528 62678
rect 233476 62614 233528 62620
rect 233474 61416 233530 61425
rect 233474 61351 233530 61360
rect 233488 61318 233516 61351
rect 233476 61312 233528 61318
rect 233476 61254 233528 61260
rect 233474 60056 233530 60065
rect 233474 59991 233530 60000
rect 233488 59958 233516 59991
rect 233476 59952 233528 59958
rect 233476 59894 233528 59900
rect 233580 59890 233608 62711
rect 234408 62610 234436 65431
rect 234396 62604 234448 62610
rect 234396 62546 234448 62552
rect 233568 59884 233620 59890
rect 233568 59826 233620 59832
rect 233658 58968 233714 58977
rect 233658 58903 233714 58912
rect 233474 58696 233530 58705
rect 233474 58631 233530 58640
rect 233488 57034 233516 58631
rect 233566 57200 233622 57209
rect 233566 57135 233622 57144
rect 233476 57028 233528 57034
rect 233476 56970 233528 56976
rect 233474 56112 233530 56121
rect 233474 56047 233530 56056
rect 233488 55810 233516 56047
rect 233476 55804 233528 55810
rect 233476 55746 233528 55752
rect 233580 55742 233608 57135
rect 233672 57102 233700 58903
rect 233660 57096 233712 57102
rect 233660 57038 233712 57044
rect 233568 55736 233620 55742
rect 233568 55678 233620 55684
rect 233474 55296 233530 55305
rect 233474 55231 233530 55240
rect 233488 55062 233516 55231
rect 233476 55056 233528 55062
rect 233476 54998 233528 55004
rect 233474 54480 233530 54489
rect 233474 54415 233476 54424
rect 233528 54415 233530 54424
rect 233476 54386 233528 54392
rect 233476 53696 233528 53702
rect 233476 53638 233528 53644
rect 233488 53537 233516 53638
rect 233474 53528 233530 53537
rect 233474 53463 233530 53472
rect 233476 52948 233528 52954
rect 233476 52890 233528 52896
rect 233488 52449 233516 52890
rect 233474 52440 233530 52449
rect 233474 52375 233530 52384
rect 232096 51588 232148 51594
rect 232096 51530 232148 51536
rect 228692 51520 228744 51526
rect 228692 51462 228744 51468
rect 232108 48194 232136 51530
rect 233566 50808 233622 50817
rect 233566 50743 233622 50752
rect 233474 50400 233530 50409
rect 233580 50370 233608 50743
rect 233474 50335 233530 50344
rect 233568 50364 233620 50370
rect 233488 50302 233516 50335
rect 233568 50306 233620 50312
rect 233476 50296 233528 50302
rect 233476 50238 233528 50244
rect 233474 49040 233530 49049
rect 233474 48975 233530 48984
rect 233488 48942 233516 48975
rect 233476 48936 233528 48942
rect 233476 48878 233528 48884
rect 241124 48194 241460 48210
rect 232096 48188 232148 48194
rect 232096 48130 232148 48136
rect 238628 48188 238680 48194
rect 238628 48130 238680 48136
rect 241112 48188 241460 48194
rect 241164 48182 241460 48188
rect 241112 48130 241164 48136
rect 238640 48097 238668 48130
rect 238626 48088 238682 48097
rect 260430 48088 260486 48097
rect 238626 48023 238682 48032
rect 250508 48046 250996 48074
rect 260136 48046 260430 48074
rect 250508 47961 250536 48046
rect 250494 47952 250550 47961
rect 238424 47910 238668 47938
rect 244588 47910 244924 47938
rect 247716 47910 248052 47938
rect 233474 47816 233530 47825
rect 233474 47751 233530 47760
rect 233488 47514 233516 47751
rect 233476 47508 233528 47514
rect 233476 47450 233528 47456
rect 238640 45950 238668 47910
rect 244896 46057 244924 47910
rect 248024 47281 248052 47910
rect 250494 47887 250550 47896
rect 248010 47272 248066 47281
rect 248010 47207 248066 47216
rect 244882 46048 244938 46057
rect 244882 45983 244938 45992
rect 238628 45944 238680 45950
rect 238628 45886 238680 45892
rect 250968 45882 250996 48046
rect 260430 48023 260486 48032
rect 262822 48088 262878 48097
rect 262878 48046 263264 48074
rect 262822 48023 262878 48032
rect 257302 47952 257358 47961
rect 253880 47910 254032 47938
rect 257008 47910 257302 47938
rect 250956 45876 251008 45882
rect 250956 45818 251008 45824
rect 254004 45814 254032 47910
rect 257302 47887 257358 47896
rect 262546 46048 262602 46057
rect 262546 45983 262602 45992
rect 262560 45814 262588 45983
rect 262836 45921 262864 48023
rect 262822 45912 262878 45921
rect 262822 45847 262878 45856
rect 253992 45808 254044 45814
rect 253992 45750 254044 45756
rect 262548 45808 262600 45814
rect 262548 45750 262600 45756
rect 262836 45338 262864 45847
rect 263100 45808 263152 45814
rect 263100 45750 263152 45756
rect 262824 45332 262876 45338
rect 262824 45274 262876 45280
rect 263112 44794 263140 45750
rect 263100 44788 263152 44794
rect 263100 44730 263152 44736
rect 261076 16636 261128 16642
rect 261076 16578 261128 16584
rect 248196 16568 248248 16574
rect 248196 16510 248248 16516
rect 235316 16500 235368 16506
rect 235316 16442 235368 16448
rect 228600 12284 228652 12290
rect 228600 12226 228652 12232
rect 235328 9304 235356 16442
rect 248208 9304 248236 16510
rect 261088 9304 261116 16578
rect 265872 12358 265900 388470
rect 266700 382906 266728 392398
rect 283984 389276 284036 389282
rect 283984 389218 284036 389224
rect 279016 389072 279068 389078
rect 279016 389014 279068 389020
rect 279028 386714 279056 389014
rect 283996 386714 284024 389218
rect 288952 389140 289004 389146
rect 288952 389082 289004 389088
rect 288964 386714 288992 389082
rect 294196 389004 294248 389010
rect 294196 388946 294248 388952
rect 294208 386714 294236 388946
rect 299452 386714 299480 393230
rect 302120 393129 302148 396344
rect 319784 393809 319812 396344
rect 319770 393800 319826 393809
rect 319770 393735 319826 393744
rect 337540 393430 337568 396344
rect 355204 393838 355232 396344
rect 355192 393832 355244 393838
rect 355192 393774 355244 393780
rect 358596 393832 358648 393838
rect 358596 393774 358648 393780
rect 337528 393424 337580 393430
rect 337528 393366 337580 393372
rect 358504 393424 358556 393430
rect 358504 393366 358556 393372
rect 304592 393356 304644 393362
rect 304592 393298 304644 393304
rect 302106 393120 302162 393129
rect 302106 393055 302162 393064
rect 304604 386714 304632 393298
rect 314620 389752 314672 389758
rect 314620 389694 314672 389700
rect 309008 388392 309060 388398
rect 309008 388334 309060 388340
rect 279028 386686 279364 386714
rect 283996 386686 284332 386714
rect 288964 386686 289300 386714
rect 294208 386686 294360 386714
rect 299328 386686 299480 386714
rect 304296 386686 304632 386714
rect 309020 386714 309048 388334
rect 314632 386714 314660 389694
rect 315632 388460 315684 388466
rect 315632 388402 315684 388408
rect 309020 386686 309356 386714
rect 314324 386686 314660 386714
rect 266700 382878 266820 382906
rect 266792 373234 266820 382878
rect 315644 378554 315672 388402
rect 319126 384824 319182 384833
rect 319126 384759 319182 384768
rect 319034 382104 319090 382113
rect 319034 382039 319090 382048
rect 315816 378668 315868 378674
rect 315816 378610 315868 378616
rect 315828 378554 315856 378610
rect 315644 378526 315856 378554
rect 266596 373228 266648 373234
rect 266596 373170 266648 373176
rect 266780 373228 266832 373234
rect 266780 373170 266832 373176
rect 266608 373114 266636 373170
rect 266608 373086 266820 373114
rect 266792 363578 266820 373086
rect 278076 370910 278412 370938
rect 277544 368332 277596 368338
rect 277544 368274 277596 368280
rect 266596 363572 266648 363578
rect 266596 363514 266648 363520
rect 266780 363572 266832 363578
rect 266780 363514 266832 363520
rect 266608 356574 266636 363514
rect 267332 357928 267384 357934
rect 267332 357870 267384 357876
rect 267344 357225 267372 357870
rect 267330 357216 267386 357225
rect 267330 357151 267386 357160
rect 266596 356568 266648 356574
rect 266596 356510 266648 356516
rect 266780 356568 266832 356574
rect 266780 356510 266832 356516
rect 267884 356568 267936 356574
rect 267884 356510 267936 356516
rect 266792 355214 266820 356510
rect 267896 356137 267924 356510
rect 267882 356128 267938 356137
rect 267882 356063 267938 356072
rect 266780 355208 266832 355214
rect 266780 355150 266832 355156
rect 266872 355208 266924 355214
rect 267884 355208 267936 355214
rect 266872 355150 266924 355156
rect 267882 355176 267884 355185
rect 267936 355176 267938 355185
rect 266884 349450 266912 355150
rect 267424 355140 267476 355146
rect 267882 355111 267938 355120
rect 267424 355082 267476 355088
rect 267436 354097 267464 355082
rect 267422 354088 267478 354097
rect 267422 354023 267478 354032
rect 267884 353848 267936 353854
rect 267884 353790 267936 353796
rect 267896 353009 267924 353790
rect 267882 353000 267938 353009
rect 267882 352935 267938 352944
rect 267884 352420 267936 352426
rect 267884 352362 267936 352368
rect 267896 352057 267924 352362
rect 267882 352048 267938 352057
rect 267882 351983 267938 351992
rect 274782 351368 274838 351377
rect 274782 351303 274838 351312
rect 267516 351060 267568 351066
rect 267516 351002 267568 351008
rect 267528 349881 267556 351002
rect 267698 350960 267754 350969
rect 267698 350895 267754 350904
rect 267712 350386 267740 350895
rect 267700 350380 267752 350386
rect 267700 350322 267752 350328
rect 267514 349872 267570 349881
rect 267514 349807 267570 349816
rect 274796 349706 274824 351303
rect 277556 351066 277584 368274
rect 278384 367658 278412 370910
rect 280408 370910 280560 370938
rect 282984 370910 283044 370938
rect 285284 370910 285528 370938
rect 288012 370910 288624 370938
rect 280408 368338 280436 370910
rect 280396 368332 280448 368338
rect 280396 368274 280448 368280
rect 282984 367658 283012 370910
rect 278372 367652 278424 367658
rect 278372 367594 278424 367600
rect 279660 367652 279712 367658
rect 279660 367594 279712 367600
rect 282972 367652 283024 367658
rect 282972 367594 283024 367600
rect 283800 367652 283852 367658
rect 283800 367594 283852 367600
rect 279672 355078 279700 367594
rect 283812 355078 283840 367594
rect 285284 367289 285312 370910
rect 285270 367280 285326 367289
rect 285270 367215 285326 367224
rect 288596 355078 288624 370910
rect 290068 370910 290496 370938
rect 293072 370910 293408 370938
rect 279660 355072 279712 355078
rect 279660 355014 279712 355020
rect 280396 355072 280448 355078
rect 280396 355014 280448 355020
rect 283800 355072 283852 355078
rect 283800 355014 283852 355020
rect 285364 355072 285416 355078
rect 285364 355014 285416 355020
rect 288584 355072 288636 355078
rect 288584 355014 288636 355020
rect 280408 351748 280436 355014
rect 285376 351748 285404 355014
rect 290068 352426 290096 370910
rect 293380 367658 293408 370910
rect 294208 370910 295556 370938
rect 298040 370910 298284 370938
rect 293368 367652 293420 367658
rect 293368 367594 293420 367600
rect 290332 355072 290384 355078
rect 290332 355014 290384 355020
rect 290056 352420 290108 352426
rect 290056 352362 290108 352368
rect 290344 351748 290372 355014
rect 294208 353854 294236 370910
rect 298256 367658 298284 370910
rect 299820 370910 300524 370938
rect 303008 370910 303344 370938
rect 294288 367652 294340 367658
rect 294288 367594 294340 367600
rect 298244 367652 298296 367658
rect 298244 367594 298296 367600
rect 299716 367652 299768 367658
rect 299716 367594 299768 367600
rect 294196 353848 294248 353854
rect 294196 353790 294248 353796
rect 294300 351898 294328 367594
rect 294300 351870 294972 351898
rect 284994 351640 285050 351649
rect 294944 351626 294972 351870
rect 299728 351626 299756 367594
rect 299820 355146 299848 370910
rect 303316 367658 303344 370910
rect 305340 370910 305584 370938
rect 308068 370910 308404 370938
rect 303304 367652 303356 367658
rect 303304 367594 303356 367600
rect 305236 367652 305288 367658
rect 305236 367594 305288 367600
rect 299808 355140 299860 355146
rect 299808 355082 299860 355088
rect 305248 351762 305276 367594
rect 305340 355214 305368 370910
rect 308376 367658 308404 370910
rect 309388 370910 310552 370938
rect 313036 370910 313464 370938
rect 308364 367652 308416 367658
rect 308364 367594 308416 367600
rect 309284 367652 309336 367658
rect 309284 367594 309336 367600
rect 305328 355208 305380 355214
rect 305328 355150 305380 355156
rect 309296 355078 309324 367594
rect 309388 356574 309416 370910
rect 309376 356568 309428 356574
rect 309376 356510 309428 356516
rect 313436 355078 313464 370910
rect 314908 370910 315520 370938
rect 314908 357934 314936 370910
rect 314896 357928 314948 357934
rect 314896 357870 314948 357876
rect 309284 355072 309336 355078
rect 309284 355014 309336 355020
rect 310388 355072 310440 355078
rect 310388 355014 310440 355020
rect 313424 355072 313476 355078
rect 313424 355014 313476 355020
rect 315356 355072 315408 355078
rect 315356 355014 315408 355020
rect 305248 351734 305354 351762
rect 310400 351748 310428 355014
rect 315368 351748 315396 355014
rect 294944 351598 295418 351626
rect 299728 351598 300386 351626
rect 284994 351575 284996 351584
rect 285048 351575 285050 351584
rect 284996 351546 285048 351552
rect 277544 351060 277596 351066
rect 277544 351002 277596 351008
rect 274966 350416 275022 350425
rect 274966 350351 275022 350360
rect 267884 349700 267936 349706
rect 267884 349642 267936 349648
rect 274784 349700 274836 349706
rect 274784 349642 274836 349648
rect 266884 349422 267004 349450
rect 266976 344169 267004 349422
rect 267896 348929 267924 349642
rect 274874 349600 274930 349609
rect 274874 349535 274930 349544
rect 267882 348920 267938 348929
rect 267882 348855 267938 348864
rect 267884 348272 267936 348278
rect 267884 348214 267936 348220
rect 267896 347841 267924 348214
rect 267882 347832 267938 347841
rect 267882 347767 267938 347776
rect 274888 346918 274916 349535
rect 274980 348278 275008 350351
rect 275058 348648 275114 348657
rect 275058 348583 275114 348592
rect 274968 348272 275020 348278
rect 274968 348214 275020 348220
rect 267884 346912 267936 346918
rect 267882 346880 267884 346889
rect 274876 346912 274928 346918
rect 267936 346880 267938 346889
rect 267424 346844 267476 346850
rect 274876 346854 274928 346860
rect 274966 346880 275022 346889
rect 267882 346815 267938 346824
rect 275072 346850 275100 348583
rect 275150 347832 275206 347841
rect 275150 347767 275206 347776
rect 274966 346815 275022 346824
rect 275060 346844 275112 346850
rect 267424 346786 267476 346792
rect 267436 345801 267464 346786
rect 274874 346064 274930 346073
rect 274874 345999 274930 346008
rect 267422 345792 267478 345801
rect 267422 345727 267478 345736
rect 274888 345626 274916 345999
rect 270736 345620 270788 345626
rect 270736 345562 270788 345568
rect 274876 345620 274928 345626
rect 274876 345562 274928 345568
rect 267884 345552 267936 345558
rect 267884 345494 267936 345500
rect 267896 344713 267924 345494
rect 267882 344704 267938 344713
rect 267882 344639 267938 344648
rect 266962 344160 267018 344169
rect 266688 344124 266740 344130
rect 266962 344095 267018 344104
rect 267146 344160 267202 344169
rect 267146 344095 267202 344104
rect 266688 344066 266740 344072
rect 266700 343761 266728 344066
rect 266686 343752 266742 343761
rect 266686 343687 266742 343696
rect 267160 339370 267188 344095
rect 267608 342764 267660 342770
rect 267608 342706 267660 342712
rect 267620 341585 267648 342706
rect 270748 342702 270776 345562
rect 274874 345112 274930 345121
rect 274874 345047 274930 345056
rect 274888 342770 274916 345047
rect 274980 344130 275008 346815
rect 275060 346786 275112 346792
rect 275164 345558 275192 347767
rect 275152 345552 275204 345558
rect 275152 345494 275204 345500
rect 275058 344296 275114 344305
rect 275058 344231 275114 344240
rect 274968 344124 275020 344130
rect 274968 344066 275020 344072
rect 274876 342764 274928 342770
rect 274876 342706 274928 342712
rect 267884 342696 267936 342702
rect 267882 342664 267884 342673
rect 270736 342696 270788 342702
rect 267936 342664 267938 342673
rect 270736 342638 270788 342644
rect 267882 342599 267938 342608
rect 267606 341576 267662 341585
rect 267606 341511 267662 341520
rect 274966 341576 275022 341585
rect 274966 341511 275022 341520
rect 267884 341404 267936 341410
rect 267884 341346 267936 341352
rect 267896 340633 267924 341346
rect 267882 340624 267938 340633
rect 267882 340559 267938 340568
rect 274874 340624 274930 340633
rect 274874 340559 274930 340568
rect 274888 340118 274916 340559
rect 272024 340112 272076 340118
rect 272024 340054 272076 340060
rect 274876 340112 274928 340118
rect 274876 340054 274928 340060
rect 267884 340044 267936 340050
rect 267884 339986 267936 339992
rect 267896 339545 267924 339986
rect 267882 339536 267938 339545
rect 267882 339471 267938 339480
rect 267148 339364 267200 339370
rect 267148 339306 267200 339312
rect 267792 338684 267844 338690
rect 267792 338626 267844 338632
rect 267516 338616 267568 338622
rect 267516 338558 267568 338564
rect 267528 337505 267556 338558
rect 267514 337496 267570 337505
rect 267514 337431 267570 337440
rect 267332 337256 267384 337262
rect 267332 337198 267384 337204
rect 267344 336417 267372 337198
rect 267330 336408 267386 336417
rect 267330 336343 267386 336352
rect 266780 335964 266832 335970
rect 266780 335906 266832 335912
rect 266792 331249 266820 335906
rect 267332 334468 267384 334474
rect 267332 334410 267384 334416
rect 267344 333289 267372 334410
rect 267804 334377 267832 338626
rect 267882 338584 267938 338593
rect 267882 338519 267884 338528
rect 267936 338519 267938 338528
rect 267884 338490 267936 338496
rect 270828 337324 270880 337330
rect 270828 337266 270880 337272
rect 270736 336032 270788 336038
rect 270736 335974 270788 335980
rect 267884 335896 267936 335902
rect 267884 335838 267936 335844
rect 267896 335465 267924 335838
rect 267882 335456 267938 335465
rect 267882 335391 267938 335400
rect 267790 334368 267846 334377
rect 267790 334303 267846 334312
rect 267330 333280 267386 333289
rect 267330 333215 267386 333224
rect 270748 333114 270776 335974
rect 270840 334474 270868 337266
rect 272036 337262 272064 340054
rect 274874 338856 274930 338865
rect 274874 338791 274930 338800
rect 274888 338690 274916 338791
rect 274876 338684 274928 338690
rect 274876 338626 274928 338632
rect 274980 338622 275008 341511
rect 275072 341410 275100 344231
rect 275150 343344 275206 343353
rect 275150 343279 275206 343288
rect 275060 341404 275112 341410
rect 275060 341346 275112 341352
rect 275164 340050 275192 343279
rect 275242 342392 275298 342401
rect 275242 342327 275298 342336
rect 275152 340044 275204 340050
rect 275152 339986 275204 339992
rect 275058 339808 275114 339817
rect 275058 339743 275114 339752
rect 274968 338616 275020 338622
rect 274968 338558 275020 338564
rect 274874 338040 274930 338049
rect 274874 337975 274930 337984
rect 274888 337330 274916 337975
rect 274876 337324 274928 337330
rect 274876 337266 274928 337272
rect 272024 337256 272076 337262
rect 272024 337198 272076 337204
rect 274966 337088 275022 337097
rect 274966 337023 275022 337032
rect 274874 336272 274930 336281
rect 274874 336207 274930 336216
rect 274888 335970 274916 336207
rect 274980 336038 275008 337023
rect 274968 336032 275020 336038
rect 274968 335974 275020 335980
rect 274876 335964 274928 335970
rect 274876 335906 274928 335912
rect 275072 335902 275100 339743
rect 275256 338554 275284 342327
rect 275244 338548 275296 338554
rect 275244 338490 275296 338496
rect 275060 335896 275112 335902
rect 275060 335838 275112 335844
rect 270828 334468 270880 334474
rect 270828 334410 270880 334416
rect 279580 333794 279608 335836
rect 280304 333856 280356 333862
rect 280304 333798 280356 333804
rect 279568 333788 279620 333794
rect 279568 333730 279620 333736
rect 267148 333108 267200 333114
rect 267148 333050 267200 333056
rect 270736 333108 270788 333114
rect 270736 333050 270788 333056
rect 267160 332337 267188 333050
rect 267146 332328 267202 332337
rect 267146 332263 267202 332272
rect 266778 331240 266834 331249
rect 266778 331175 266834 331184
rect 267882 330288 267938 330297
rect 267882 330223 267938 330232
rect 267896 329170 267924 330223
rect 267884 329164 267936 329170
rect 267884 329106 267936 329112
rect 280316 324818 280344 333798
rect 282892 333153 282920 335836
rect 285928 335822 286218 335850
rect 288688 335822 289530 335850
rect 282878 333144 282934 333153
rect 282878 333079 282934 333088
rect 281776 327464 281828 327470
rect 281776 327406 281828 327412
rect 281788 327062 281816 327406
rect 282892 327062 282920 333079
rect 285928 328966 285956 335822
rect 285916 328960 285968 328966
rect 285916 328902 285968 328908
rect 285928 328286 285956 328902
rect 285916 328280 285968 328286
rect 285916 328222 285968 328228
rect 288688 327538 288716 335822
rect 292724 333924 292776 333930
rect 292724 333866 292776 333872
rect 288676 327532 288728 327538
rect 288676 327474 288728 327480
rect 288688 327130 288716 327474
rect 288676 327124 288728 327130
rect 288676 327066 288728 327072
rect 281776 327056 281828 327062
rect 281776 326998 281828 327004
rect 282880 327056 282932 327062
rect 282880 326998 282932 327004
rect 292736 324818 292764 333866
rect 292920 331657 292948 335836
rect 296232 333153 296260 335836
rect 296218 333144 296274 333153
rect 296218 333079 296274 333088
rect 296232 332201 296260 333079
rect 296218 332192 296274 332201
rect 296218 332127 296274 332136
rect 292906 331648 292962 331657
rect 292906 331583 292962 331592
rect 299544 331550 299572 335836
rect 302870 335822 303160 335850
rect 299532 331544 299584 331550
rect 299532 331486 299584 331492
rect 299544 329034 299572 331486
rect 299532 329028 299584 329034
rect 299532 328970 299584 328976
rect 303132 328966 303160 335822
rect 306260 334474 306288 335836
rect 306248 334468 306300 334474
rect 306248 334410 306300 334416
rect 305144 333992 305196 333998
rect 305144 333934 305196 333940
rect 303120 328960 303172 328966
rect 303120 328902 303172 328908
rect 303132 327606 303160 328902
rect 303120 327600 303172 327606
rect 303120 327542 303172 327548
rect 279108 324812 279160 324818
rect 279108 324754 279160 324760
rect 280304 324812 280356 324818
rect 280304 324754 280356 324760
rect 291528 324812 291580 324818
rect 291528 324754 291580 324760
rect 292724 324812 292776 324818
rect 292724 324754 292776 324760
rect 279120 321692 279148 324754
rect 291540 321692 291568 324754
rect 305156 324070 305184 333934
rect 306260 333561 306288 334410
rect 309572 333862 309600 335836
rect 312884 333930 312912 335836
rect 316196 333998 316224 335836
rect 316184 333992 316236 333998
rect 316184 333934 316236 333940
rect 312872 333924 312924 333930
rect 312872 333866 312924 333872
rect 309560 333856 309612 333862
rect 309560 333798 309612 333804
rect 306246 333552 306302 333561
rect 306246 333487 306302 333496
rect 316552 329096 316604 329102
rect 316552 329038 316604 329044
rect 304040 324064 304092 324070
rect 304040 324006 304092 324012
rect 305144 324064 305196 324070
rect 305144 324006 305196 324012
rect 304052 321692 304080 324006
rect 316564 321692 316592 329038
rect 319048 328966 319076 382039
rect 319140 334474 319168 384759
rect 319218 380200 319274 380209
rect 319218 380135 319274 380144
rect 319128 334468 319180 334474
rect 319128 334410 319180 334416
rect 319232 334082 319260 380135
rect 319310 377480 319366 377489
rect 319310 377415 319366 377424
rect 319140 334054 319260 334082
rect 319140 331754 319168 334054
rect 319324 333153 319352 377415
rect 319402 374760 319458 374769
rect 319402 374695 319458 374704
rect 319310 333144 319366 333153
rect 319310 333079 319366 333088
rect 319128 331748 319180 331754
rect 319128 331690 319180 331696
rect 319140 330462 319168 331690
rect 319416 331657 319444 374695
rect 320322 372176 320378 372185
rect 320322 372111 320378 372120
rect 320336 371806 320364 372111
rect 320324 371800 320376 371806
rect 320324 371742 320376 371748
rect 328420 357928 328472 357934
rect 328420 357870 328472 357876
rect 328432 357497 328460 357870
rect 328418 357488 328474 357497
rect 328418 357423 328474 357432
rect 328328 356568 328380 356574
rect 328328 356510 328380 356516
rect 328340 356137 328368 356510
rect 328326 356128 328382 356137
rect 328326 356063 328382 356072
rect 328420 355208 328472 355214
rect 328418 355176 328420 355185
rect 328472 355176 328474 355185
rect 328418 355111 328474 355120
rect 328512 355140 328564 355146
rect 328512 355082 328564 355088
rect 328524 354641 328552 355082
rect 328510 354632 328566 354641
rect 328510 354567 328566 354576
rect 328052 353848 328104 353854
rect 328052 353790 328104 353796
rect 328064 353417 328092 353790
rect 328050 353408 328106 353417
rect 328050 353343 328106 353352
rect 328512 352420 328564 352426
rect 328512 352362 328564 352368
rect 328524 352329 328552 352362
rect 328510 352320 328566 352329
rect 328510 352255 328566 352264
rect 320598 351368 320654 351377
rect 320598 351303 320654 351312
rect 320612 351134 320640 351303
rect 320600 351128 320652 351134
rect 320600 351070 320652 351076
rect 327224 351128 327276 351134
rect 327224 351070 327276 351076
rect 321610 350416 321666 350425
rect 321610 350351 321666 350360
rect 321624 349774 321652 350351
rect 321612 349768 321664 349774
rect 321612 349710 321664 349716
rect 327132 349768 327184 349774
rect 327132 349710 327184 349716
rect 320690 349600 320746 349609
rect 320690 349535 320746 349544
rect 320704 348346 320732 349535
rect 321610 348648 321666 348657
rect 321610 348583 321666 348592
rect 321624 348482 321652 348583
rect 321612 348476 321664 348482
rect 321612 348418 321664 348424
rect 327040 348476 327092 348482
rect 327040 348418 327092 348424
rect 320692 348340 320744 348346
rect 320692 348282 320744 348288
rect 321058 347832 321114 347841
rect 321058 347767 321114 347776
rect 321072 346986 321100 347767
rect 321060 346980 321112 346986
rect 321060 346922 321112 346928
rect 323176 346980 323228 346986
rect 323176 346922 323228 346928
rect 320506 346880 320562 346889
rect 320506 346815 320562 346824
rect 320520 345626 320548 346815
rect 321610 346064 321666 346073
rect 321610 345999 321666 346008
rect 321624 345762 321652 345999
rect 321612 345756 321664 345762
rect 321612 345698 321664 345704
rect 320508 345620 320560 345626
rect 320508 345562 320560 345568
rect 323188 345558 323216 346922
rect 327052 346481 327080 348418
rect 327144 348249 327172 349710
rect 327236 349609 327264 351070
rect 327868 351060 327920 351066
rect 327868 351002 327920 351008
rect 327498 350960 327554 350969
rect 327498 350895 327554 350904
rect 327512 350386 327540 350895
rect 327880 350425 327908 351002
rect 327866 350416 327922 350425
rect 327500 350380 327552 350386
rect 327866 350351 327922 350360
rect 327500 350322 327552 350328
rect 327222 349600 327278 349609
rect 327222 349535 327278 349544
rect 327224 348340 327276 348346
rect 327224 348282 327276 348288
rect 327130 348240 327186 348249
rect 327130 348175 327186 348184
rect 327236 346889 327264 348282
rect 327222 346880 327278 346889
rect 327222 346815 327278 346824
rect 327038 346472 327094 346481
rect 327038 346407 327094 346416
rect 326948 345756 327000 345762
rect 326948 345698 327000 345704
rect 323268 345620 323320 345626
rect 323268 345562 323320 345568
rect 323176 345552 323228 345558
rect 323176 345494 323228 345500
rect 323280 345370 323308 345562
rect 323188 345342 323308 345370
rect 320966 345112 321022 345121
rect 320966 345047 321022 345056
rect 320980 344538 321008 345047
rect 320968 344532 321020 344538
rect 320968 344474 321020 344480
rect 321610 344296 321666 344305
rect 321610 344231 321612 344240
rect 321664 344231 321666 344240
rect 321612 344202 321664 344208
rect 323188 344130 323216 345342
rect 323268 344532 323320 344538
rect 323268 344474 323320 344480
rect 323176 344124 323228 344130
rect 323176 344066 323228 344072
rect 321610 343344 321666 343353
rect 321610 343279 321666 343288
rect 321624 342906 321652 343279
rect 321612 342900 321664 342906
rect 321612 342842 321664 342848
rect 323280 342770 323308 344474
rect 323268 342764 323320 342770
rect 323268 342706 323320 342712
rect 326960 342673 326988 345698
rect 328052 345552 328104 345558
rect 328052 345494 328104 345500
rect 328064 345121 328092 345494
rect 328050 345112 328106 345121
rect 328050 345047 328106 345056
rect 327408 344260 327460 344266
rect 327408 344202 327460 344208
rect 327224 342900 327276 342906
rect 327224 342842 327276 342848
rect 326946 342664 327002 342673
rect 326946 342599 327002 342608
rect 321058 342392 321114 342401
rect 321058 342327 321114 342336
rect 321072 341546 321100 342327
rect 321610 341576 321666 341585
rect 321060 341540 321112 341546
rect 321610 341511 321666 341520
rect 327132 341540 327184 341546
rect 321060 341482 321112 341488
rect 321624 341478 321652 341511
rect 327132 341482 327184 341488
rect 321612 341472 321664 341478
rect 321612 341414 321664 341420
rect 327040 341472 327092 341478
rect 327040 341414 327092 341420
rect 320598 340624 320654 340633
rect 320598 340559 320654 340568
rect 320612 340118 320640 340559
rect 320600 340112 320652 340118
rect 320600 340054 320652 340060
rect 320506 339808 320562 339817
rect 320506 339743 320562 339752
rect 320414 338856 320470 338865
rect 320414 338791 320416 338800
rect 320468 338791 320470 338800
rect 320416 338762 320468 338768
rect 320520 338690 320548 339743
rect 326580 338820 326632 338826
rect 326580 338762 326632 338768
rect 320508 338684 320560 338690
rect 320508 338626 320560 338632
rect 320414 338040 320470 338049
rect 320414 337975 320470 337984
rect 320428 337330 320456 337975
rect 320416 337324 320468 337330
rect 320416 337266 320468 337272
rect 320414 337088 320470 337097
rect 320414 337023 320470 337032
rect 320428 336106 320456 337023
rect 320506 336272 320562 336281
rect 320506 336207 320562 336216
rect 320416 336100 320468 336106
rect 320416 336042 320468 336048
rect 319680 334468 319732 334474
rect 319680 334410 319732 334416
rect 319692 333182 319720 334410
rect 319680 333176 319732 333182
rect 319680 333118 319732 333124
rect 319862 333144 319918 333153
rect 319862 333079 319918 333088
rect 319876 331822 319904 333079
rect 319864 331816 319916 331822
rect 319864 331758 319916 331764
rect 320520 331754 320548 336207
rect 326592 334377 326620 338762
rect 327052 338185 327080 341414
rect 327144 338593 327172 341482
rect 327236 339953 327264 342842
rect 327420 341313 327448 344202
rect 328512 344124 328564 344130
rect 328512 344066 328564 344072
rect 328524 344033 328552 344066
rect 328510 344024 328566 344033
rect 328510 343959 328566 343968
rect 328052 342764 328104 342770
rect 328052 342706 328104 342712
rect 328064 342129 328092 342706
rect 328050 342120 328106 342129
rect 328050 342055 328106 342064
rect 327406 341304 327462 341313
rect 327406 341239 327462 341248
rect 327868 340112 327920 340118
rect 327868 340054 327920 340060
rect 327222 339944 327278 339953
rect 327222 339879 327278 339888
rect 327224 338684 327276 338690
rect 327224 338626 327276 338632
rect 327130 338584 327186 338593
rect 327130 338519 327186 338528
rect 327038 338176 327094 338185
rect 327038 338111 327094 338120
rect 326764 337324 326816 337330
rect 326764 337266 326816 337272
rect 326578 334368 326634 334377
rect 326578 334303 326634 334312
rect 326776 333969 326804 337266
rect 327236 335873 327264 338626
rect 327880 337097 327908 340054
rect 327866 337088 327922 337097
rect 327866 337023 327922 337032
rect 327316 336100 327368 336106
rect 327316 336042 327368 336048
rect 327222 335864 327278 335873
rect 327222 335799 327278 335808
rect 326762 333960 326818 333969
rect 326762 333895 326818 333904
rect 323820 333788 323872 333794
rect 323820 333730 323872 333736
rect 320508 331748 320560 331754
rect 320508 331690 320560 331696
rect 319402 331648 319458 331657
rect 319402 331583 319458 331592
rect 319678 331648 319734 331657
rect 319678 331583 319734 331592
rect 319692 330530 319720 331583
rect 319680 330524 319732 330530
rect 319680 330466 319732 330472
rect 319128 330456 319180 330462
rect 319128 330398 319180 330404
rect 319586 330288 319642 330297
rect 319586 330223 319642 330232
rect 319600 329238 319628 330223
rect 319588 329232 319640 329238
rect 319588 329174 319640 329180
rect 319036 328960 319088 328966
rect 319036 328902 319088 328908
rect 270274 313560 270330 313569
rect 270274 313495 270330 313504
rect 270288 313122 270316 313495
rect 270276 313116 270328 313122
rect 270276 313058 270328 313064
rect 270368 297204 270420 297210
rect 270368 297146 270420 297152
rect 270380 296841 270408 297146
rect 270366 296832 270422 296841
rect 270366 296767 270422 296776
rect 269264 286324 269316 286330
rect 269264 286266 269316 286272
rect 269276 280249 269304 286266
rect 269262 280240 269318 280249
rect 269262 280175 269318 280184
rect 276452 269670 276480 271916
rect 276440 269664 276492 269670
rect 276440 269606 276492 269612
rect 283536 269534 283564 271916
rect 290712 269670 290740 271916
rect 290700 269664 290752 269670
rect 290700 269606 290752 269612
rect 283524 269528 283576 269534
rect 283524 269470 283576 269476
rect 284536 269052 284588 269058
rect 284536 268994 284588 269000
rect 268620 268984 268672 268990
rect 268620 268926 268672 268932
rect 267240 263544 267292 263550
rect 267240 263486 267292 263492
rect 266594 256168 266650 256177
rect 266594 256103 266650 256112
rect 266608 255934 266636 256103
rect 266596 255928 266648 255934
rect 266596 255870 266648 255876
rect 266594 254672 266650 254681
rect 266594 254607 266650 254616
rect 266608 254574 266636 254607
rect 266596 254568 266648 254574
rect 266596 254510 266648 254516
rect 266594 253312 266650 253321
rect 266594 253247 266650 253256
rect 266608 253146 266636 253247
rect 266596 253140 266648 253146
rect 266596 253082 266648 253088
rect 266594 251952 266650 251961
rect 266594 251887 266650 251896
rect 266608 251786 266636 251887
rect 266596 251780 266648 251786
rect 266596 251722 266648 251728
rect 266596 250284 266648 250290
rect 266596 250226 266648 250232
rect 266608 249105 266636 250226
rect 266594 249096 266650 249105
rect 266594 249031 266650 249040
rect 266596 248924 266648 248930
rect 266596 248866 266648 248872
rect 266608 247745 266636 248866
rect 266594 247736 266650 247745
rect 266594 247671 266650 247680
rect 266596 246136 266648 246142
rect 266596 246078 266648 246084
rect 266608 244889 266636 246078
rect 266594 244880 266650 244889
rect 266594 244815 266650 244824
rect 266596 244776 266648 244782
rect 266596 244718 266648 244724
rect 266608 243529 266636 244718
rect 266594 243520 266650 243529
rect 266594 243455 266650 243464
rect 266778 239304 266834 239313
rect 266778 239239 266834 239248
rect 266792 239206 266820 239239
rect 266780 239200 266832 239206
rect 266780 239142 266832 239148
rect 267252 236593 267280 263486
rect 267422 263104 267478 263113
rect 267422 263039 267478 263048
rect 267330 258888 267386 258897
rect 267330 258823 267386 258832
rect 267344 252398 267372 258823
rect 267332 252392 267384 252398
rect 267332 252334 267384 252340
rect 267330 250592 267386 250601
rect 267330 250527 267386 250536
rect 267344 237234 267372 250527
rect 267436 250222 267464 263039
rect 267514 261744 267570 261753
rect 267514 261679 267570 261688
rect 267424 250216 267476 250222
rect 267424 250158 267476 250164
rect 267528 248862 267556 261679
rect 267606 260384 267662 260393
rect 267606 260319 267662 260328
rect 267516 248856 267568 248862
rect 267516 248798 267568 248804
rect 267620 248794 267648 260319
rect 267790 257528 267846 257537
rect 267790 257463 267846 257472
rect 267804 252482 267832 257463
rect 267884 254500 267936 254506
rect 267884 254442 267936 254448
rect 267712 252454 267832 252482
rect 267608 248788 267660 248794
rect 267608 248730 267660 248736
rect 267712 246210 267740 252454
rect 267792 252392 267844 252398
rect 267792 252334 267844 252340
rect 267804 247570 267832 252334
rect 267792 247564 267844 247570
rect 267792 247506 267844 247512
rect 267896 246385 267924 254442
rect 267882 246376 267938 246385
rect 267882 246311 267938 246320
rect 267700 246204 267752 246210
rect 267700 246146 267752 246152
rect 267884 242192 267936 242198
rect 267882 242160 267884 242169
rect 267936 242160 267938 242169
rect 267882 242095 267938 242104
rect 267882 240664 267938 240673
rect 267882 240599 267884 240608
rect 267936 240599 267938 240608
rect 267884 240570 267936 240576
rect 267608 239268 267660 239274
rect 267608 239210 267660 239216
rect 267620 237953 267648 239210
rect 267606 237944 267662 237953
rect 267606 237879 267662 237888
rect 267332 237228 267384 237234
rect 267332 237170 267384 237176
rect 267238 236584 267294 236593
rect 267238 236519 267294 236528
rect 268632 175694 268660 268926
rect 284548 257772 284576 268994
rect 290712 268990 290740 269606
rect 297796 269058 297824 271916
rect 304972 269398 305000 271916
rect 312056 269398 312084 271916
rect 303764 269392 303816 269398
rect 303764 269334 303816 269340
rect 304960 269392 305012 269398
rect 304960 269334 305012 269340
rect 310756 269392 310808 269398
rect 310756 269334 310808 269340
rect 312044 269392 312096 269398
rect 312044 269334 312096 269340
rect 297784 269052 297836 269058
rect 297784 268994 297836 269000
rect 290700 268984 290752 268990
rect 290700 268926 290752 268932
rect 303776 261306 303804 269334
rect 310768 264094 310796 269334
rect 310756 264088 310808 264094
rect 310756 264030 310808 264036
rect 310768 263550 310796 264030
rect 310756 263544 310808 263550
rect 310756 263486 310808 263492
rect 297876 261300 297928 261306
rect 297876 261242 297928 261248
rect 303764 261300 303816 261306
rect 303764 261242 303816 261248
rect 297888 257772 297916 261242
rect 319232 260694 319260 271916
rect 311216 260688 311268 260694
rect 311216 260630 311268 260636
rect 319220 260688 319272 260694
rect 319220 260630 319272 260636
rect 311228 257772 311256 260630
rect 321060 258580 321112 258586
rect 321060 258522 321112 258528
rect 321072 257401 321100 258522
rect 276162 257392 276218 257401
rect 276162 257327 276218 257336
rect 321058 257392 321114 257401
rect 321058 257327 321114 257336
rect 274966 256440 275022 256449
rect 274966 256375 275022 256384
rect 271380 255928 271432 255934
rect 271380 255870 271432 255876
rect 271392 246074 271420 255870
rect 274874 255624 274930 255633
rect 274874 255559 274930 255568
rect 272760 254568 272812 254574
rect 272760 254510 272812 254516
rect 271472 251780 271524 251786
rect 271472 251722 271524 251728
rect 271380 246068 271432 246074
rect 271380 246010 271432 246016
rect 271484 242198 271512 251722
rect 272772 244782 272800 254510
rect 274888 254506 274916 255559
rect 274876 254500 274928 254506
rect 274876 254442 274928 254448
rect 272852 253140 272904 253146
rect 272852 253082 272904 253088
rect 272760 244776 272812 244782
rect 272760 244718 272812 244724
rect 272864 243422 272892 253082
rect 274874 252904 274930 252913
rect 274874 252839 274930 252848
rect 274888 251786 274916 252839
rect 274876 251780 274928 251786
rect 274876 251722 274928 251728
rect 274876 250216 274928 250222
rect 274876 250158 274928 250164
rect 274888 250057 274916 250158
rect 274874 250048 274930 250057
rect 274874 249983 274930 249992
rect 274980 248930 275008 256375
rect 275794 254672 275850 254681
rect 275794 254607 275850 254616
rect 275610 252088 275666 252097
rect 275610 252023 275666 252032
rect 275518 251136 275574 251145
rect 275518 251071 275574 251080
rect 274968 248924 275020 248930
rect 274968 248866 275020 248872
rect 274876 248856 274928 248862
rect 274874 248824 274876 248833
rect 274928 248824 274930 248833
rect 274874 248759 274930 248768
rect 274968 248788 275020 248794
rect 274968 248730 275020 248736
rect 274980 248289 275008 248730
rect 274966 248280 275022 248289
rect 274966 248215 275022 248224
rect 274876 247564 274928 247570
rect 274876 247506 274928 247512
rect 274888 247337 274916 247506
rect 274874 247328 274930 247337
rect 274874 247263 274930 247272
rect 274876 246204 274928 246210
rect 274876 246146 274928 246152
rect 274888 246113 274916 246146
rect 274874 246104 274930 246113
rect 274874 246039 274930 246048
rect 274968 246068 275020 246074
rect 274968 246010 275020 246016
rect 274980 245569 275008 246010
rect 274966 245560 275022 245569
rect 274966 245495 275022 245504
rect 274876 244776 274928 244782
rect 274876 244718 274928 244724
rect 274888 244617 274916 244718
rect 274874 244608 274930 244617
rect 274874 244543 274930 244552
rect 272852 243416 272904 243422
rect 275428 243416 275480 243422
rect 272852 243358 272904 243364
rect 275426 243384 275428 243393
rect 275480 243384 275482 243393
rect 275426 243319 275482 243328
rect 271472 242192 271524 242198
rect 271472 242134 271524 242140
rect 275532 239206 275560 251071
rect 275624 240634 275652 252023
rect 275702 250320 275758 250329
rect 275702 250255 275758 250264
rect 275612 240628 275664 240634
rect 275612 240570 275664 240576
rect 275716 239274 275744 250255
rect 275808 246142 275836 254607
rect 275886 253856 275942 253865
rect 275886 253791 275942 253800
rect 275796 246136 275848 246142
rect 275796 246078 275848 246084
rect 275900 244646 275928 253791
rect 275980 251916 276032 251922
rect 275980 251858 276032 251864
rect 275888 244640 275940 244646
rect 275888 244582 275940 244588
rect 275992 242849 276020 251858
rect 276176 250290 276204 257327
rect 321060 257220 321112 257226
rect 321060 257162 321112 257168
rect 321072 256449 321100 257162
rect 321058 256440 321114 256449
rect 321058 256375 321114 256384
rect 320600 255860 320652 255866
rect 320600 255802 320652 255808
rect 320612 254681 320640 255802
rect 321612 255792 321664 255798
rect 321612 255734 321664 255740
rect 321624 255633 321652 255734
rect 321610 255624 321666 255633
rect 321610 255559 321666 255568
rect 320598 254672 320654 254681
rect 320598 254607 320654 254616
rect 320508 254500 320560 254506
rect 320508 254442 320560 254448
rect 320520 252913 320548 254442
rect 321612 253956 321664 253962
rect 321612 253898 321664 253904
rect 321624 253865 321652 253898
rect 321610 253856 321666 253865
rect 321610 253791 321666 253800
rect 320506 252904 320562 252913
rect 320506 252839 320562 252848
rect 321610 252088 321666 252097
rect 321610 252023 321666 252032
rect 321624 251922 321652 252023
rect 321612 251916 321664 251922
rect 321612 251858 321664 251864
rect 321610 251136 321666 251145
rect 321610 251071 321666 251080
rect 321624 251038 321652 251071
rect 321612 251032 321664 251038
rect 321612 250974 321664 250980
rect 321058 250320 321114 250329
rect 276164 250284 276216 250290
rect 321058 250255 321114 250264
rect 276164 250226 276216 250232
rect 321072 249542 321100 250255
rect 321060 249536 321112 249542
rect 321060 249478 321112 249484
rect 321610 249368 321666 249377
rect 321610 249303 321666 249312
rect 321624 249134 321652 249303
rect 321612 249128 321664 249134
rect 321612 249070 321664 249076
rect 321610 248416 321666 248425
rect 321610 248351 321666 248360
rect 321624 247706 321652 248351
rect 321612 247700 321664 247706
rect 321612 247642 321664 247648
rect 321794 247600 321850 247609
rect 321794 247535 321796 247544
rect 321848 247535 321850 247544
rect 321796 247506 321848 247512
rect 321808 247475 321836 247506
rect 321426 246648 321482 246657
rect 321426 246583 321482 246592
rect 321440 246278 321468 246583
rect 321428 246272 321480 246278
rect 321428 246214 321480 246220
rect 321610 245832 321666 245841
rect 321610 245767 321666 245776
rect 321624 244850 321652 245767
rect 321704 244912 321756 244918
rect 321702 244880 321704 244889
rect 323176 244912 323228 244918
rect 321756 244880 321758 244889
rect 321612 244844 321664 244850
rect 323176 244854 323228 244860
rect 321702 244815 321758 244824
rect 321612 244786 321664 244792
rect 321610 244064 321666 244073
rect 321610 243999 321666 244008
rect 321624 243490 321652 243999
rect 321612 243484 321664 243490
rect 321612 243426 321664 243432
rect 323188 243422 323216 244854
rect 323176 243416 323228 243422
rect 323176 243358 323228 243364
rect 321610 243112 321666 243121
rect 321610 243047 321666 243056
rect 275978 242840 276034 242849
rect 275978 242775 276034 242784
rect 320506 242296 320562 242305
rect 321624 242266 321652 243047
rect 320506 242231 320562 242240
rect 321612 242260 321664 242266
rect 320520 242130 320548 242231
rect 321612 242202 321664 242208
rect 320508 242124 320560 242130
rect 320508 242066 320560 242072
rect 279672 239342 279700 241860
rect 283260 239449 283288 241860
rect 283246 239440 283302 239449
rect 283246 239375 283302 239384
rect 279660 239336 279712 239342
rect 279660 239278 279712 239284
rect 280304 239336 280356 239342
rect 280304 239278 280356 239284
rect 275704 239268 275756 239274
rect 275704 239210 275756 239216
rect 275520 239200 275572 239206
rect 275520 239142 275572 239148
rect 279108 230292 279160 230298
rect 279108 230234 279160 230240
rect 279120 227716 279148 230234
rect 280316 227646 280344 239278
rect 286940 236321 286968 241860
rect 290528 238594 290556 241860
rect 294208 239857 294236 241860
rect 297796 241738 297824 241860
rect 301476 241738 301504 241860
rect 296968 241710 297824 241738
rect 301108 241710 301504 241738
rect 305064 241738 305092 241860
rect 308744 241738 308772 241860
rect 312332 241738 312360 241860
rect 316026 241846 316132 241874
rect 305064 241710 305184 241738
rect 294194 239848 294250 239857
rect 294194 239783 294250 239792
rect 290056 238588 290108 238594
rect 290056 238530 290108 238536
rect 290516 238588 290568 238594
rect 290516 238530 290568 238536
rect 290068 238497 290096 238530
rect 290054 238488 290110 238497
rect 290054 238423 290110 238432
rect 296968 236350 296996 241710
rect 296956 236344 297008 236350
rect 286926 236312 286982 236321
rect 296956 236286 297008 236292
rect 298244 236344 298296 236350
rect 298244 236286 298296 236292
rect 286926 236247 286982 236256
rect 286940 235874 286968 236247
rect 298256 235942 298284 236286
rect 298244 235936 298296 235942
rect 298244 235878 298296 235884
rect 286928 235868 286980 235874
rect 286928 235810 286980 235816
rect 301108 234961 301136 241710
rect 305156 240401 305184 241710
rect 308008 241710 308772 241738
rect 312148 241710 312360 241738
rect 305142 240392 305198 240401
rect 305142 240327 305198 240336
rect 301094 234952 301150 234961
rect 301094 234887 301150 234896
rect 301108 234446 301136 234887
rect 301096 234440 301148 234446
rect 301096 234382 301148 234388
rect 304040 230428 304092 230434
rect 304040 230370 304092 230376
rect 291528 230360 291580 230366
rect 291528 230302 291580 230308
rect 291540 227716 291568 230302
rect 304052 227716 304080 230370
rect 305156 227714 305184 240327
rect 308008 230298 308036 241710
rect 312148 230366 312176 241710
rect 316104 239886 316132 241846
rect 314896 239880 314948 239886
rect 314896 239822 314948 239828
rect 316092 239880 316144 239886
rect 316092 239822 316144 239828
rect 314908 230434 314936 239822
rect 316276 237228 316328 237234
rect 316276 237170 316328 237176
rect 316288 236622 316316 237170
rect 316276 236616 316328 236622
rect 316276 236558 316328 236564
rect 314896 230428 314948 230434
rect 314896 230370 314948 230376
rect 312136 230360 312188 230366
rect 312136 230302 312188 230308
rect 307996 230292 308048 230298
rect 307996 230234 308048 230240
rect 316288 227730 316316 236558
rect 323832 233766 323860 333730
rect 325384 333176 325436 333182
rect 325384 333118 325436 333124
rect 325200 331816 325252 331822
rect 325200 331758 325252 331764
rect 324740 328960 324792 328966
rect 324740 328902 324792 328908
rect 324556 322772 324608 322778
rect 324556 322714 324608 322720
rect 324568 320369 324596 322714
rect 324752 320738 324780 328902
rect 325108 327124 325160 327130
rect 325108 327066 325160 327072
rect 325120 324886 325148 327066
rect 325108 324880 325160 324886
rect 325108 324822 325160 324828
rect 324740 320732 324792 320738
rect 324740 320674 324792 320680
rect 324554 320360 324610 320369
rect 324554 320295 324610 320304
rect 324752 317241 324780 320674
rect 325120 320058 325148 324822
rect 325212 322234 325240 331758
rect 325292 330456 325344 330462
rect 325292 330398 325344 330404
rect 325200 322228 325252 322234
rect 325200 322170 325252 322176
rect 325108 320052 325160 320058
rect 325108 319994 325160 320000
rect 324738 317232 324794 317241
rect 324738 317167 324794 317176
rect 325212 310985 325240 322170
rect 325304 319378 325332 330398
rect 325396 322778 325424 333118
rect 327328 333017 327356 336042
rect 327314 333008 327370 333017
rect 327314 332943 327370 332952
rect 328512 331748 328564 331754
rect 328512 331690 328564 331696
rect 328524 331521 328552 331690
rect 328510 331512 328566 331521
rect 328510 331447 328566 331456
rect 325752 330524 325804 330530
rect 325752 330466 325804 330472
rect 325660 328280 325712 328286
rect 325660 328222 325712 328228
rect 325568 327056 325620 327062
rect 325568 326998 325620 327004
rect 325384 322772 325436 322778
rect 325384 322714 325436 322720
rect 325396 322166 325424 322714
rect 325384 322160 325436 322166
rect 325384 322102 325436 322108
rect 325580 320194 325608 326998
rect 325672 320806 325700 328222
rect 325764 323526 325792 330466
rect 330088 329838 331298 329866
rect 331468 329838 332034 329866
rect 326580 326920 326632 326926
rect 326580 326862 326632 326868
rect 325752 323520 325804 323526
rect 325752 323462 325804 323468
rect 325660 320800 325712 320806
rect 325660 320742 325712 320748
rect 325568 320188 325620 320194
rect 325568 320130 325620 320136
rect 325568 320052 325620 320058
rect 325568 319994 325620 320000
rect 325476 319440 325528 319446
rect 325476 319382 325528 319388
rect 325292 319372 325344 319378
rect 325292 319314 325344 319320
rect 325292 314476 325344 314482
rect 325292 314418 325344 314424
rect 325198 310976 325254 310985
rect 325198 310911 325254 310920
rect 325106 305536 325162 305545
rect 325106 305471 325162 305480
rect 325120 298473 325148 305471
rect 325106 298464 325162 298473
rect 325106 298399 325162 298408
rect 324554 292208 324610 292217
rect 324554 292143 324610 292152
rect 323820 233760 323872 233766
rect 323820 233702 323872 233708
rect 305144 227708 305196 227714
rect 316288 227702 316578 227730
rect 322992 227708 323044 227714
rect 305144 227650 305196 227656
rect 322992 227650 323044 227656
rect 280304 227640 280356 227646
rect 280304 227582 280356 227588
rect 323004 226393 323032 227650
rect 322990 226384 323046 226393
rect 322990 226319 323046 226328
rect 322532 224172 322584 224178
rect 322532 224114 322584 224120
rect 272942 219584 272998 219593
rect 272942 219519 272998 219528
rect 272956 219282 272984 219519
rect 272944 219276 272996 219282
rect 272944 219218 272996 219224
rect 272944 203364 272996 203370
rect 272944 203306 272996 203312
rect 272956 202865 272984 203306
rect 272942 202856 272998 202865
rect 272942 202791 272998 202800
rect 273128 192416 273180 192422
rect 273128 192358 273180 192364
rect 273140 186273 273168 192358
rect 273126 186264 273182 186273
rect 273126 186199 273182 186208
rect 276452 175830 276480 177940
rect 276440 175824 276492 175830
rect 276440 175766 276492 175772
rect 283536 175762 283564 177940
rect 283524 175756 283576 175762
rect 283524 175698 283576 175704
rect 290712 175694 290740 177940
rect 268620 175688 268672 175694
rect 268620 175630 268672 175636
rect 290700 175688 290752 175694
rect 290700 175630 290752 175636
rect 297796 175150 297824 177940
rect 285824 175144 285876 175150
rect 285824 175086 285876 175092
rect 297784 175144 297836 175150
rect 297784 175086 297836 175092
rect 267240 169568 267292 169574
rect 267240 169510 267292 169516
rect 267146 164912 267202 164921
rect 267146 164847 267202 164856
rect 267054 162192 267110 162201
rect 267054 162127 267110 162136
rect 266872 162088 266924 162094
rect 266872 162030 266924 162036
rect 266596 160728 266648 160734
rect 266594 160696 266596 160705
rect 266648 160696 266650 160705
rect 266594 160631 266650 160640
rect 266594 159336 266650 159345
rect 266594 159271 266596 159280
rect 266648 159271 266650 159280
rect 266596 159242 266648 159248
rect 266596 158008 266648 158014
rect 266594 157976 266596 157985
rect 266648 157976 266650 157985
rect 266594 157911 266650 157920
rect 266594 155120 266650 155129
rect 266594 155055 266650 155064
rect 266608 155022 266636 155055
rect 266596 155016 266648 155022
rect 266596 154958 266648 154964
rect 266884 153769 266912 162030
rect 266964 160796 267016 160802
rect 266964 160738 267016 160744
rect 266870 153760 266926 153769
rect 266870 153695 266926 153704
rect 266976 152409 267004 160738
rect 267068 154954 267096 162127
rect 267056 154948 267108 154954
rect 267056 154890 267108 154896
rect 267160 153730 267188 164847
rect 267148 153724 267200 153730
rect 267148 153666 267200 153672
rect 266962 152400 267018 152409
rect 266962 152335 267018 152344
rect 266594 150904 266650 150913
rect 266594 150839 266596 150848
rect 266648 150839 266650 150848
rect 266596 150810 266648 150816
rect 266594 149544 266650 149553
rect 266594 149479 266650 149488
rect 266608 149446 266636 149479
rect 266596 149440 266648 149446
rect 266596 149382 266648 149388
rect 266596 148216 266648 148222
rect 266594 148184 266596 148193
rect 266648 148184 266650 148193
rect 266594 148119 266650 148128
rect 266780 145428 266832 145434
rect 266780 145370 266832 145376
rect 266792 145337 266820 145370
rect 266778 145328 266834 145337
rect 266778 145263 266834 145272
rect 267252 142617 267280 169510
rect 267422 169128 267478 169137
rect 267422 169063 267478 169072
rect 267332 160796 267384 160802
rect 267332 160738 267384 160744
rect 267344 160666 267372 160738
rect 267332 160660 267384 160666
rect 267332 160602 267384 160608
rect 267330 156616 267386 156625
rect 267330 156551 267386 156560
rect 267238 142608 267294 142617
rect 267238 142543 267294 142552
rect 267344 142034 267372 156551
rect 267436 156450 267464 169063
rect 267698 167768 267754 167777
rect 267698 167703 267754 167712
rect 267514 166408 267570 166417
rect 267514 166343 267570 166352
rect 267424 156444 267476 156450
rect 267424 156386 267476 156392
rect 267528 153662 267556 166343
rect 267712 155090 267740 167703
rect 285836 166310 285864 175086
rect 304972 166854 305000 177940
rect 312056 170254 312084 177940
rect 312044 170248 312096 170254
rect 312044 170190 312096 170196
rect 312056 169574 312084 170190
rect 312044 169568 312096 169574
rect 312044 169510 312096 169516
rect 319232 166854 319260 177940
rect 297876 166848 297928 166854
rect 297876 166790 297928 166796
rect 304960 166848 305012 166854
rect 304960 166790 305012 166796
rect 311216 166848 311268 166854
rect 311216 166790 311268 166796
rect 319220 166848 319272 166854
rect 319220 166790 319272 166796
rect 284536 166304 284588 166310
rect 284536 166246 284588 166252
rect 285824 166304 285876 166310
rect 285824 166246 285876 166252
rect 284548 163796 284576 166246
rect 297888 163796 297916 166790
rect 311228 163796 311256 166790
rect 321796 164808 321848 164814
rect 321796 164750 321848 164756
rect 267882 163552 267938 163561
rect 267882 163487 267938 163496
rect 321612 163516 321664 163522
rect 267792 155152 267844 155158
rect 267792 155094 267844 155100
rect 267700 155084 267752 155090
rect 267700 155026 267752 155032
rect 267700 154948 267752 154954
rect 267700 154890 267752 154896
rect 267516 153656 267568 153662
rect 267516 153598 267568 153604
rect 267712 150942 267740 154890
rect 267700 150936 267752 150942
rect 267700 150878 267752 150884
rect 267804 143977 267832 155094
rect 267896 152370 267924 163487
rect 321612 163458 321664 163464
rect 321624 163425 321652 163458
rect 274506 163416 274562 163425
rect 321610 163416 321666 163425
rect 274506 163351 274562 163360
rect 320968 163380 321020 163386
rect 274324 160728 274376 160734
rect 274324 160670 274376 160676
rect 271380 160660 271432 160666
rect 271380 160602 271432 160608
rect 267884 152364 267936 152370
rect 267884 152306 267936 152312
rect 271392 150874 271420 160602
rect 274232 159300 274284 159306
rect 274232 159242 274284 159248
rect 274138 158928 274194 158937
rect 274138 158863 274194 158872
rect 271380 150868 271432 150874
rect 271380 150810 271432 150816
rect 274152 148222 274180 158863
rect 274244 149553 274272 159242
rect 274336 150641 274364 160670
rect 274416 158008 274468 158014
rect 274416 157950 274468 157956
rect 274322 150632 274378 150641
rect 274322 150567 274378 150576
rect 274230 149544 274286 149553
rect 274230 149479 274286 149488
rect 274428 148873 274456 157950
rect 274520 155022 274548 163351
rect 321610 163351 321666 163360
rect 320968 163322 321020 163328
rect 320980 162473 321008 163322
rect 274874 162464 274930 162473
rect 274874 162399 274930 162408
rect 320966 162464 321022 162473
rect 320966 162399 321022 162408
rect 274888 162094 274916 162399
rect 274876 162088 274928 162094
rect 274876 162030 274928 162036
rect 321704 162088 321756 162094
rect 321704 162030 321756 162036
rect 274874 161648 274930 161657
rect 274874 161583 274930 161592
rect 274888 160802 274916 161583
rect 320784 161340 320836 161346
rect 320784 161282 320836 161288
rect 274876 160796 274928 160802
rect 274876 160738 274928 160744
rect 320796 160705 320824 161282
rect 274874 160696 274930 160705
rect 274874 160631 274876 160640
rect 274928 160631 274930 160640
rect 320782 160696 320838 160705
rect 320782 160631 320838 160640
rect 274876 160602 274928 160608
rect 321716 159889 321744 162030
rect 321808 161929 321836 164750
rect 321794 161920 321850 161929
rect 321794 161855 321850 161864
rect 275702 159880 275758 159889
rect 275702 159815 275758 159824
rect 321702 159880 321758 159889
rect 321702 159815 321758 159824
rect 275518 158112 275574 158121
rect 275518 158047 275574 158056
rect 274876 156444 274928 156450
rect 274876 156386 274928 156392
rect 274888 156081 274916 156386
rect 274966 156344 275022 156353
rect 274966 156279 275022 156288
rect 274874 156072 274930 156081
rect 274874 156007 274930 156016
rect 274980 155158 275008 156279
rect 274968 155152 275020 155158
rect 274968 155094 275020 155100
rect 274876 155084 274928 155090
rect 274876 155026 274928 155032
rect 274508 155016 274560 155022
rect 274888 154993 274916 155026
rect 274508 154958 274560 154964
rect 274874 154984 274930 154993
rect 274874 154919 274930 154928
rect 274968 153724 275020 153730
rect 274968 153666 275020 153672
rect 274876 153656 274928 153662
rect 274874 153624 274876 153633
rect 274928 153624 274930 153633
rect 274874 153559 274930 153568
rect 274980 153361 275008 153666
rect 274966 153352 275022 153361
rect 274966 153287 275022 153296
rect 274876 152364 274928 152370
rect 274876 152306 274928 152312
rect 274888 152137 274916 152306
rect 274874 152128 274930 152137
rect 274874 152063 274930 152072
rect 274876 150936 274928 150942
rect 274874 150904 274876 150913
rect 274928 150904 274930 150913
rect 274874 150839 274930 150848
rect 274414 148864 274470 148873
rect 274414 148799 274470 148808
rect 274140 148216 274192 148222
rect 274140 148158 274192 148164
rect 275532 146794 275560 158047
rect 275610 157160 275666 157169
rect 275610 157095 275666 157104
rect 267884 146788 267936 146794
rect 267884 146730 267936 146736
rect 275520 146788 275572 146794
rect 275520 146730 275572 146736
rect 267896 146697 267924 146730
rect 267882 146688 267938 146697
rect 267882 146623 267938 146632
rect 275624 145434 275652 157095
rect 275716 149446 275744 159815
rect 321058 158928 321114 158937
rect 321058 158863 321114 158872
rect 321072 158082 321100 158863
rect 321612 158212 321664 158218
rect 321612 158154 321664 158160
rect 321624 158121 321652 158154
rect 321610 158112 321666 158121
rect 321060 158076 321112 158082
rect 321610 158047 321666 158056
rect 321060 158018 321112 158024
rect 321612 157260 321664 157266
rect 321612 157202 321664 157208
rect 321624 157169 321652 157202
rect 321610 157160 321666 157169
rect 321610 157095 321666 157104
rect 321610 156344 321666 156353
rect 321610 156279 321666 156288
rect 321624 155974 321652 156279
rect 321612 155968 321664 155974
rect 321612 155910 321664 155916
rect 321610 155392 321666 155401
rect 321610 155327 321666 155336
rect 321624 155158 321652 155327
rect 321612 155152 321664 155158
rect 321612 155094 321664 155100
rect 320874 154440 320930 154449
rect 320874 154375 320930 154384
rect 320888 153798 320916 154375
rect 320876 153792 320928 153798
rect 320876 153734 320928 153740
rect 321610 153624 321666 153633
rect 321610 153559 321666 153568
rect 320506 152672 320562 152681
rect 320506 152607 320562 152616
rect 320520 152506 320548 152607
rect 320508 152500 320560 152506
rect 320508 152442 320560 152448
rect 321624 152438 321652 153559
rect 321612 152432 321664 152438
rect 321612 152374 321664 152380
rect 320782 151856 320838 151865
rect 320782 151791 320838 151800
rect 320796 151418 320824 151791
rect 320784 151412 320836 151418
rect 320784 151354 320836 151360
rect 321058 150904 321114 150913
rect 321058 150839 321114 150848
rect 321072 149650 321100 150839
rect 321610 150088 321666 150097
rect 321610 150023 321666 150032
rect 321624 149786 321652 150023
rect 321612 149780 321664 149786
rect 321612 149722 321664 149728
rect 321060 149644 321112 149650
rect 321060 149586 321112 149592
rect 275704 149440 275756 149446
rect 275704 149382 275756 149388
rect 321610 149136 321666 149145
rect 321610 149071 321666 149080
rect 321624 148426 321652 149071
rect 321612 148420 321664 148426
rect 321612 148362 321664 148368
rect 321702 148320 321758 148329
rect 321758 148278 321836 148306
rect 321702 148255 321758 148264
rect 279672 145434 279700 147884
rect 283260 147762 283288 147884
rect 286940 147762 286968 147884
rect 283168 147734 283288 147762
rect 285928 147734 286968 147762
rect 275612 145428 275664 145434
rect 275612 145370 275664 145376
rect 279660 145428 279712 145434
rect 279660 145370 279712 145376
rect 280304 144816 280356 144822
rect 280304 144758 280356 144764
rect 267790 143968 267846 143977
rect 267790 143903 267846 143912
rect 267332 142028 267384 142034
rect 267332 141970 267384 141976
rect 280316 136186 280344 144758
rect 283168 138537 283196 147734
rect 283154 138528 283210 138537
rect 283154 138463 283210 138472
rect 284442 138528 284498 138537
rect 284442 138463 284498 138472
rect 284456 137886 284484 138463
rect 284444 137880 284496 137886
rect 284444 137822 284496 137828
rect 279108 136180 279160 136186
rect 279108 136122 279160 136128
rect 280304 136180 280356 136186
rect 280304 136122 280356 136128
rect 279120 133740 279148 136122
rect 285928 135817 285956 147734
rect 290528 144754 290556 147884
rect 292724 144884 292776 144890
rect 292724 144826 292776 144832
rect 290516 144748 290568 144754
rect 290516 144690 290568 144696
rect 290528 144521 290556 144690
rect 290514 144512 290570 144521
rect 290514 144447 290570 144456
rect 292736 136322 292764 144826
rect 294208 144770 294236 147884
rect 297796 147762 297824 147884
rect 301476 147762 301504 147884
rect 296968 147734 297824 147762
rect 301108 147734 301504 147762
rect 294208 144742 294328 144770
rect 294300 143394 294328 144742
rect 294288 143388 294340 143394
rect 294288 143330 294340 143336
rect 294300 143161 294328 143330
rect 294286 143152 294342 143161
rect 294286 143087 294342 143096
rect 296968 137857 296996 147734
rect 301108 141121 301136 147734
rect 305064 142102 305092 147884
rect 308744 144822 308772 147884
rect 312332 144890 312360 147884
rect 312320 144884 312372 144890
rect 312320 144826 312372 144832
rect 308732 144816 308784 144822
rect 308732 144758 308784 144764
rect 316012 144142 316040 147884
rect 312780 144136 312832 144142
rect 312780 144078 312832 144084
rect 316000 144136 316052 144142
rect 316000 144078 316052 144084
rect 305052 142096 305104 142102
rect 305052 142038 305104 142044
rect 301094 141112 301150 141121
rect 301094 141047 301150 141056
rect 301108 140606 301136 141047
rect 301096 140600 301148 140606
rect 301096 140542 301148 140548
rect 296954 137848 297010 137857
rect 296954 137783 297010 137792
rect 312792 136458 312820 144078
rect 321808 144074 321836 148278
rect 321796 144068 321848 144074
rect 321796 144010 321848 144016
rect 316276 142028 316328 142034
rect 316276 141970 316328 141976
rect 316288 141354 316316 141970
rect 316276 141348 316328 141354
rect 316276 141290 316328 141296
rect 304040 136452 304092 136458
rect 304040 136394 304092 136400
rect 312780 136452 312832 136458
rect 312780 136394 312832 136400
rect 291528 136316 291580 136322
rect 291528 136258 291580 136264
rect 292724 136316 292776 136322
rect 292724 136258 292776 136264
rect 285914 135808 285970 135817
rect 285914 135743 285970 135752
rect 286742 135808 286798 135817
rect 286742 135743 286798 135752
rect 286756 135098 286784 135743
rect 286744 135092 286796 135098
rect 286744 135034 286796 135040
rect 291540 133740 291568 136258
rect 304052 133740 304080 136394
rect 316288 133754 316316 141290
rect 316288 133726 316578 133754
rect 270366 125472 270422 125481
rect 270366 125407 270422 125416
rect 270380 125306 270408 125407
rect 270368 125300 270420 125306
rect 270368 125242 270420 125248
rect 270000 117956 270052 117962
rect 270000 117898 270052 117904
rect 270012 108889 270040 117898
rect 269998 108880 270054 108889
rect 269998 108815 270054 108824
rect 267240 98576 267292 98582
rect 267240 98518 267292 98524
rect 267252 93006 267280 98518
rect 267240 93000 267292 93006
rect 267240 92942 267292 92948
rect 270368 93000 270420 93006
rect 270368 92942 270420 92948
rect 270380 92297 270408 92942
rect 270366 92288 270422 92297
rect 270366 92223 270422 92232
rect 276360 83814 276466 83842
rect 283168 83814 283550 83842
rect 290344 83814 290726 83842
rect 297520 83814 297810 83842
rect 304880 83814 304986 83842
rect 311872 83814 312070 83842
rect 319140 83814 319246 83842
rect 276360 81990 276388 83814
rect 276348 81984 276400 81990
rect 276348 81926 276400 81932
rect 276360 81310 276388 81926
rect 283168 81922 283196 83814
rect 283156 81916 283208 81922
rect 283156 81858 283208 81864
rect 290344 81854 290372 83814
rect 290332 81848 290384 81854
rect 290332 81790 290384 81796
rect 297520 81378 297548 83814
rect 304880 83706 304908 83814
rect 304880 83678 305092 83706
rect 285824 81372 285876 81378
rect 285824 81314 285876 81320
rect 297508 81372 297560 81378
rect 297508 81314 297560 81320
rect 276348 81304 276400 81310
rect 276348 81246 276400 81252
rect 266596 76408 266648 76414
rect 266596 76350 266648 76356
rect 266608 75297 266636 76350
rect 266594 75288 266650 75297
rect 266594 75223 266650 75232
rect 266594 74200 266650 74209
rect 266594 74135 266650 74144
rect 266608 73762 266636 74135
rect 266596 73756 266648 73762
rect 266596 73698 266648 73704
rect 274876 73756 274928 73762
rect 274876 73698 274928 73704
rect 266594 73248 266650 73257
rect 266594 73183 266650 73192
rect 266608 72402 266636 73183
rect 266596 72396 266648 72402
rect 266596 72338 266648 72344
rect 274692 72396 274744 72402
rect 274692 72338 274744 72344
rect 266686 72160 266742 72169
rect 266686 72095 266742 72104
rect 266594 71072 266650 71081
rect 266594 71007 266596 71016
rect 266648 71007 266650 71016
rect 266596 70978 266648 70984
rect 266700 70974 266728 72095
rect 272024 71036 272076 71042
rect 272024 70978 272076 70984
rect 266688 70968 266740 70974
rect 266688 70910 266740 70916
rect 266594 70120 266650 70129
rect 266594 70055 266650 70064
rect 266608 69614 266636 70055
rect 266596 69608 266648 69614
rect 266596 69550 266648 69556
rect 266594 69032 266650 69041
rect 266594 68967 266650 68976
rect 266608 68254 266636 68967
rect 266596 68248 266648 68254
rect 266596 68190 266648 68196
rect 266686 67944 266742 67953
rect 266686 67879 266742 67888
rect 266594 66992 266650 67001
rect 266594 66927 266650 66936
rect 266608 66826 266636 66927
rect 266700 66894 266728 67879
rect 267240 67568 267292 67574
rect 267240 67510 267292 67516
rect 266688 66888 266740 66894
rect 266688 66830 266740 66836
rect 266596 66820 266648 66826
rect 266596 66762 266648 66768
rect 266594 65904 266650 65913
rect 266594 65839 266650 65848
rect 266608 65466 266636 65839
rect 266596 65460 266648 65466
rect 266596 65402 266648 65408
rect 266594 64952 266650 64961
rect 266594 64887 266650 64896
rect 266608 64106 266636 64887
rect 266596 64100 266648 64106
rect 266596 64042 266648 64048
rect 266686 63864 266742 63873
rect 266686 63799 266742 63808
rect 266594 62776 266650 62785
rect 266594 62711 266596 62720
rect 266648 62711 266650 62720
rect 266596 62682 266648 62688
rect 266700 62678 266728 63799
rect 266688 62672 266740 62678
rect 266688 62614 266740 62620
rect 266594 61824 266650 61833
rect 266594 61759 266650 61768
rect 266608 61318 266636 61759
rect 266596 61312 266648 61318
rect 266596 61254 266648 61260
rect 266594 60736 266650 60745
rect 266594 60671 266650 60680
rect 266608 59958 266636 60671
rect 266596 59952 266648 59958
rect 266596 59894 266648 59900
rect 267252 55577 267280 67510
rect 272036 66758 272064 70978
rect 274704 68497 274732 72338
rect 274784 70968 274836 70974
rect 274784 70910 274836 70916
rect 274690 68488 274746 68497
rect 274690 68423 274746 68432
rect 274692 68248 274744 68254
rect 274692 68190 274744 68196
rect 272668 66888 272720 66894
rect 272668 66830 272720 66836
rect 272024 66752 272076 66758
rect 272024 66694 272076 66700
rect 272680 65398 272708 66830
rect 274232 66820 274284 66826
rect 274232 66762 274284 66768
rect 272668 65392 272720 65398
rect 272668 65334 272720 65340
rect 273404 64100 273456 64106
rect 273404 64042 273456 64048
rect 272852 62740 272904 62746
rect 272852 62682 272904 62688
rect 272760 61312 272812 61318
rect 272760 61254 272812 61260
rect 272668 59952 272720 59958
rect 272668 59894 272720 59900
rect 267330 59648 267386 59657
rect 267330 59583 267386 59592
rect 267344 58598 267372 59583
rect 267882 58696 267938 58705
rect 267882 58631 267884 58640
rect 267936 58631 267938 58640
rect 272116 58660 272168 58666
rect 267884 58602 267936 58608
rect 272116 58602 272168 58608
rect 267332 58592 267384 58598
rect 267332 58534 267384 58540
rect 267698 57608 267754 57617
rect 267698 57543 267754 57552
rect 267712 57442 267740 57543
rect 267700 57436 267752 57442
rect 267700 57378 267752 57384
rect 272128 57034 272156 58602
rect 272300 58592 272352 58598
rect 272300 58534 272352 58540
rect 272208 57436 272260 57442
rect 272208 57378 272260 57384
rect 272116 57028 272168 57034
rect 272116 56970 272168 56976
rect 267330 56656 267386 56665
rect 267330 56591 267386 56600
rect 267344 55810 267372 56591
rect 267332 55804 267384 55810
rect 267332 55746 267384 55752
rect 272116 55804 272168 55810
rect 272116 55746 272168 55752
rect 267238 55568 267294 55577
rect 267238 55503 267294 55512
rect 267882 54480 267938 54489
rect 267882 54415 267884 54424
rect 267936 54415 267938 54424
rect 267884 54386 267936 54392
rect 272128 54382 272156 55746
rect 272220 55742 272248 57378
rect 272312 57102 272340 58534
rect 272680 58530 272708 59894
rect 272772 59890 272800 61254
rect 272760 59884 272812 59890
rect 272760 59826 272812 59832
rect 272864 59822 272892 62682
rect 273416 62610 273444 64042
rect 274244 63193 274272 66762
rect 274704 64961 274732 68190
rect 274796 67681 274824 70910
rect 274888 69449 274916 73698
rect 285836 72402 285864 81314
rect 305064 73762 305092 83678
rect 311872 80170 311900 83814
rect 319140 80630 319168 83814
rect 318300 80624 318352 80630
rect 318300 80566 318352 80572
rect 319128 80624 319180 80630
rect 319128 80566 319180 80572
rect 311872 80142 312084 80170
rect 312056 76414 312084 80142
rect 312044 76408 312096 76414
rect 312044 76350 312096 76356
rect 304868 73756 304920 73762
rect 304868 73698 304920 73704
rect 305052 73756 305104 73762
rect 305052 73698 305104 73704
rect 304880 72402 304908 73698
rect 318312 72674 318340 80566
rect 321796 73756 321848 73762
rect 321796 73698 321848 73704
rect 311216 72668 311268 72674
rect 311216 72610 311268 72616
rect 318300 72668 318352 72674
rect 318300 72610 318352 72616
rect 284536 72396 284588 72402
rect 284536 72338 284588 72344
rect 285824 72396 285876 72402
rect 285824 72338 285876 72344
rect 297876 72396 297928 72402
rect 297876 72338 297928 72344
rect 304868 72396 304920 72402
rect 304868 72338 304920 72344
rect 284548 69820 284576 72338
rect 297888 69820 297916 72338
rect 311228 69820 311256 72610
rect 321244 70968 321296 70974
rect 321244 70910 321296 70916
rect 274968 69608 275020 69614
rect 274968 69550 275020 69556
rect 274874 69440 274930 69449
rect 274874 69375 274930 69384
rect 274782 67672 274838 67681
rect 274782 67607 274838 67616
rect 274876 66752 274928 66758
rect 274874 66720 274876 66729
rect 274928 66720 274930 66729
rect 274874 66655 274930 66664
rect 274980 65913 275008 69550
rect 317392 67630 317604 67658
rect 317392 66758 317420 67630
rect 317576 67574 317604 67630
rect 317564 67568 317616 67574
rect 317564 67510 317616 67516
rect 317380 66752 317432 66758
rect 321256 66729 321284 70910
rect 321702 69440 321758 69449
rect 321808 69426 321836 73698
rect 321758 69398 321836 69426
rect 321702 69375 321758 69384
rect 321612 69132 321664 69138
rect 321612 69074 321664 69080
rect 321624 68497 321652 69074
rect 321610 68488 321666 68497
rect 321610 68423 321666 68432
rect 321610 67672 321666 67681
rect 321610 67607 321666 67616
rect 321624 67098 321652 67607
rect 321612 67092 321664 67098
rect 321612 67034 321664 67040
rect 317380 66694 317432 66700
rect 321242 66720 321298 66729
rect 321242 66655 321298 66664
rect 321612 66004 321664 66010
rect 321612 65946 321664 65952
rect 321624 65913 321652 65946
rect 274966 65904 275022 65913
rect 274966 65839 275022 65848
rect 321610 65904 321666 65913
rect 321610 65839 321666 65848
rect 274784 65460 274836 65466
rect 274784 65402 274836 65408
rect 274690 64952 274746 64961
rect 274690 64887 274746 64896
rect 274230 63184 274286 63193
rect 274230 63119 274286 63128
rect 273404 62604 273456 62610
rect 273404 62546 273456 62552
rect 274796 62377 274824 65402
rect 274876 65392 274928 65398
rect 274876 65334 274928 65340
rect 274888 64145 274916 65334
rect 321610 64952 321666 64961
rect 321610 64887 321666 64896
rect 321624 64650 321652 64887
rect 321612 64644 321664 64650
rect 321612 64586 321664 64592
rect 321612 64168 321664 64174
rect 274874 64136 274930 64145
rect 274874 64071 274930 64080
rect 321610 64136 321612 64145
rect 321664 64136 321666 64145
rect 321610 64071 321666 64080
rect 320508 63692 320560 63698
rect 320508 63634 320560 63640
rect 320520 62785 320548 63634
rect 320506 62776 320562 62785
rect 320506 62711 320562 62720
rect 274876 62672 274928 62678
rect 274876 62614 274928 62620
rect 274782 62368 274838 62377
rect 274782 62303 274838 62312
rect 274888 60473 274916 62614
rect 274968 62604 275020 62610
rect 274968 62546 275020 62552
rect 321060 62604 321112 62610
rect 321060 62546 321112 62552
rect 274980 61425 275008 62546
rect 318390 61824 318446 61833
rect 318390 61759 318446 61768
rect 318404 61425 318432 61759
rect 320692 61584 320744 61590
rect 320690 61552 320692 61561
rect 320744 61552 320746 61561
rect 320690 61487 320746 61496
rect 321072 61425 321100 62546
rect 274966 61416 275022 61425
rect 274966 61351 275022 61360
rect 318390 61416 318446 61425
rect 318390 61351 318446 61360
rect 321058 61416 321114 61425
rect 321058 61351 321114 61360
rect 274874 60464 274930 60473
rect 274874 60399 274930 60408
rect 321060 60292 321112 60298
rect 321060 60234 321112 60240
rect 321072 59929 321100 60234
rect 321058 59920 321114 59929
rect 275428 59884 275480 59890
rect 321058 59855 321114 59864
rect 275428 59826 275480 59832
rect 272852 59816 272904 59822
rect 272852 59758 272904 59764
rect 275440 58705 275468 59826
rect 275704 59816 275756 59822
rect 275704 59758 275756 59764
rect 275716 59657 275744 59758
rect 275702 59648 275758 59657
rect 275702 59583 275758 59592
rect 320506 59648 320562 59657
rect 320506 59583 320562 59592
rect 320520 58734 320548 59583
rect 320508 58728 320560 58734
rect 275426 58696 275482 58705
rect 275426 58631 275482 58640
rect 320414 58696 320470 58705
rect 320508 58670 320560 58676
rect 320414 58631 320470 58640
rect 320428 58598 320456 58631
rect 320416 58592 320468 58598
rect 320416 58534 320468 58540
rect 272668 58524 272720 58530
rect 272668 58466 272720 58472
rect 275704 58524 275756 58530
rect 275704 58466 275756 58472
rect 275716 57889 275744 58466
rect 275702 57880 275758 57889
rect 275702 57815 275758 57824
rect 320414 57880 320470 57889
rect 320414 57815 320416 57824
rect 320468 57815 320470 57824
rect 320416 57786 320468 57792
rect 317564 57164 317616 57170
rect 317564 57106 317616 57112
rect 272300 57096 272352 57102
rect 272300 57038 272352 57044
rect 275704 57096 275756 57102
rect 275704 57038 275756 57044
rect 275244 57028 275296 57034
rect 275244 56970 275296 56976
rect 275256 56121 275284 56970
rect 275716 56937 275744 57038
rect 275702 56928 275758 56937
rect 275702 56863 275758 56872
rect 275242 56112 275298 56121
rect 275242 56047 275298 56056
rect 272208 55736 272260 55742
rect 272208 55678 272260 55684
rect 275428 55736 275480 55742
rect 275428 55678 275480 55684
rect 275440 55169 275468 55678
rect 275426 55160 275482 55169
rect 275426 55095 275482 55104
rect 317576 55062 317604 57106
rect 320506 56928 320562 56937
rect 320506 56863 320562 56872
rect 320416 56552 320468 56558
rect 320416 56494 320468 56500
rect 320428 56121 320456 56494
rect 320520 56354 320548 56863
rect 320508 56348 320560 56354
rect 320508 56290 320560 56296
rect 320414 56112 320470 56121
rect 320414 56047 320470 56056
rect 320416 55668 320468 55674
rect 320416 55610 320468 55616
rect 320428 55169 320456 55610
rect 320414 55160 320470 55169
rect 320414 55095 320470 55104
rect 317564 55056 317616 55062
rect 317564 54998 317616 55004
rect 272116 54376 272168 54382
rect 275704 54376 275756 54382
rect 272116 54318 272168 54324
rect 275702 54344 275704 54353
rect 275756 54344 275758 54353
rect 275702 54279 275758 54288
rect 320414 54344 320470 54353
rect 320414 54279 320470 54288
rect 320428 54246 320456 54279
rect 320416 54240 320468 54246
rect 320416 54182 320468 54188
rect 311584 54172 311636 54178
rect 311584 54114 311636 54120
rect 267884 53696 267936 53702
rect 267884 53638 267936 53644
rect 267896 53537 267924 53638
rect 267882 53528 267938 53537
rect 267882 53463 267938 53472
rect 267884 53016 267936 53022
rect 267884 52958 267936 52964
rect 267896 52449 267924 52958
rect 267882 52440 267938 52449
rect 267882 52375 267938 52384
rect 279028 51594 279056 53908
rect 279016 51588 279068 51594
rect 279016 51530 279068 51536
rect 281328 51361 281356 53908
rect 267514 51352 267570 51361
rect 267514 51287 267570 51296
rect 281314 51352 281370 51361
rect 281314 51287 281370 51296
rect 266778 50400 266834 50409
rect 267528 50370 267556 51287
rect 280304 50908 280356 50914
rect 280304 50850 280356 50856
rect 266778 50335 266834 50344
rect 267516 50364 267568 50370
rect 266792 50302 266820 50335
rect 267516 50306 267568 50312
rect 266780 50296 266832 50302
rect 266780 50238 266832 50244
rect 276164 49548 276216 49554
rect 276164 49490 276216 49496
rect 267882 49312 267938 49321
rect 267882 49247 267938 49256
rect 267896 48942 267924 49247
rect 267884 48936 267936 48942
rect 267884 48878 267936 48884
rect 267882 48360 267938 48369
rect 267882 48295 267938 48304
rect 267896 47514 267924 48295
rect 276072 48188 276124 48194
rect 276072 48130 276124 48136
rect 276084 47961 276112 48130
rect 275794 47952 275850 47961
rect 275794 47887 275850 47896
rect 276070 47952 276126 47961
rect 276070 47887 276126 47896
rect 267884 47508 267936 47514
rect 267884 47450 267936 47456
rect 275520 45876 275572 45882
rect 275520 45818 275572 45824
rect 275532 23345 275560 45818
rect 275808 28105 275836 47887
rect 275980 46760 276032 46766
rect 275980 46702 276032 46708
rect 275992 46601 276020 46702
rect 275978 46592 276034 46601
rect 275978 46527 276034 46536
rect 275888 45332 275940 45338
rect 275888 45274 275940 45280
rect 275900 33681 275928 45274
rect 275886 33672 275942 33681
rect 275886 33607 275942 33616
rect 275992 30825 276020 46527
rect 276176 45882 276204 49490
rect 276164 45876 276216 45882
rect 276164 45818 276216 45824
rect 276072 45400 276124 45406
rect 276072 45342 276124 45348
rect 276084 44794 276112 45342
rect 276072 44788 276124 44794
rect 276072 44730 276124 44736
rect 275978 30816 276034 30825
rect 275978 30751 276034 30760
rect 275794 28096 275850 28105
rect 275794 28031 275850 28040
rect 276084 26065 276112 44730
rect 280316 37382 280344 50850
rect 283720 48097 283748 53908
rect 284444 50976 284496 50982
rect 284444 50918 284496 50924
rect 283706 48088 283762 48097
rect 283706 48023 283762 48032
rect 284350 48088 284406 48097
rect 284350 48023 284406 48032
rect 281592 47508 281644 47514
rect 281592 47450 281644 47456
rect 279108 37376 279160 37382
rect 279108 37318 279160 37324
rect 280304 37376 280356 37382
rect 280304 37318 280356 37324
rect 279120 34732 279148 37318
rect 281604 34732 281632 47450
rect 284364 45814 284392 48023
rect 284352 45808 284404 45814
rect 284352 45750 284404 45756
rect 284456 34746 284484 50918
rect 286020 47417 286048 53908
rect 288412 49554 288440 53908
rect 289964 51044 290016 51050
rect 289964 50986 290016 50992
rect 288400 49548 288452 49554
rect 288400 49490 288452 49496
rect 286560 48936 286612 48942
rect 286560 48878 286612 48884
rect 286006 47408 286062 47417
rect 286006 47343 286008 47352
rect 286060 47343 286062 47352
rect 286008 47314 286060 47320
rect 286020 47283 286048 47314
rect 284102 34718 284484 34746
rect 286572 34732 286600 48878
rect 289976 37790 290004 50986
rect 290712 45406 290740 53908
rect 291528 50296 291580 50302
rect 291528 50238 291580 50244
rect 290700 45400 290752 45406
rect 290700 45342 290752 45348
rect 289044 37784 289096 37790
rect 289044 37726 289096 37732
rect 289964 37784 290016 37790
rect 289964 37726 290016 37732
rect 289056 34732 289084 37726
rect 291540 34732 291568 50238
rect 293104 48194 293132 53908
rect 294104 51112 294156 51118
rect 294104 51054 294156 51060
rect 293092 48188 293144 48194
rect 293092 48130 293144 48136
rect 294116 34732 294144 51054
rect 295496 47446 295524 53908
rect 297810 53894 298284 53922
rect 296588 50364 296640 50370
rect 296588 50306 296640 50312
rect 295484 47440 295536 47446
rect 295484 47382 295536 47388
rect 295496 46766 295524 47382
rect 295484 46760 295536 46766
rect 295484 46702 295536 46708
rect 296600 34732 296628 50306
rect 298256 46086 298284 53894
rect 299624 51180 299676 51186
rect 299624 51122 299676 51128
rect 298244 46080 298296 46086
rect 298244 46022 298296 46028
rect 299636 34610 299664 51122
rect 300188 50914 300216 53908
rect 301646 53120 301702 53129
rect 301646 53055 301702 53064
rect 301660 53022 301688 53055
rect 301648 53016 301700 53022
rect 301648 52958 301700 52964
rect 302488 50982 302516 53908
rect 304880 51050 304908 53908
rect 306616 53696 306668 53702
rect 306616 53638 306668 53644
rect 306628 53129 306656 53638
rect 306614 53120 306670 53129
rect 306614 53055 306670 53064
rect 307272 51118 307300 53908
rect 309572 51186 309600 53908
rect 309560 51180 309612 51186
rect 309560 51122 309612 51128
rect 307260 51112 307312 51118
rect 307260 51054 307312 51060
rect 304868 51044 304920 51050
rect 304868 50986 304920 50992
rect 302476 50976 302528 50982
rect 302476 50918 302528 50924
rect 300176 50908 300228 50914
rect 300176 50850 300228 50856
rect 305144 50908 305196 50914
rect 305144 50850 305196 50856
rect 305156 37790 305184 50850
rect 306614 47408 306670 47417
rect 306614 47343 306670 47352
rect 304040 37784 304092 37790
rect 301554 37752 301610 37761
rect 304040 37726 304092 37732
rect 305144 37784 305196 37790
rect 305144 37726 305196 37732
rect 301554 37687 301610 37696
rect 301568 34732 301596 37687
rect 304052 34732 304080 37726
rect 306628 34732 306656 47343
rect 309100 36764 309152 36770
rect 309100 36706 309152 36712
rect 309112 34732 309140 36706
rect 311596 34732 311624 54114
rect 311964 50914 311992 53908
rect 314264 51526 314292 53908
rect 316656 51526 316684 53908
rect 312780 51520 312832 51526
rect 312780 51462 312832 51468
rect 314252 51520 314304 51526
rect 314252 51462 314304 51468
rect 314804 51520 314856 51526
rect 314804 51462 314856 51468
rect 316644 51520 316696 51526
rect 316644 51462 316696 51468
rect 311952 50908 312004 50914
rect 311952 50850 312004 50856
rect 312792 36770 312820 51462
rect 314816 37178 314844 51462
rect 317472 46148 317524 46154
rect 317472 46090 317524 46096
rect 317484 44862 317512 46090
rect 322544 45950 322572 224114
rect 323820 222880 323872 222886
rect 323820 222822 323872 222828
rect 322624 222812 322676 222818
rect 322624 222754 322676 222760
rect 322636 131290 322664 222754
rect 322808 221384 322860 221390
rect 322808 221326 322860 221332
rect 322716 220500 322768 220506
rect 322716 220442 322768 220448
rect 322728 139858 322756 220442
rect 322820 145434 322848 221326
rect 323176 152500 323228 152506
rect 323176 152442 323228 152448
rect 323188 150942 323216 152442
rect 323268 151412 323320 151418
rect 323268 151354 323320 151360
rect 323176 150936 323228 150942
rect 323176 150878 323228 150884
rect 323176 149644 323228 149650
rect 323176 149586 323228 149592
rect 323188 148222 323216 149586
rect 323280 149582 323308 151354
rect 323268 149576 323320 149582
rect 323268 149518 323320 149524
rect 323176 148216 323228 148222
rect 323176 148158 323228 148164
rect 322808 145428 322860 145434
rect 322808 145370 322860 145376
rect 322716 139852 322768 139858
rect 322716 139794 322768 139800
rect 322624 131284 322676 131290
rect 322624 131226 322676 131232
rect 323832 51594 323860 222822
rect 324568 198785 324596 292143
rect 325212 262802 325240 310911
rect 325304 292217 325332 314418
rect 325384 309716 325436 309722
rect 325384 309658 325436 309664
rect 325290 292208 325346 292217
rect 325290 292143 325346 292152
rect 325290 285952 325346 285961
rect 325290 285887 325346 285896
rect 325200 262796 325252 262802
rect 325200 262738 325252 262744
rect 324648 261436 324700 261442
rect 324648 261378 324700 261384
rect 324660 258586 324688 261378
rect 324648 258580 324700 258586
rect 324648 258522 324700 258528
rect 325200 238588 325252 238594
rect 325200 238530 325252 238536
rect 324832 235936 324884 235942
rect 324832 235878 324884 235884
rect 324646 234408 324702 234417
rect 324646 234343 324702 234352
rect 324660 229686 324688 234343
rect 324844 231046 324872 235878
rect 324924 234440 324976 234446
rect 324924 234382 324976 234388
rect 324936 233834 324964 234382
rect 324924 233828 324976 233834
rect 324924 233770 324976 233776
rect 324832 231040 324884 231046
rect 324832 230982 324884 230988
rect 324648 229680 324700 229686
rect 324648 229622 324700 229628
rect 324936 229498 324964 233770
rect 324660 229470 324964 229498
rect 324660 223265 324688 229470
rect 324738 226384 324794 226393
rect 324738 226319 324740 226328
rect 324792 226319 324794 226328
rect 324740 226290 324792 226296
rect 325212 224246 325240 238530
rect 324924 224240 324976 224246
rect 324924 224182 324976 224188
rect 325200 224240 325252 224246
rect 325200 224182 325252 224188
rect 324646 223256 324702 223265
rect 324646 223191 324702 223200
rect 324936 213881 324964 224182
rect 325200 221452 325252 221458
rect 325200 221394 325252 221400
rect 324922 213872 324978 213881
rect 324922 213807 324978 213816
rect 324554 198776 324610 198785
rect 324554 198711 324610 198720
rect 324556 188948 324608 188954
rect 324556 188890 324608 188896
rect 324568 188857 324596 188890
rect 324554 188848 324610 188857
rect 324554 188783 324610 188792
rect 324556 179904 324608 179910
rect 324556 179846 324608 179852
rect 324568 179473 324596 179846
rect 324554 179464 324610 179473
rect 324554 179399 324610 179408
rect 324556 166236 324608 166242
rect 324556 166178 324608 166184
rect 324568 163386 324596 166178
rect 324556 163380 324608 163386
rect 324556 163322 324608 163328
rect 324556 142096 324608 142102
rect 324556 142038 324608 142044
rect 324568 135846 324596 142038
rect 325108 140600 325160 140606
rect 325108 140542 325160 140548
rect 324832 137880 324884 137886
rect 324832 137822 324884 137828
rect 324556 135840 324608 135846
rect 324556 135782 324608 135788
rect 324568 132417 324596 135782
rect 324648 135092 324700 135098
rect 324648 135034 324700 135040
rect 324660 134486 324688 135034
rect 324648 134480 324700 134486
rect 324648 134422 324700 134428
rect 324660 132666 324688 134422
rect 324660 132638 324780 132666
rect 324646 132544 324702 132553
rect 324646 132479 324702 132488
rect 324554 132408 324610 132417
rect 324554 132343 324610 132352
rect 324556 132236 324608 132242
rect 324556 132178 324608 132184
rect 324568 120018 324596 132178
rect 324660 130338 324688 132479
rect 324752 132242 324780 132638
rect 324740 132236 324792 132242
rect 324740 132178 324792 132184
rect 324844 131766 324872 137822
rect 324832 131760 324884 131766
rect 324832 131702 324884 131708
rect 325120 131698 325148 140542
rect 325108 131692 325160 131698
rect 325108 131634 325160 131640
rect 324740 130400 324792 130406
rect 324740 130342 324792 130348
rect 324648 130332 324700 130338
rect 324648 130274 324700 130280
rect 324660 126025 324688 130274
rect 324646 126016 324702 126025
rect 324646 125951 324702 125960
rect 324752 123305 324780 130342
rect 325120 129833 325148 131634
rect 325106 129824 325162 129833
rect 325106 129759 325162 129768
rect 324738 123296 324794 123305
rect 324738 123231 324794 123240
rect 324476 119990 324596 120018
rect 324476 119746 324504 119990
rect 324556 119928 324608 119934
rect 324554 119896 324556 119905
rect 324608 119896 324610 119905
rect 324554 119831 324610 119840
rect 324476 119718 324596 119746
rect 324568 117321 324596 119718
rect 324554 117312 324610 117321
rect 324554 117247 324610 117256
rect 325212 98553 325240 221394
rect 325304 220642 325332 285887
rect 325396 279705 325424 309658
rect 325488 305545 325516 319382
rect 325474 305536 325530 305545
rect 325474 305471 325530 305480
rect 325580 305409 325608 319994
rect 325566 305400 325622 305409
rect 325566 305335 325622 305344
rect 325672 301601 325700 320742
rect 325764 307857 325792 323462
rect 325844 320188 325896 320194
rect 325844 320130 325896 320136
rect 325856 319446 325884 320130
rect 325844 319440 325896 319446
rect 325844 319382 325896 319388
rect 325844 319304 325896 319310
rect 325844 319246 325896 319252
rect 325856 314113 325884 319246
rect 325842 314104 325898 314113
rect 325842 314039 325898 314048
rect 325750 307848 325806 307857
rect 325750 307783 325806 307792
rect 325658 301592 325714 301601
rect 325658 301527 325714 301536
rect 325476 295912 325528 295918
rect 325476 295854 325528 295860
rect 325382 279696 325438 279705
rect 325382 279631 325438 279640
rect 325488 276577 325516 295854
rect 325568 283536 325620 283542
rect 325568 283478 325620 283484
rect 325474 276568 325530 276577
rect 325474 276503 325530 276512
rect 325580 273449 325608 283478
rect 325844 282856 325896 282862
rect 325842 282824 325844 282833
rect 325896 282824 325898 282833
rect 325842 282759 325898 282768
rect 325566 273440 325622 273449
rect 325566 273375 325622 273384
rect 325844 262796 325896 262802
rect 325844 262738 325896 262744
rect 325856 239721 325884 262738
rect 325842 239712 325898 239721
rect 325842 239647 325898 239656
rect 325384 235868 325436 235874
rect 325384 235810 325436 235816
rect 325396 227034 325424 235810
rect 325752 231040 325804 231046
rect 325752 230982 325804 230988
rect 325476 229680 325528 229686
rect 325476 229622 325528 229628
rect 325384 227028 325436 227034
rect 325384 226970 325436 226976
rect 325292 220636 325344 220642
rect 325292 220578 325344 220584
rect 325384 220568 325436 220574
rect 325384 220510 325436 220516
rect 325292 215876 325344 215882
rect 325292 215818 325344 215824
rect 325304 185729 325332 215818
rect 325396 191985 325424 220510
rect 325488 207625 325516 229622
rect 325660 227028 325712 227034
rect 325660 226970 325712 226976
rect 325568 222948 325620 222954
rect 325568 222890 325620 222896
rect 325474 207616 325530 207625
rect 325474 207551 325530 207560
rect 325580 204497 325608 222890
rect 325672 210753 325700 226970
rect 325764 220137 325792 230982
rect 325856 224314 325884 239647
rect 326592 232270 326620 326862
rect 330088 282862 330116 329838
rect 331468 320534 331496 329838
rect 331456 320528 331508 320534
rect 331456 320470 331508 320476
rect 332848 320262 332876 329852
rect 333676 326586 333704 329852
rect 334320 329838 334426 329866
rect 334216 326852 334268 326858
rect 334216 326794 334268 326800
rect 332928 326580 332980 326586
rect 332928 326522 332980 326528
rect 333664 326580 333716 326586
rect 333664 326522 333716 326528
rect 332940 320602 332968 326522
rect 332928 320596 332980 320602
rect 332928 320538 332980 320544
rect 332836 320256 332888 320262
rect 332836 320198 332888 320204
rect 334228 320058 334256 326794
rect 334320 320126 334348 329838
rect 335240 326858 335268 329852
rect 335608 329838 336082 329866
rect 335228 326852 335280 326858
rect 335228 326794 335280 326800
rect 335608 320330 335636 329838
rect 336804 326926 336832 329852
rect 336988 329838 337646 329866
rect 335688 326920 335740 326926
rect 335688 326862 335740 326868
rect 336792 326920 336844 326926
rect 336792 326862 336844 326868
rect 335596 320324 335648 320330
rect 335596 320266 335648 320272
rect 334308 320120 334360 320126
rect 334308 320062 334360 320068
rect 334216 320052 334268 320058
rect 334216 319994 334268 320000
rect 335700 319990 335728 326862
rect 336988 320398 337016 329838
rect 337160 327600 337212 327606
rect 337160 327542 337212 327548
rect 337068 326512 337120 326518
rect 337068 326454 337120 326460
rect 336976 320392 337028 320398
rect 336976 320334 337028 320340
rect 335688 319984 335740 319990
rect 335688 319926 335740 319932
rect 337080 316810 337108 326454
rect 337172 320670 337200 327542
rect 337160 320664 337212 320670
rect 337160 320606 337212 320612
rect 337528 320664 337580 320670
rect 337528 320606 337580 320612
rect 337540 316810 337568 320606
rect 338460 320466 338488 329852
rect 339196 327441 339224 329852
rect 340024 327441 340052 329852
rect 339182 327432 339238 327441
rect 340010 327432 340066 327441
rect 339182 327367 339238 327376
rect 339644 327396 339696 327402
rect 340010 327367 340066 327376
rect 339644 327338 339696 327344
rect 338540 326920 338592 326926
rect 338540 326862 338592 326868
rect 338448 320460 338500 320466
rect 338448 320402 338500 320408
rect 338552 319786 338580 326862
rect 339368 326852 339420 326858
rect 339368 326794 339420 326800
rect 338540 319780 338592 319786
rect 338540 319722 338592 319728
rect 338724 319644 338776 319650
rect 338724 319586 338776 319592
rect 338736 316810 338764 319586
rect 339380 316810 339408 326794
rect 339460 319780 339512 319786
rect 339460 319722 339512 319728
rect 337080 316782 337232 316810
rect 337540 316782 337784 316810
rect 338428 316782 338764 316810
rect 339072 316782 339408 316810
rect 339472 316810 339500 319722
rect 339656 319650 339684 327338
rect 339920 327056 339972 327062
rect 339920 326998 339972 327004
rect 339932 320670 339960 326998
rect 340852 326722 340880 329852
rect 341300 327532 341352 327538
rect 341300 327474 341352 327480
rect 341024 327464 341076 327470
rect 341024 327406 341076 327412
rect 340840 326716 340892 326722
rect 340840 326658 340892 326664
rect 339920 320664 339972 320670
rect 339920 320606 339972 320612
rect 340564 320664 340616 320670
rect 340564 320606 340616 320612
rect 340472 320528 340524 320534
rect 340472 320470 340524 320476
rect 339644 319644 339696 319650
rect 339644 319586 339696 319592
rect 340484 316810 340512 320470
rect 339472 316782 339624 316810
rect 340268 316782 340512 316810
rect 340576 316810 340604 320606
rect 341036 320534 341064 327406
rect 341208 327124 341260 327130
rect 341208 327066 341260 327072
rect 341024 320528 341076 320534
rect 341024 320470 341076 320476
rect 341220 319514 341248 327066
rect 341208 319508 341260 319514
rect 341208 319450 341260 319456
rect 341312 316810 341340 327474
rect 341588 326654 341616 329852
rect 342416 327334 342444 329852
rect 342404 327328 342456 327334
rect 342404 327270 342456 327276
rect 343244 326790 343272 329852
rect 343232 326784 343284 326790
rect 343232 326726 343284 326732
rect 341576 326648 341628 326654
rect 341576 326590 341628 326596
rect 343980 326586 344008 329852
rect 344808 327198 344836 329852
rect 345256 327668 345308 327674
rect 345256 327610 345308 327616
rect 344796 327192 344848 327198
rect 344796 327134 344848 327140
rect 343968 326580 344020 326586
rect 343968 326522 344020 326528
rect 343968 324880 344020 324886
rect 343968 324822 344020 324828
rect 343876 322840 343928 322846
rect 343876 322782 343928 322788
rect 343888 322234 343916 322782
rect 343876 322228 343928 322234
rect 343876 322170 343928 322176
rect 342496 322092 342548 322098
rect 342496 322034 342548 322040
rect 342508 320806 342536 322034
rect 342496 320800 342548 320806
rect 342496 320742 342548 320748
rect 342956 320800 343008 320806
rect 342956 320742 343008 320748
rect 341760 319508 341812 319514
rect 341760 319450 341812 319456
rect 341772 316810 341800 319450
rect 342496 319440 342548 319446
rect 342496 319382 342548 319388
rect 342508 316810 342536 319382
rect 342968 316810 342996 320742
rect 343980 317082 344008 324822
rect 344796 324132 344848 324138
rect 344796 324074 344848 324080
rect 344808 323526 344836 324074
rect 344796 323520 344848 323526
rect 344796 323462 344848 323468
rect 343934 317054 344008 317082
rect 340576 316782 340912 316810
rect 341312 316782 341464 316810
rect 341772 316782 342108 316810
rect 342508 316782 342752 316810
rect 342968 316782 343304 316810
rect 343934 316796 343962 317054
rect 344808 316810 344836 323462
rect 345164 322840 345216 322846
rect 345164 322782 345216 322788
rect 344592 316782 344836 316810
rect 345176 316810 345204 322782
rect 345268 322098 345296 327610
rect 345636 327266 345664 329852
rect 346096 329838 346478 329866
rect 346096 327674 346124 329838
rect 346084 327668 346136 327674
rect 346084 327610 346136 327616
rect 345624 327260 345676 327266
rect 345624 327202 345676 327208
rect 347200 324886 347228 329852
rect 348042 329838 348148 329866
rect 348016 325220 348068 325226
rect 348016 325162 348068 325168
rect 347188 324880 347240 324886
rect 347188 324822 347240 324828
rect 348028 322846 348056 325162
rect 348120 324138 348148 329838
rect 348488 329838 348870 329866
rect 349408 329838 349606 329866
rect 349684 329838 350434 329866
rect 348488 325226 348516 329838
rect 348476 325220 348528 325226
rect 348476 325162 348528 325168
rect 348108 324132 348160 324138
rect 348108 324074 348160 324080
rect 348016 322840 348068 322846
rect 348016 322782 348068 322788
rect 347004 322160 347056 322166
rect 347004 322102 347056 322108
rect 345256 322092 345308 322098
rect 345256 322034 345308 322040
rect 346452 320732 346504 320738
rect 346452 320674 346504 320680
rect 345716 319372 345768 319378
rect 345716 319314 345768 319320
rect 345728 316810 345756 319314
rect 346464 317082 346492 320674
rect 346418 317054 346492 317082
rect 345176 316782 345236 316810
rect 345728 316782 345788 316810
rect 346418 316796 346446 317054
rect 347016 316674 347044 322102
rect 348568 320596 348620 320602
rect 348568 320538 348620 320544
rect 348016 320256 348068 320262
rect 348016 320198 348068 320204
rect 347280 320188 347332 320194
rect 347280 320130 347332 320136
rect 347292 316810 347320 320130
rect 348028 316810 348056 320198
rect 348580 316810 348608 320538
rect 349408 320210 349436 329838
rect 349684 327418 349712 329838
rect 349500 327390 349712 327418
rect 349500 320738 349528 327390
rect 351248 322166 351276 329852
rect 351984 326518 352012 329852
rect 352812 327606 352840 329852
rect 352800 327600 352852 327606
rect 352800 327542 352852 327548
rect 353640 327402 353668 329852
rect 353628 327396 353680 327402
rect 353628 327338 353680 327344
rect 354376 326858 354404 329852
rect 355204 326926 355232 329852
rect 356032 327470 356060 329852
rect 356020 327464 356072 327470
rect 356020 327406 356072 327412
rect 355560 327328 355612 327334
rect 355560 327270 355612 327276
rect 355192 326920 355244 326926
rect 355192 326862 355244 326868
rect 354364 326852 354416 326858
rect 354364 326794 354416 326800
rect 352800 326716 352852 326722
rect 352800 326658 352852 326664
rect 351972 326512 352024 326518
rect 351972 326454 352024 326460
rect 351236 322160 351288 322166
rect 351236 322102 351288 322108
rect 349488 320732 349540 320738
rect 349488 320674 349540 320680
rect 352812 320602 352840 326658
rect 354180 326648 354232 326654
rect 354180 326590 354232 326596
rect 352800 320596 352852 320602
rect 352800 320538 352852 320544
rect 352248 320528 352300 320534
rect 352248 320470 352300 320476
rect 352892 320528 352944 320534
rect 352892 320470 352944 320476
rect 351604 320460 351656 320466
rect 351604 320402 351656 320408
rect 350408 320392 350460 320398
rect 350408 320334 350460 320340
rect 349408 320182 349528 320210
rect 349396 320120 349448 320126
rect 349396 320062 349448 320068
rect 349408 316810 349436 320062
rect 349500 319990 349528 320182
rect 349764 320052 349816 320058
rect 349764 319994 349816 320000
rect 349488 319984 349540 319990
rect 349488 319926 349540 319932
rect 349500 319378 349528 319926
rect 349488 319372 349540 319378
rect 349488 319314 349540 319320
rect 349776 316810 349804 319994
rect 350420 316810 350448 320334
rect 350960 320324 351012 320330
rect 350960 320266 351012 320272
rect 350972 316810 351000 320266
rect 351616 316810 351644 320402
rect 352260 316810 352288 320470
rect 347292 316782 347628 316810
rect 348028 316782 348272 316810
rect 348580 316782 348916 316810
rect 349408 316782 349468 316810
rect 349776 316782 350112 316810
rect 350420 316782 350756 316810
rect 350972 316782 351308 316810
rect 351616 316782 351952 316810
rect 352260 316782 352596 316810
rect 347016 316646 347076 316674
rect 352904 316590 352932 320470
rect 352892 316584 352944 316590
rect 352892 316526 352944 316532
rect 334214 309752 334270 309761
rect 334214 309687 334216 309696
rect 334268 309687 334270 309696
rect 334216 309658 334268 309664
rect 352892 306996 352944 307002
rect 352892 306938 352944 306944
rect 352904 301494 352932 306938
rect 352892 301488 352944 301494
rect 352892 301430 352944 301436
rect 352800 301352 352852 301358
rect 352800 301294 352852 301300
rect 352812 297249 352840 301294
rect 352798 297240 352854 297249
rect 352798 297175 352854 297184
rect 353994 297240 354050 297249
rect 353994 297175 354050 297184
rect 334214 296288 334270 296297
rect 334214 296223 334270 296232
rect 334228 295918 334256 296223
rect 334216 295912 334268 295918
rect 334216 295854 334268 295860
rect 353536 295844 353588 295850
rect 353536 295786 353588 295792
rect 353548 295170 353576 295786
rect 353536 295164 353588 295170
rect 353536 295106 353588 295112
rect 334214 283640 334270 283649
rect 334214 283575 334270 283584
rect 334228 283542 334256 283575
rect 334216 283536 334268 283542
rect 334216 283478 334268 283484
rect 330076 282856 330128 282862
rect 330076 282798 330128 282804
rect 328420 264088 328472 264094
rect 328420 264030 328472 264036
rect 328432 263521 328460 264030
rect 330088 263906 330116 282798
rect 352984 279388 353036 279394
rect 352984 279330 353036 279336
rect 337324 276934 337660 276962
rect 336884 274832 336936 274838
rect 336884 274774 336936 274780
rect 334124 274764 334176 274770
rect 334124 274706 334176 274712
rect 332744 274628 332796 274634
rect 332744 274570 332796 274576
rect 330088 263878 330852 263906
rect 330824 263634 330852 263878
rect 332756 263770 332784 274570
rect 334136 265590 334164 274706
rect 335412 274696 335464 274702
rect 335412 274638 335464 274644
rect 335424 265590 335452 274638
rect 335504 274560 335556 274566
rect 335504 274502 335556 274508
rect 333388 265584 333440 265590
rect 333388 265526 333440 265532
rect 334124 265584 334176 265590
rect 334124 265526 334176 265532
rect 334400 265584 334452 265590
rect 334400 265526 334452 265532
rect 335412 265584 335464 265590
rect 335412 265526 335464 265532
rect 332402 263742 332784 263770
rect 333400 263756 333428 265526
rect 334412 263756 334440 265526
rect 335516 263756 335544 274502
rect 336896 263770 336924 274774
rect 337632 273954 337660 276934
rect 338138 276690 338166 276948
rect 338980 276934 339316 276962
rect 339808 276934 340144 276962
rect 340636 276934 340972 276962
rect 341464 276934 341800 276962
rect 342292 276934 342444 276962
rect 343212 276934 343548 276962
rect 344040 276934 344376 276962
rect 344868 276934 345204 276962
rect 338138 276662 338212 276690
rect 338184 274090 338212 276662
rect 338264 275036 338316 275042
rect 338264 274978 338316 274984
rect 338172 274084 338224 274090
rect 338172 274026 338224 274032
rect 337620 273948 337672 273954
rect 337620 273890 337672 273896
rect 338276 263906 338304 274978
rect 339288 274022 339316 276934
rect 339644 274968 339696 274974
rect 339644 274910 339696 274916
rect 339276 274016 339328 274022
rect 339276 273958 339328 273964
rect 338540 266196 338592 266202
rect 338540 266138 338592 266144
rect 337908 263878 338304 263906
rect 337908 263770 337936 263878
rect 336542 263742 336924 263770
rect 337554 263742 337936 263770
rect 338552 263756 338580 266138
rect 339656 263756 339684 274910
rect 340116 273886 340144 276934
rect 340104 273880 340156 273886
rect 340104 273822 340156 273828
rect 340944 273818 340972 276934
rect 341024 274900 341076 274906
rect 341024 274842 341076 274848
rect 340932 273812 340984 273818
rect 340932 273754 340984 273760
rect 341036 263770 341064 274842
rect 341772 274566 341800 276934
rect 342416 274702 342444 276934
rect 343520 274770 343548 276934
rect 343508 274764 343560 274770
rect 343508 274706 343560 274712
rect 342404 274696 342456 274702
rect 342404 274638 342456 274644
rect 344348 274634 344376 276934
rect 344336 274628 344388 274634
rect 344336 274570 344388 274576
rect 341760 274560 341812 274566
rect 341760 274502 341812 274508
rect 345176 274498 345204 276934
rect 345360 276934 345696 276962
rect 346188 276934 346524 276962
rect 347016 276934 347352 276962
rect 348028 276934 348272 276962
rect 348764 276934 349100 276962
rect 349592 276934 349928 276962
rect 350420 276934 350756 276962
rect 351248 276934 351584 276962
rect 352168 276934 352412 276962
rect 345164 274492 345216 274498
rect 345164 274434 345216 274440
rect 345360 274430 345388 276934
rect 346188 274838 346216 276934
rect 347016 275110 347044 276934
rect 347004 275104 347056 275110
rect 347004 275046 347056 275052
rect 346176 274832 346228 274838
rect 346176 274774 346228 274780
rect 345900 274696 345952 274702
rect 345900 274638 345952 274644
rect 345348 274424 345400 274430
rect 345348 274366 345400 274372
rect 342588 274084 342640 274090
rect 342588 274026 342640 274032
rect 341944 274016 341996 274022
rect 341944 273958 341996 273964
rect 341116 273948 341168 273954
rect 341116 273890 341168 273896
rect 341128 263906 341156 273890
rect 341852 273880 341904 273886
rect 341852 273822 341904 273828
rect 341760 273812 341812 273818
rect 341760 273754 341812 273760
rect 341772 266542 341800 273754
rect 341760 266536 341812 266542
rect 341760 266478 341812 266484
rect 341864 265658 341892 273822
rect 341852 265652 341904 265658
rect 341852 265594 341904 265600
rect 341956 265590 341984 273958
rect 341944 265584 341996 265590
rect 341944 265526 341996 265532
rect 341128 263878 341340 263906
rect 340682 263742 341064 263770
rect 341312 263770 341340 263878
rect 342600 263770 342628 274026
rect 345808 266536 345860 266542
rect 345808 266478 345860 266484
rect 344796 265652 344848 265658
rect 344796 265594 344848 265600
rect 343784 265584 343836 265590
rect 343784 265526 343836 265532
rect 341312 263742 341694 263770
rect 342600 263742 342706 263770
rect 343796 263756 343824 265526
rect 344808 263756 344836 265594
rect 345820 263756 345848 266478
rect 345912 265658 345940 274638
rect 345992 274560 346044 274566
rect 345992 274502 346044 274508
rect 345900 265652 345952 265658
rect 345900 265594 345952 265600
rect 346004 265590 346032 274502
rect 348028 274294 348056 276934
rect 348764 275178 348792 276934
rect 348752 275172 348804 275178
rect 348752 275114 348804 275120
rect 349592 275042 349620 276934
rect 349580 275036 349632 275042
rect 349580 274978 349632 274984
rect 348200 274764 348252 274770
rect 348200 274706 348252 274712
rect 348016 274288 348068 274294
rect 348016 274230 348068 274236
rect 347924 265652 347976 265658
rect 347924 265594 347976 265600
rect 345992 265584 346044 265590
rect 345992 265526 346044 265532
rect 346820 265584 346872 265590
rect 346820 265526 346872 265532
rect 346832 263756 346860 265526
rect 347936 263756 347964 265594
rect 348212 263906 348240 274706
rect 349580 274628 349632 274634
rect 349580 274570 349632 274576
rect 349488 271772 349540 271778
rect 349488 271714 349540 271720
rect 349500 266202 349528 271714
rect 349488 266196 349540 266202
rect 349488 266138 349540 266144
rect 348212 263878 348424 263906
rect 348396 263770 348424 263878
rect 349592 263770 349620 274570
rect 350420 271778 350448 276934
rect 351248 274974 351276 276934
rect 351236 274968 351288 274974
rect 351236 274910 351288 274916
rect 352168 274906 352196 276934
rect 352156 274900 352208 274906
rect 352156 274842 352208 274848
rect 352996 272458 353024 279330
rect 352800 272452 352852 272458
rect 352800 272394 352852 272400
rect 352984 272452 353036 272458
rect 352984 272394 353036 272400
rect 350408 271772 350460 271778
rect 350408 271714 350460 271720
rect 352062 266776 352118 266785
rect 352062 266711 352118 266720
rect 350958 266640 351014 266649
rect 350958 266575 351014 266584
rect 348396 263742 348962 263770
rect 349592 263742 349974 263770
rect 350972 263756 351000 266575
rect 352076 263756 352104 266711
rect 352812 263770 352840 272394
rect 353548 263906 353576 295106
rect 354008 291022 354036 297175
rect 354192 295850 354220 326590
rect 354916 306248 354968 306254
rect 354916 306190 354968 306196
rect 354180 295844 354232 295850
rect 354180 295786 354232 295792
rect 353996 291016 354048 291022
rect 353996 290958 354048 290964
rect 354272 285508 354324 285514
rect 354272 285450 354324 285456
rect 354284 285281 354312 285450
rect 354270 285272 354326 285281
rect 354270 285207 354326 285216
rect 354928 267902 354956 306190
rect 355572 300678 355600 327270
rect 356768 327062 356796 329852
rect 357596 327538 357624 329852
rect 357584 327532 357636 327538
rect 357584 327474 357636 327480
rect 358320 327192 358372 327198
rect 358320 327134 358372 327140
rect 356756 327056 356808 327062
rect 356756 326998 356808 327004
rect 355652 326784 355704 326790
rect 355652 326726 355704 326732
rect 355664 306254 355692 326726
rect 356940 326580 356992 326586
rect 356940 326522 356992 326528
rect 356202 314104 356258 314113
rect 356202 314039 356258 314048
rect 356216 313802 356244 314039
rect 356204 313796 356256 313802
rect 356204 313738 356256 313744
rect 356952 310334 356980 326522
rect 358332 315910 358360 327134
rect 358424 327130 358452 329852
rect 358412 327124 358464 327130
rect 358412 327066 358464 327072
rect 357676 315904 357728 315910
rect 357676 315846 357728 315852
rect 358320 315904 358372 315910
rect 358320 315846 358372 315852
rect 356940 310328 356992 310334
rect 356940 310270 356992 310276
rect 356952 309722 356980 310270
rect 356296 309716 356348 309722
rect 356296 309658 356348 309664
rect 356940 309716 356992 309722
rect 356940 309658 356992 309664
rect 356202 308664 356258 308673
rect 356202 308599 356258 308608
rect 356216 308294 356244 308599
rect 356204 308288 356256 308294
rect 356204 308230 356256 308236
rect 355652 306248 355704 306254
rect 355652 306190 355704 306196
rect 356202 304176 356258 304185
rect 356202 304111 356204 304120
rect 356256 304111 356258 304120
rect 356204 304082 356256 304088
rect 355560 300672 355612 300678
rect 355560 300614 355612 300620
rect 355572 300066 355600 300614
rect 355008 300060 355060 300066
rect 355008 300002 355060 300008
rect 355560 300060 355612 300066
rect 355560 300002 355612 300008
rect 354916 267896 354968 267902
rect 354916 267838 354968 267844
rect 353548 263878 353852 263906
rect 353824 263770 353852 263878
rect 355020 263770 355048 300002
rect 356202 298872 356258 298881
rect 356202 298807 356258 298816
rect 356216 298638 356244 298807
rect 356204 298632 356256 298638
rect 356204 298574 356256 298580
rect 356202 293840 356258 293849
rect 356202 293775 356204 293784
rect 356256 293775 356258 293784
rect 356204 293746 356256 293752
rect 356202 289080 356258 289089
rect 356202 289015 356258 289024
rect 356216 288982 356244 289015
rect 356204 288976 356256 288982
rect 356204 288918 356256 288924
rect 356202 283776 356258 283785
rect 356202 283711 356258 283720
rect 356216 283474 356244 283711
rect 356204 283468 356256 283474
rect 356204 283410 356256 283416
rect 356202 279424 356258 279433
rect 356202 279359 356258 279368
rect 356216 279326 356244 279359
rect 356204 279320 356256 279326
rect 356204 279262 356256 279268
rect 355836 267896 355888 267902
rect 355836 267838 355888 267844
rect 356308 267850 356336 309658
rect 355848 263770 355876 267838
rect 356308 267822 356980 267850
rect 356952 263770 356980 267822
rect 357688 263906 357716 315846
rect 357688 263878 357900 263906
rect 357872 263770 357900 263878
rect 352812 263742 353102 263770
rect 353824 263742 354114 263770
rect 355020 263742 355126 263770
rect 355848 263742 356230 263770
rect 356952 263742 357242 263770
rect 357872 263742 358254 263770
rect 330824 263606 331390 263634
rect 328418 263512 328474 263521
rect 328418 263447 328474 263456
rect 358412 263476 358464 263482
rect 358412 263418 358464 263424
rect 327682 261744 327738 261753
rect 327682 261679 327738 261688
rect 327696 261442 327724 261679
rect 327684 261436 327736 261442
rect 327684 261378 327736 261384
rect 327958 260384 328014 260393
rect 327958 260319 328014 260328
rect 327222 258888 327278 258897
rect 327222 258823 327278 258832
rect 327130 257528 327186 257537
rect 327130 257463 327186 257472
rect 327144 255866 327172 257463
rect 327132 255860 327184 255866
rect 327132 255802 327184 255808
rect 327236 255798 327264 258823
rect 327972 257226 328000 260319
rect 327960 257220 328012 257226
rect 327960 257162 328012 257168
rect 328510 256168 328566 256177
rect 328510 256103 328566 256112
rect 327224 255792 327276 255798
rect 327224 255734 327276 255740
rect 328418 254672 328474 254681
rect 328418 254607 328474 254616
rect 328432 254506 328460 254607
rect 328420 254500 328472 254506
rect 328420 254442 328472 254448
rect 328524 253962 328552 256103
rect 328512 253956 328564 253962
rect 328512 253898 328564 253904
rect 327130 253312 327186 253321
rect 327130 253247 327186 253256
rect 327144 251922 327172 253247
rect 327222 251952 327278 251961
rect 327132 251916 327184 251922
rect 327222 251887 327278 251896
rect 327132 251858 327184 251864
rect 327236 251038 327264 251887
rect 327224 251032 327276 251038
rect 327224 250974 327276 250980
rect 327222 250592 327278 250601
rect 327222 250527 327278 250536
rect 327236 249542 327264 250527
rect 327224 249536 327276 249542
rect 327224 249478 327276 249484
rect 328420 249128 328472 249134
rect 328418 249096 328420 249105
rect 328472 249096 328474 249105
rect 328418 249031 328474 249040
rect 328418 247736 328474 247745
rect 328418 247671 328420 247680
rect 328472 247671 328474 247680
rect 328420 247642 328472 247648
rect 328420 247564 328472 247570
rect 328420 247506 328472 247512
rect 328432 246929 328460 247506
rect 328418 246920 328474 246929
rect 328418 246855 328474 246864
rect 327868 246204 327920 246210
rect 327868 246146 327920 246152
rect 327880 245569 327908 246146
rect 327866 245560 327922 245569
rect 327866 245495 327922 245504
rect 327868 244776 327920 244782
rect 327868 244718 327920 244724
rect 327880 244073 327908 244718
rect 327866 244064 327922 244073
rect 327866 243999 327922 244008
rect 327224 243484 327276 243490
rect 327224 243426 327276 243432
rect 327236 240673 327264 243426
rect 327868 243416 327920 243422
rect 327868 243358 327920 243364
rect 327880 242713 327908 243358
rect 327866 242704 327922 242713
rect 327866 242639 327922 242648
rect 328052 242260 328104 242266
rect 328052 242202 328104 242208
rect 327868 242124 327920 242130
rect 327868 242066 327920 242072
rect 327222 240664 327278 240673
rect 327222 240599 327278 240608
rect 327880 238633 327908 242066
rect 328064 239313 328092 242202
rect 328050 239304 328106 239313
rect 328050 239239 328106 239248
rect 327866 238624 327922 238633
rect 327866 238559 327922 238568
rect 328420 236616 328472 236622
rect 328418 236584 328420 236593
rect 328472 236584 328474 236593
rect 328418 236519 328474 236528
rect 330088 235862 331390 235890
rect 332402 235862 332784 235890
rect 326580 232264 326632 232270
rect 326580 232206 326632 232212
rect 325844 224308 325896 224314
rect 325844 224250 325896 224256
rect 325750 220128 325806 220137
rect 325750 220063 325806 220072
rect 325856 217009 325884 224250
rect 325842 217000 325898 217009
rect 325842 216935 325898 216944
rect 325658 210744 325714 210753
rect 325658 210679 325714 210688
rect 325566 204488 325622 204497
rect 325566 204423 325622 204432
rect 325476 202072 325528 202078
rect 325476 202014 325528 202020
rect 325382 191976 325438 191985
rect 325382 191911 325438 191920
rect 325290 185720 325346 185729
rect 325290 185655 325346 185664
rect 325488 182601 325516 202014
rect 330088 188954 330116 235862
rect 332756 224994 332784 235862
rect 333400 232474 333428 235876
rect 334412 232474 334440 235876
rect 333388 232468 333440 232474
rect 333388 232410 333440 232416
rect 334124 232468 334176 232474
rect 334124 232410 334176 232416
rect 334400 232468 334452 232474
rect 334400 232410 334452 232416
rect 335412 232468 335464 232474
rect 335412 232410 335464 232416
rect 332744 224988 332796 224994
rect 332744 224930 332796 224936
rect 334136 224926 334164 232410
rect 335424 225062 335452 232410
rect 335412 225056 335464 225062
rect 335412 224998 335464 225004
rect 334124 224920 334176 224926
rect 334124 224862 334176 224868
rect 335516 224858 335544 235876
rect 336542 235862 336924 235890
rect 337554 235862 338304 235890
rect 335504 224852 335556 224858
rect 335504 224794 335556 224800
rect 336896 224586 336924 235862
rect 337160 225260 337212 225266
rect 337160 225202 337212 225208
rect 336884 224580 336936 224586
rect 336884 224522 336936 224528
rect 337172 222834 337200 225202
rect 337712 225124 337764 225130
rect 337712 225066 337764 225072
rect 337724 222834 337752 225066
rect 338276 224450 338304 235862
rect 338552 232474 338580 235876
rect 339564 235862 339670 235890
rect 340682 235862 341064 235890
rect 338540 232468 338592 232474
rect 338540 232410 338592 232416
rect 339564 226642 339592 235862
rect 340932 233556 340984 233562
rect 340932 233498 340984 233504
rect 340840 233420 340892 233426
rect 340840 233362 340892 233368
rect 339644 232468 339696 232474
rect 339644 232410 339696 232416
rect 339472 226614 339592 226642
rect 338356 225464 338408 225470
rect 338356 225406 338408 225412
rect 338264 224444 338316 224450
rect 338264 224386 338316 224392
rect 338368 222834 338396 225406
rect 339000 225192 339052 225198
rect 339000 225134 339052 225140
rect 339012 222834 339040 225134
rect 339472 224382 339500 226614
rect 339656 224790 339684 232410
rect 339644 224784 339696 224790
rect 339644 224726 339696 224732
rect 339552 224716 339604 224722
rect 339552 224658 339604 224664
rect 339460 224376 339512 224382
rect 339460 224318 339512 224324
rect 339564 222834 339592 224658
rect 340852 223242 340880 233362
rect 340760 223214 340880 223242
rect 337172 222806 337232 222834
rect 337724 222806 337784 222834
rect 338368 222806 338428 222834
rect 339012 222806 339072 222834
rect 339564 222806 339624 222834
rect 340760 222562 340788 223214
rect 340944 223106 340972 233498
rect 341036 225146 341064 235862
rect 341128 235862 341694 235890
rect 342508 235862 342706 235890
rect 343520 235862 343810 235890
rect 341128 225266 341156 235862
rect 341116 225260 341168 225266
rect 341116 225202 341168 225208
rect 341208 225260 341260 225266
rect 341208 225202 341260 225208
rect 341220 225146 341248 225202
rect 341036 225118 341248 225146
rect 342036 225192 342088 225198
rect 342036 225134 342088 225140
rect 341392 224512 341444 224518
rect 341392 224454 341444 224460
rect 340898 223078 340972 223106
rect 340898 222820 340926 223078
rect 341404 222834 341432 224454
rect 342048 222834 342076 225134
rect 342508 225130 342536 235862
rect 342680 232468 342732 232474
rect 342680 232410 342732 232416
rect 342496 225124 342548 225130
rect 342496 225066 342548 225072
rect 342692 224722 342720 232410
rect 343232 229680 343284 229686
rect 343232 229622 343284 229628
rect 342680 224716 342732 224722
rect 342680 224658 342732 224664
rect 342726 223084 342778 223090
rect 342726 223026 342778 223032
rect 342738 222954 342766 223026
rect 342726 222948 342778 222954
rect 342726 222890 342778 222896
rect 341404 222806 341464 222834
rect 342048 222806 342108 222834
rect 342738 222820 342766 222890
rect 343244 222834 343272 229622
rect 343520 225470 343548 235862
rect 344808 232474 344836 235876
rect 345360 235862 345834 235890
rect 345256 233828 345308 233834
rect 345256 233770 345308 233776
rect 344796 232468 344848 232474
rect 344796 232410 344848 232416
rect 343784 230292 343836 230298
rect 343784 230234 343836 230240
rect 343796 229686 343824 230234
rect 343784 229680 343836 229686
rect 343784 229622 343836 229628
rect 345268 228938 345296 233770
rect 345256 228932 345308 228938
rect 345256 228874 345308 228880
rect 345164 227708 345216 227714
rect 345164 227650 345216 227656
rect 345176 227034 345204 227650
rect 343876 227028 343928 227034
rect 343876 226970 343928 226976
rect 345164 227028 345216 227034
rect 345164 226970 345216 226976
rect 343508 225464 343560 225470
rect 343508 225406 343560 225412
rect 343888 222834 343916 226970
rect 345360 224654 345388 235862
rect 346544 234440 346596 234446
rect 346544 234382 346596 234388
rect 346556 233834 346584 234382
rect 346544 233828 346596 233834
rect 346544 233770 346596 233776
rect 346832 233426 346860 235876
rect 347936 233562 347964 235876
rect 348028 235862 348962 235890
rect 347924 233556 347976 233562
rect 347924 233498 347976 233504
rect 346820 233420 346872 233426
rect 346820 233362 346872 233368
rect 345716 231720 345768 231726
rect 345716 231662 345768 231668
rect 345728 231046 345756 231662
rect 345440 231040 345492 231046
rect 345440 230982 345492 230988
rect 345716 231040 345768 231046
rect 345716 230982 345768 230988
rect 345348 224648 345400 224654
rect 345348 224590 345400 224596
rect 345164 224308 345216 224314
rect 345164 224250 345216 224256
rect 344520 224240 344572 224246
rect 344520 224182 344572 224188
rect 344532 222834 344560 224182
rect 345176 222834 345204 224250
rect 345452 222834 345480 230982
rect 346084 228932 346136 228938
rect 346084 228874 346136 228880
rect 346096 222834 346124 228874
rect 347188 226348 347240 226354
rect 347188 226290 347240 226296
rect 347200 225742 347228 226290
rect 347188 225736 347240 225742
rect 347188 225678 347240 225684
rect 343244 222806 343304 222834
rect 343888 222806 343948 222834
rect 344532 222806 344592 222834
rect 345176 222806 345236 222834
rect 345452 222806 345788 222834
rect 346096 222806 346432 222834
rect 347200 222698 347228 225678
rect 347280 224988 347332 224994
rect 347280 224930 347332 224936
rect 347292 222834 347320 224930
rect 347924 224920 347976 224926
rect 347924 224862 347976 224868
rect 347936 224330 347964 224862
rect 348028 224518 348056 235862
rect 349960 232474 349988 235876
rect 350972 232513 351000 235876
rect 352076 232513 352104 235876
rect 352720 235862 353102 235890
rect 353548 235862 354114 235890
rect 355020 235862 355126 235890
rect 355848 235862 356230 235890
rect 356308 235862 357242 235890
rect 357688 235862 358254 235890
rect 350958 232504 351014 232513
rect 348108 232468 348160 232474
rect 348108 232410 348160 232416
rect 349948 232468 350000 232474
rect 350958 232439 351014 232448
rect 352062 232504 352118 232513
rect 352062 232439 352118 232448
rect 349948 232410 350000 232416
rect 348120 225198 348148 232410
rect 350960 225464 351012 225470
rect 350960 225406 351012 225412
rect 348108 225192 348160 225198
rect 348108 225134 348160 225140
rect 348568 225056 348620 225062
rect 348568 224998 348620 225004
rect 348016 224512 348068 224518
rect 348016 224454 348068 224460
rect 347936 224302 348056 224330
rect 348028 222834 348056 224302
rect 348580 222834 348608 224998
rect 349396 224852 349448 224858
rect 349396 224794 349448 224800
rect 349408 222834 349436 224794
rect 349764 224580 349816 224586
rect 349764 224522 349816 224528
rect 349776 222834 349804 224522
rect 350684 224444 350736 224450
rect 350684 224386 350736 224392
rect 350696 223106 350724 224386
rect 350696 223078 350770 223106
rect 347292 222806 347628 222834
rect 348028 222806 348272 222834
rect 348580 222806 348916 222834
rect 349408 222806 349468 222834
rect 349776 222806 350112 222834
rect 350742 222820 350770 223078
rect 350972 222834 351000 225406
rect 352248 225260 352300 225266
rect 352248 225202 352300 225208
rect 351604 224376 351656 224382
rect 351604 224318 351656 224324
rect 351616 222834 351644 224318
rect 352260 222834 352288 225202
rect 350972 222806 351308 222834
rect 351616 222806 351952 222834
rect 352260 222806 352596 222834
rect 347076 222670 347228 222698
rect 340268 222534 340788 222562
rect 334214 216184 334270 216193
rect 334214 216119 334270 216128
rect 334228 215882 334256 216119
rect 334216 215876 334268 215882
rect 334216 215818 334268 215824
rect 334214 202856 334270 202865
rect 334214 202791 334270 202800
rect 334228 202078 334256 202791
rect 334216 202072 334268 202078
rect 334216 202014 334268 202020
rect 352720 195822 352748 235862
rect 352892 233080 352944 233086
rect 352892 233022 352944 233028
rect 352800 218664 352852 218670
rect 352800 218606 352852 218612
rect 352708 195816 352760 195822
rect 352708 195758 352760 195764
rect 334214 189528 334270 189537
rect 334214 189463 334270 189472
rect 330076 188948 330128 188954
rect 330076 188890 330128 188896
rect 326580 188268 326632 188274
rect 326580 188210 326632 188216
rect 325474 182592 325530 182601
rect 325474 182527 325530 182536
rect 326592 179910 326620 188210
rect 326580 179904 326632 179910
rect 326580 179846 326632 179852
rect 328420 170248 328472 170254
rect 328420 170190 328472 170196
rect 328432 169137 328460 170190
rect 330088 169930 330116 188890
rect 334228 188274 334256 189463
rect 334216 188268 334268 188274
rect 334216 188210 334268 188216
rect 337324 182822 337660 182850
rect 338152 182822 338304 182850
rect 338980 182822 339316 182850
rect 339808 182822 340144 182850
rect 340636 182822 340972 182850
rect 341464 182822 341708 182850
rect 342292 182822 342444 182850
rect 343212 182822 343548 182850
rect 344040 182822 344376 182850
rect 344868 182822 345204 182850
rect 337632 181338 337660 182822
rect 337620 181332 337672 181338
rect 337620 181274 337672 181280
rect 338276 181202 338304 182822
rect 338264 181196 338316 181202
rect 338264 181138 338316 181144
rect 336884 181060 336936 181066
rect 336884 181002 336936 181008
rect 334124 180992 334176 180998
rect 334124 180934 334176 180940
rect 332744 180720 332796 180726
rect 332744 180662 332796 180668
rect 330088 169902 330852 169930
rect 330824 169658 330852 169902
rect 332756 169794 332784 180662
rect 334136 173042 334164 180934
rect 335412 180788 335464 180794
rect 335412 180730 335464 180736
rect 333388 173036 333440 173042
rect 333388 172978 333440 172984
rect 334124 173036 334176 173042
rect 334124 172978 334176 172984
rect 332402 169766 332784 169794
rect 333400 169780 333428 172978
rect 335424 172090 335452 180730
rect 335504 180652 335556 180658
rect 335504 180594 335556 180600
rect 334400 172084 334452 172090
rect 334400 172026 334452 172032
rect 335412 172084 335464 172090
rect 335412 172026 335464 172032
rect 334412 169780 334440 172026
rect 335516 169780 335544 180594
rect 336896 169794 336924 181002
rect 338264 180584 338316 180590
rect 338264 180526 338316 180532
rect 336542 169766 336924 169794
rect 338276 169658 338304 180526
rect 339288 180522 339316 182822
rect 340116 181134 340144 182822
rect 340104 181128 340156 181134
rect 340104 181070 340156 181076
rect 339644 180992 339696 180998
rect 339644 180934 339696 180940
rect 339276 180516 339328 180522
rect 339276 180458 339328 180464
rect 338540 172356 338592 172362
rect 338540 172298 338592 172304
rect 338552 169780 338580 172298
rect 339656 169780 339684 180934
rect 340944 180454 340972 182822
rect 341116 181332 341168 181338
rect 341116 181274 341168 181280
rect 341024 180856 341076 180862
rect 341024 180798 341076 180804
rect 340932 180448 340984 180454
rect 340932 180390 340984 180396
rect 341036 169794 341064 180798
rect 340682 169766 341064 169794
rect 330824 169630 331390 169658
rect 337554 169630 338304 169658
rect 341128 169658 341156 181274
rect 341680 180114 341708 182822
rect 341852 181196 341904 181202
rect 341852 181138 341904 181144
rect 341760 180516 341812 180522
rect 341760 180458 341812 180464
rect 341668 180108 341720 180114
rect 341668 180050 341720 180056
rect 341772 172974 341800 180458
rect 341864 173042 341892 181138
rect 342416 179978 342444 182822
rect 343520 180182 343548 182822
rect 343876 181128 343928 181134
rect 343876 181070 343928 181076
rect 343508 180176 343560 180182
rect 343508 180118 343560 180124
rect 342404 179972 342456 179978
rect 342404 179914 342456 179920
rect 341852 173036 341904 173042
rect 341852 172978 341904 172984
rect 342680 173036 342732 173042
rect 342680 172978 342732 172984
rect 341760 172968 341812 172974
rect 341760 172910 341812 172916
rect 342692 169780 342720 172978
rect 343784 172968 343836 172974
rect 343784 172910 343836 172916
rect 343796 169780 343824 172910
rect 343888 169658 343916 181070
rect 344348 180046 344376 182822
rect 345176 181338 345204 182822
rect 345360 182822 345696 182850
rect 346188 182822 346524 182850
rect 347016 182822 347352 182850
rect 348028 182822 348272 182850
rect 348764 182822 349100 182850
rect 349592 182822 349928 182850
rect 350756 182822 350816 182850
rect 345164 181332 345216 181338
rect 345164 181274 345216 181280
rect 345360 180726 345388 182822
rect 346188 181270 346216 182822
rect 346176 181264 346228 181270
rect 346176 181206 346228 181212
rect 347016 180794 347044 182822
rect 347004 180788 347056 180794
rect 347004 180730 347056 180736
rect 345348 180720 345400 180726
rect 345348 180662 345400 180668
rect 348028 180658 348056 182822
rect 348764 181066 348792 182822
rect 348752 181060 348804 181066
rect 348752 181002 348804 181008
rect 348016 180652 348068 180658
rect 348016 180594 348068 180600
rect 349592 180590 349620 182822
rect 349580 180584 349632 180590
rect 349580 180526 349632 180532
rect 344612 180448 344664 180454
rect 344612 180390 344664 180396
rect 344336 180040 344388 180046
rect 344336 179982 344388 179988
rect 344520 179972 344572 179978
rect 344520 179914 344572 179920
rect 344532 171886 344560 179914
rect 344520 171880 344572 171886
rect 344520 171822 344572 171828
rect 344624 171750 344652 180390
rect 348016 180176 348068 180182
rect 348016 180118 348068 180124
rect 344704 180108 344756 180114
rect 344704 180050 344756 180056
rect 344716 171818 344744 180050
rect 347280 180040 347332 180046
rect 347280 179982 347332 179988
rect 347292 173042 347320 179982
rect 347280 173036 347332 173042
rect 347280 172978 347332 172984
rect 347924 171880 347976 171886
rect 347924 171822 347976 171828
rect 344704 171812 344756 171818
rect 344704 171754 344756 171760
rect 346820 171812 346872 171818
rect 346820 171754 346872 171760
rect 344612 171744 344664 171750
rect 344612 171686 344664 171692
rect 345808 171744 345860 171750
rect 345808 171686 345860 171692
rect 345820 169780 345848 171686
rect 346832 169780 346860 171754
rect 347936 169780 347964 171822
rect 348028 169658 348056 180118
rect 350788 177682 350816 182822
rect 351248 182822 351584 182850
rect 352168 182822 352412 182850
rect 351248 180998 351276 182822
rect 352168 181746 352196 182822
rect 352156 181740 352208 181746
rect 352156 181682 352208 181688
rect 351236 180992 351288 180998
rect 351236 180934 351288 180940
rect 350696 177654 350816 177682
rect 349948 173036 350000 173042
rect 349948 172978 350000 172984
rect 349960 169780 349988 172978
rect 350696 172362 350724 177654
rect 350958 172664 351014 172673
rect 350958 172599 351014 172608
rect 352062 172664 352118 172673
rect 352062 172599 352118 172608
rect 350684 172356 350736 172362
rect 350684 172298 350736 172304
rect 350972 169780 351000 172599
rect 352076 169780 352104 172599
rect 352720 169794 352748 195758
rect 352812 191826 352840 218606
rect 352904 218602 352932 233022
rect 353076 227640 353128 227646
rect 353076 227582 353128 227588
rect 352892 218596 352944 218602
rect 352892 218538 352944 218544
rect 352984 217236 353036 217242
rect 352984 217178 353036 217184
rect 352812 191798 352932 191826
rect 352800 191668 352852 191674
rect 352800 191610 352852 191616
rect 352812 191441 352840 191610
rect 352798 191432 352854 191441
rect 352798 191367 352854 191376
rect 352800 186160 352852 186166
rect 352800 186102 352852 186108
rect 352812 184097 352840 186102
rect 352798 184088 352854 184097
rect 352798 184023 352854 184032
rect 352904 182193 352932 191798
rect 352890 182184 352946 182193
rect 352890 182119 352946 182128
rect 352996 182057 353024 217178
rect 353088 214318 353116 227582
rect 353168 226280 353220 226286
rect 353168 226222 353220 226228
rect 353180 215814 353208 226222
rect 353260 226212 353312 226218
rect 353260 226154 353312 226160
rect 353168 215808 353220 215814
rect 353168 215750 353220 215756
rect 353272 215746 353300 226154
rect 353352 226144 353404 226150
rect 353352 226086 353404 226092
rect 353364 217106 353392 226086
rect 353444 220636 353496 220642
rect 353444 220578 353496 220584
rect 353352 217100 353404 217106
rect 353352 217042 353404 217048
rect 353260 215740 353312 215746
rect 353260 215682 353312 215688
rect 353076 214312 353128 214318
rect 353076 214254 353128 214260
rect 353456 213094 353484 220578
rect 353444 213088 353496 213094
rect 353444 213030 353496 213036
rect 353548 201330 353576 235862
rect 354916 228932 354968 228938
rect 354916 228874 354968 228880
rect 354928 210986 354956 228874
rect 354916 210980 354968 210986
rect 354916 210922 354968 210928
rect 353536 201324 353588 201330
rect 353536 201266 353588 201272
rect 352982 182048 353038 182057
rect 352982 181983 353038 181992
rect 353548 169930 353576 201266
rect 354928 172634 354956 210922
rect 355020 206838 355048 235862
rect 355848 228938 355876 235862
rect 355836 228932 355888 228938
rect 355836 228874 355888 228880
rect 355098 220264 355154 220273
rect 355098 220199 355154 220208
rect 355112 213978 355140 220199
rect 356308 215921 356336 235862
rect 356294 215912 356350 215921
rect 356294 215847 356350 215856
rect 356202 215232 356258 215241
rect 356202 215167 356258 215176
rect 356216 214114 356244 215167
rect 356204 214108 356256 214114
rect 356204 214050 356256 214056
rect 355100 213972 355152 213978
rect 355100 213914 355152 213920
rect 356202 210200 356258 210209
rect 356202 210135 356258 210144
rect 356216 209626 356244 210135
rect 356204 209620 356256 209626
rect 356204 209562 356256 209568
rect 355008 206832 355060 206838
rect 355008 206774 355060 206780
rect 354916 172628 354968 172634
rect 354916 172570 354968 172576
rect 353548 169902 353852 169930
rect 353824 169794 353852 169902
rect 355020 169794 355048 206774
rect 356202 205304 356258 205313
rect 356202 205239 356258 205248
rect 356216 204798 356244 205239
rect 356204 204792 356256 204798
rect 356204 204734 356256 204740
rect 356202 200272 356258 200281
rect 356202 200207 356258 200216
rect 356216 199290 356244 200207
rect 356204 199284 356256 199290
rect 356204 199226 356256 199232
rect 356202 195240 356258 195249
rect 356202 195175 356258 195184
rect 356216 195142 356244 195175
rect 356204 195136 356256 195142
rect 356204 195078 356256 195084
rect 356202 190208 356258 190217
rect 356202 190143 356258 190152
rect 356216 189634 356244 190143
rect 356204 189628 356256 189634
rect 356204 189570 356256 189576
rect 356202 185312 356258 185321
rect 356202 185247 356258 185256
rect 356216 184058 356244 185247
rect 356204 184052 356256 184058
rect 356204 183994 356256 184000
rect 355836 172628 355888 172634
rect 355836 172570 355888 172576
rect 355848 169794 355876 172570
rect 356308 169930 356336 215847
rect 357688 214046 357716 235862
rect 358320 231040 358372 231046
rect 358320 230982 358372 230988
rect 358332 229634 358360 230982
rect 358240 229606 358360 229634
rect 358240 224858 358268 229606
rect 358044 224852 358096 224858
rect 358044 224794 358096 224800
rect 358228 224852 358280 224858
rect 358228 224794 358280 224800
rect 358056 220001 358084 224794
rect 358042 219992 358098 220001
rect 358042 219927 358098 219936
rect 358226 219992 358282 220001
rect 358226 219927 358282 219936
rect 358240 215542 358268 219927
rect 358424 215678 358452 263418
rect 358516 239954 358544 393366
rect 358608 240022 358636 393774
rect 372960 393226 372988 396344
rect 372948 393220 373000 393226
rect 372948 393162 373000 393168
rect 390624 393158 390652 396344
rect 408380 393362 408408 396344
rect 408368 393356 408420 393362
rect 408368 393298 408420 393304
rect 426044 393294 426072 396344
rect 426032 393288 426084 393294
rect 426032 393230 426084 393236
rect 390612 393152 390664 393158
rect 390612 393094 390664 393100
rect 429434 390536 429490 390545
rect 429434 390471 429490 390480
rect 429448 389758 429476 390471
rect 429436 389752 429488 389758
rect 429436 389694 429488 389700
rect 429436 378668 429488 378674
rect 429436 378610 429488 378616
rect 429448 378033 429476 378610
rect 429434 378024 429490 378033
rect 429434 377959 429490 377968
rect 362460 371800 362512 371806
rect 362460 371742 362512 371748
rect 359700 327260 359752 327266
rect 359700 327202 359752 327208
rect 358596 240016 358648 240022
rect 358596 239958 358648 239964
rect 358504 239948 358556 239954
rect 358504 239890 358556 239896
rect 359712 235126 359740 327202
rect 360712 262796 360764 262802
rect 360712 262738 360764 262744
rect 360436 262048 360488 262054
rect 360436 261990 360488 261996
rect 359700 235120 359752 235126
rect 359700 235062 359752 235068
rect 360448 226014 360476 261990
rect 360620 259328 360672 259334
rect 360620 259270 360672 259276
rect 360632 259169 360660 259270
rect 360618 259160 360674 259169
rect 360618 259095 360674 259104
rect 360526 256032 360582 256041
rect 360526 255967 360582 255976
rect 360540 231726 360568 255967
rect 360632 234446 360660 259095
rect 360724 252913 360752 262738
rect 360802 262288 360858 262297
rect 360802 262223 360858 262232
rect 360816 262054 360844 262223
rect 360804 262048 360856 262054
rect 360804 261990 360856 261996
rect 361172 256540 361224 256546
rect 361172 256482 361224 256488
rect 361184 256041 361212 256482
rect 361170 256032 361226 256041
rect 361170 255967 361226 255976
rect 361172 253072 361224 253078
rect 361172 253014 361224 253020
rect 361184 252913 361212 253014
rect 360710 252904 360766 252913
rect 360710 252839 360766 252848
rect 361170 252904 361226 252913
rect 361170 252839 361226 252848
rect 360710 249776 360766 249785
rect 360710 249711 360766 249720
rect 360724 249610 360752 249711
rect 360712 249604 360764 249610
rect 360712 249546 360764 249552
rect 360620 234440 360672 234446
rect 360620 234382 360672 234388
rect 360528 231720 360580 231726
rect 360528 231662 360580 231668
rect 360436 226008 360488 226014
rect 360436 225950 360488 225956
rect 359700 225872 359752 225878
rect 359700 225814 359752 225820
rect 358412 215672 358464 215678
rect 358412 215614 358464 215620
rect 358228 215536 358280 215542
rect 358228 215478 358280 215484
rect 358412 215536 358464 215542
rect 358412 215478 358464 215484
rect 357676 214040 357728 214046
rect 357676 213982 357728 213988
rect 357688 169930 357716 213982
rect 358424 211705 358452 215478
rect 358410 211696 358466 211705
rect 358410 211631 358466 211640
rect 358594 211696 358650 211705
rect 358594 211631 358650 211640
rect 358608 202078 358636 211631
rect 358412 202072 358464 202078
rect 358412 202014 358464 202020
rect 358596 202072 358648 202078
rect 358596 202014 358648 202020
rect 358424 185570 358452 202014
rect 358240 185542 358452 185570
rect 358240 185434 358268 185542
rect 358240 185406 358360 185434
rect 358332 175966 358360 185406
rect 358320 175960 358372 175966
rect 358320 175902 358372 175908
rect 358320 175824 358372 175830
rect 358320 175766 358372 175772
rect 358332 173058 358360 175766
rect 358332 173030 358452 173058
rect 358424 171614 358452 173030
rect 358412 171608 358464 171614
rect 358412 171550 358464 171556
rect 358596 171608 358648 171614
rect 358596 171550 358648 171556
rect 356308 169902 356796 169930
rect 357688 169902 357900 169930
rect 352720 169766 353102 169794
rect 353824 169766 354114 169794
rect 355020 169766 355126 169794
rect 355848 169766 356230 169794
rect 356768 169658 356796 169902
rect 357872 169794 357900 169902
rect 357872 169766 358254 169794
rect 341128 169630 341694 169658
rect 343888 169630 344822 169658
rect 348028 169630 348962 169658
rect 356768 169630 357242 169658
rect 328418 169128 328474 169137
rect 328418 169063 328474 169072
rect 327222 167768 327278 167777
rect 327222 167703 327278 167712
rect 327236 163522 327264 167703
rect 328418 166408 328474 166417
rect 328418 166343 328474 166352
rect 328432 166242 328460 166343
rect 328420 166236 328472 166242
rect 328420 166178 328472 166184
rect 328510 164912 328566 164921
rect 328510 164847 328566 164856
rect 328524 164814 328552 164847
rect 328512 164808 328564 164814
rect 328512 164750 328564 164756
rect 327224 163516 327276 163522
rect 327224 163458 327276 163464
rect 327222 163416 327278 163425
rect 358608 163386 358636 171550
rect 359712 168894 359740 225814
rect 360724 224994 360752 249546
rect 360802 246648 360858 246657
rect 360802 246583 360858 246592
rect 360816 227714 360844 246583
rect 360894 243520 360950 243529
rect 360894 243455 360950 243464
rect 360908 230298 360936 243455
rect 360986 240392 361042 240401
rect 360986 240327 361042 240336
rect 360896 230292 360948 230298
rect 360896 230234 360948 230240
rect 360804 227708 360856 227714
rect 360804 227650 360856 227656
rect 360712 224988 360764 224994
rect 360712 224930 360764 224936
rect 361000 224790 361028 240327
rect 361262 237400 361318 237409
rect 361262 237335 361318 237344
rect 361172 224988 361224 224994
rect 361172 224930 361224 224936
rect 360988 224784 361040 224790
rect 360988 224726 361040 224732
rect 361184 224246 361212 224930
rect 361172 224240 361224 224246
rect 361172 224182 361224 224188
rect 361080 221520 361132 221526
rect 361080 221462 361132 221468
rect 359792 220092 359844 220098
rect 359792 220034 359844 220040
rect 359804 181338 359832 220034
rect 359792 181332 359844 181338
rect 359792 181274 359844 181280
rect 359700 168888 359752 168894
rect 359700 168830 359752 168836
rect 359712 168321 359740 168830
rect 359054 168312 359110 168321
rect 359054 168247 359110 168256
rect 359698 168312 359754 168321
rect 359698 168247 359754 168256
rect 327222 163351 327278 163360
rect 358596 163380 358648 163386
rect 327236 161346 327264 163351
rect 358596 163322 358648 163328
rect 328418 162192 328474 162201
rect 328418 162127 328474 162136
rect 328432 162094 328460 162127
rect 328420 162088 328472 162094
rect 328420 162030 328472 162036
rect 327224 161340 327276 161346
rect 327224 161282 327276 161288
rect 327314 160696 327370 160705
rect 327314 160631 327370 160640
rect 327222 159336 327278 159345
rect 327222 159271 327278 159280
rect 327236 158218 327264 159271
rect 327224 158212 327276 158218
rect 327224 158154 327276 158160
rect 327328 158082 327356 160631
rect 327316 158076 327368 158082
rect 327316 158018 327368 158024
rect 327222 157976 327278 157985
rect 327222 157911 327278 157920
rect 327236 157266 327264 157911
rect 327224 157260 327276 157266
rect 327224 157202 327276 157208
rect 327222 156616 327278 156625
rect 327222 156551 327278 156560
rect 327236 155974 327264 156551
rect 358596 156444 358648 156450
rect 358596 156386 358648 156392
rect 327224 155968 327276 155974
rect 327224 155910 327276 155916
rect 328418 155120 328474 155129
rect 328418 155055 328420 155064
rect 328472 155055 328474 155064
rect 328420 155026 328472 155032
rect 328420 153792 328472 153798
rect 328418 153760 328420 153769
rect 328472 153760 328474 153769
rect 358608 153746 358636 156386
rect 358608 153718 358728 153746
rect 328418 153695 328474 153704
rect 328420 152432 328472 152438
rect 328418 152400 328420 152409
rect 328472 152400 328474 152409
rect 328418 152335 328474 152344
rect 328420 150936 328472 150942
rect 328418 150904 328420 150913
rect 328472 150904 328474 150913
rect 328418 150839 328474 150848
rect 327224 149780 327276 149786
rect 327224 149722 327276 149728
rect 327236 146697 327264 149722
rect 328420 149576 328472 149582
rect 328418 149544 328420 149553
rect 328472 149544 328474 149553
rect 328418 149479 328474 149488
rect 327868 148420 327920 148426
rect 327868 148362 327920 148368
rect 327222 146688 327278 146697
rect 327222 146623 327278 146632
rect 327880 145337 327908 148362
rect 328420 148216 328472 148222
rect 328418 148184 328420 148193
rect 328472 148184 328474 148193
rect 328418 148119 328474 148128
rect 327866 145328 327922 145337
rect 327866 145263 327922 145272
rect 326580 144748 326632 144754
rect 326580 144690 326632 144696
rect 325292 143388 325344 143394
rect 325292 143330 325344 143336
rect 325304 130406 325332 143330
rect 326592 133058 326620 144690
rect 358700 144090 358728 153718
rect 327316 144068 327368 144074
rect 327316 144010 327368 144016
rect 358516 144062 358728 144090
rect 327328 143977 327356 144010
rect 327314 143968 327370 143977
rect 327314 143903 327370 143912
rect 327314 141928 327370 141937
rect 327314 141863 327370 141872
rect 330088 141886 331390 141914
rect 332402 141886 332784 141914
rect 327328 141354 327356 141863
rect 327316 141348 327368 141354
rect 327316 141290 327368 141296
rect 326580 133052 326632 133058
rect 326580 132994 326632 133000
rect 325476 131760 325528 131766
rect 325476 131702 325528 131708
rect 325384 130468 325436 130474
rect 325384 130410 325436 130416
rect 325292 130400 325344 130406
rect 325292 130342 325344 130348
rect 325292 122036 325344 122042
rect 325292 121978 325344 121984
rect 325198 98544 325254 98553
rect 325198 98479 325254 98488
rect 324556 95108 324608 95114
rect 324556 95050 324608 95056
rect 324568 95017 324596 95050
rect 324554 95008 324610 95017
rect 324554 94943 324610 94952
rect 325304 92297 325332 121978
rect 325396 110929 325424 130410
rect 325488 113649 325516 131702
rect 326592 119934 326620 132994
rect 326580 119928 326632 119934
rect 326580 119870 326632 119876
rect 325474 113640 325530 113649
rect 325474 113575 325530 113584
rect 325382 110920 325438 110929
rect 325382 110855 325438 110864
rect 325384 108232 325436 108238
rect 325384 108174 325436 108180
rect 325290 92288 325346 92297
rect 325290 92223 325346 92232
rect 325396 88897 325424 108174
rect 325382 88888 325438 88897
rect 325382 88823 325438 88832
rect 326592 86721 326620 119870
rect 330088 95114 330116 141886
rect 332756 131154 332784 141886
rect 333400 139246 333428 141900
rect 333388 139240 333440 139246
rect 333388 139182 333440 139188
rect 334124 139240 334176 139246
rect 334124 139182 334176 139188
rect 332744 131148 332796 131154
rect 332744 131090 332796 131096
rect 334136 131086 334164 139182
rect 334412 138634 334440 141900
rect 335424 141886 335530 141914
rect 336542 141886 336924 141914
rect 337554 141886 338120 141914
rect 334400 138628 334452 138634
rect 334400 138570 334452 138576
rect 334124 131080 334176 131086
rect 334124 131022 334176 131028
rect 335424 131018 335452 141886
rect 335504 138628 335556 138634
rect 335504 138570 335556 138576
rect 335516 131290 335544 138570
rect 335504 131284 335556 131290
rect 335504 131226 335556 131232
rect 336896 131222 336924 141886
rect 338092 131358 338120 141886
rect 338264 138832 338316 138838
rect 338264 138774 338316 138780
rect 338172 138696 338224 138702
rect 338172 138638 338224 138644
rect 338080 131352 338132 131358
rect 338080 131294 338132 131300
rect 336884 131216 336936 131222
rect 336884 131158 336936 131164
rect 335412 131012 335464 131018
rect 335412 130954 335464 130960
rect 338184 130406 338212 138638
rect 337528 130400 337580 130406
rect 337528 130342 337580 130348
rect 338172 130400 338224 130406
rect 338172 130342 338224 130348
rect 337540 128722 337568 130342
rect 338276 130082 338304 138774
rect 338552 138634 338580 141900
rect 339564 141886 339670 141914
rect 340682 141886 341064 141914
rect 338540 138628 338592 138634
rect 338540 138570 338592 138576
rect 339564 131426 339592 141886
rect 339644 138628 339696 138634
rect 339644 138570 339696 138576
rect 339656 131562 339684 138570
rect 339644 131556 339696 131562
rect 339644 131498 339696 131504
rect 341036 131494 341064 141886
rect 341680 138702 341708 141900
rect 341760 138900 341812 138906
rect 341760 138842 341812 138848
rect 341668 138696 341720 138702
rect 341668 138638 341720 138644
rect 341668 131624 341720 131630
rect 341668 131566 341720 131572
rect 341024 131488 341076 131494
rect 341024 131430 341076 131436
rect 339552 131420 339604 131426
rect 339552 131362 339604 131368
rect 341024 131148 341076 131154
rect 341024 131090 341076 131096
rect 340564 130944 340616 130950
rect 340564 130886 340616 130892
rect 338724 130604 338776 130610
rect 338724 130546 338776 130552
rect 338184 130054 338304 130082
rect 338184 128722 338212 130054
rect 338736 128722 338764 130546
rect 339368 130536 339420 130542
rect 339368 130478 339420 130484
rect 339380 128722 339408 130478
rect 339552 130400 339604 130406
rect 339552 130342 339604 130348
rect 337232 128694 337568 128722
rect 337784 128694 338212 128722
rect 338428 128694 338764 128722
rect 339072 128694 339408 128722
rect 339564 128586 339592 130342
rect 340576 128722 340604 130886
rect 341036 128722 341064 131090
rect 341680 128722 341708 131566
rect 341772 130406 341800 138842
rect 342692 138838 342720 141900
rect 342680 138832 342732 138838
rect 342680 138774 342732 138780
rect 341944 138696 341996 138702
rect 341944 138638 341996 138644
rect 341852 138628 341904 138634
rect 341852 138570 341904 138576
rect 341864 130610 341892 138570
rect 341852 130604 341904 130610
rect 341852 130546 341904 130552
rect 341956 130542 341984 138638
rect 343796 138634 343824 141900
rect 344808 138702 344836 141900
rect 345820 138838 345848 141900
rect 346740 141886 346846 141914
rect 347568 141886 347950 141914
rect 348028 141886 348962 141914
rect 345808 138832 345860 138838
rect 345808 138774 345860 138780
rect 344796 138696 344848 138702
rect 344796 138638 344848 138644
rect 343784 138628 343836 138634
rect 343784 138570 343836 138576
rect 346636 136520 346688 136526
rect 346636 136462 346688 136468
rect 343876 135092 343928 135098
rect 343876 135034 343928 135040
rect 343888 134486 343916 135034
rect 343876 134480 343928 134486
rect 343876 134422 343928 134428
rect 343324 132372 343376 132378
rect 343324 132314 343376 132320
rect 343336 131766 343364 132314
rect 343324 131760 343376 131766
rect 343324 131702 343376 131708
rect 342496 130876 342548 130882
rect 342496 130818 342548 130824
rect 342404 130808 342456 130814
rect 342404 130750 342456 130756
rect 341944 130536 341996 130542
rect 341944 130478 341996 130484
rect 341760 130400 341812 130406
rect 341760 130342 341812 130348
rect 342416 128722 342444 130750
rect 340268 128694 340604 128722
rect 340912 128694 341064 128722
rect 341464 128694 341708 128722
rect 342108 128694 342444 128722
rect 342508 128722 342536 130818
rect 343336 128994 343364 131702
rect 343290 128966 343364 128994
rect 342508 128694 342752 128722
rect 343290 128708 343318 128966
rect 343888 128722 343916 134422
rect 343968 133732 344020 133738
rect 343968 133674 344020 133680
rect 343980 133058 344008 133674
rect 343968 133052 344020 133058
rect 343968 132994 344020 133000
rect 344244 133052 344296 133058
rect 344244 132994 344296 133000
rect 344256 128722 344284 132994
rect 346084 132508 346136 132514
rect 346084 132450 346136 132456
rect 346096 131698 346124 132450
rect 346084 131692 346136 131698
rect 346084 131634 346136 131640
rect 345164 130536 345216 130542
rect 345164 130478 345216 130484
rect 345176 128722 345204 130478
rect 345716 130332 345768 130338
rect 345716 130274 345768 130280
rect 343888 128694 343948 128722
rect 344256 128694 344592 128722
rect 345176 128694 345236 128722
rect 345728 128586 345756 130274
rect 346096 128722 346124 131634
rect 346648 131154 346676 136462
rect 346636 131148 346688 131154
rect 346636 131090 346688 131096
rect 346740 130950 346768 141886
rect 347568 136526 347596 141886
rect 347556 136520 347608 136526
rect 347556 136462 347608 136468
rect 347004 135840 347056 135846
rect 347004 135782 347056 135788
rect 346728 130944 346780 130950
rect 346728 130886 346780 130892
rect 347016 128722 347044 135782
rect 348028 131630 348056 141886
rect 349960 138634 349988 141900
rect 350972 139625 351000 141900
rect 352076 139625 352104 141900
rect 352720 141886 353102 141914
rect 353548 141886 354114 141914
rect 355020 141886 355126 141914
rect 355848 141886 356230 141914
rect 356308 141886 357242 141914
rect 357688 141886 358254 141914
rect 350958 139616 351014 139625
rect 350958 139551 351014 139560
rect 352062 139616 352118 139625
rect 352062 139551 352118 139560
rect 348660 138628 348712 138634
rect 348660 138570 348712 138576
rect 349948 138628 350000 138634
rect 349948 138570 350000 138576
rect 348016 131624 348068 131630
rect 348016 131566 348068 131572
rect 348568 131284 348620 131290
rect 348568 131226 348620 131232
rect 348016 131080 348068 131086
rect 348016 131022 348068 131028
rect 347280 130740 347332 130746
rect 347280 130682 347332 130688
rect 347292 128722 347320 130682
rect 348028 128722 348056 131022
rect 348580 128722 348608 131226
rect 348672 130814 348700 138570
rect 350960 131556 351012 131562
rect 350960 131498 351012 131504
rect 350408 131352 350460 131358
rect 350408 131294 350460 131300
rect 349764 131216 349816 131222
rect 349764 131158 349816 131164
rect 349396 131012 349448 131018
rect 349396 130954 349448 130960
rect 348660 130808 348712 130814
rect 348660 130750 348712 130756
rect 349408 128722 349436 130954
rect 349776 128722 349804 131158
rect 350420 128722 350448 131294
rect 350972 128722 351000 131498
rect 352248 131488 352300 131494
rect 352248 131430 352300 131436
rect 351604 131420 351656 131426
rect 351604 131362 351656 131368
rect 351616 128722 351644 131362
rect 352260 128722 352288 131430
rect 346096 128694 346432 128722
rect 347016 128694 347076 128722
rect 347292 128694 347628 128722
rect 348028 128694 348272 128722
rect 348580 128694 348916 128722
rect 349408 128694 349468 128722
rect 349776 128694 350112 128722
rect 350420 128694 350756 128722
rect 350972 128694 351308 128722
rect 351616 128694 351952 128722
rect 352260 128694 352596 128722
rect 339564 128558 339624 128586
rect 345728 128558 345788 128586
rect 334214 122208 334270 122217
rect 334214 122143 334270 122152
rect 334228 122042 334256 122143
rect 334216 122036 334268 122042
rect 334216 121978 334268 121984
rect 334214 108880 334270 108889
rect 334214 108815 334270 108824
rect 334228 108238 334256 108815
rect 334216 108232 334268 108238
rect 334216 108174 334268 108180
rect 352720 101982 352748 141886
rect 353548 107490 353576 141886
rect 354916 132440 354968 132446
rect 354916 132382 354968 132388
rect 354928 117146 354956 132382
rect 354916 117140 354968 117146
rect 354916 117082 354968 117088
rect 353536 107484 353588 107490
rect 353536 107426 353588 107432
rect 352708 101976 352760 101982
rect 352708 101918 352760 101924
rect 334214 95552 334270 95561
rect 334214 95487 334270 95496
rect 330076 95108 330128 95114
rect 330076 95050 330128 95056
rect 329340 94428 329392 94434
rect 329340 94370 329392 94376
rect 326578 86712 326634 86721
rect 326578 86647 326634 86656
rect 329352 86070 329380 94370
rect 324556 86064 324608 86070
rect 324556 86006 324608 86012
rect 329340 86064 329392 86070
rect 329340 86006 329392 86012
rect 324568 85769 324596 86006
rect 324554 85760 324610 85769
rect 324554 85695 324610 85704
rect 328420 76408 328472 76414
rect 328420 76350 328472 76356
rect 328432 75297 328460 76350
rect 330088 75954 330116 95050
rect 334228 94434 334256 95487
rect 334216 94428 334268 94434
rect 334216 94370 334268 94376
rect 337324 88846 337660 88874
rect 338152 88846 338304 88874
rect 338980 88846 339592 88874
rect 339808 88846 340144 88874
rect 340636 88846 340972 88874
rect 341464 88846 341708 88874
rect 342292 88846 342444 88874
rect 343212 88846 343548 88874
rect 344040 88846 344376 88874
rect 344868 88846 345112 88874
rect 336884 87220 336936 87226
rect 336884 87162 336936 87168
rect 334124 87016 334176 87022
rect 334124 86958 334176 86964
rect 332744 86812 332796 86818
rect 332744 86754 332796 86760
rect 330088 75926 330852 75954
rect 330824 75682 330852 75926
rect 332756 75818 332784 86754
rect 334136 79202 334164 86958
rect 335412 86948 335464 86954
rect 335412 86890 335464 86896
rect 335424 79202 335452 86890
rect 335504 86880 335556 86886
rect 335504 86822 335556 86828
rect 333388 79196 333440 79202
rect 333388 79138 333440 79144
rect 334124 79196 334176 79202
rect 334124 79138 334176 79144
rect 334400 79196 334452 79202
rect 334400 79138 334452 79144
rect 335412 79196 335464 79202
rect 335412 79138 335464 79144
rect 332402 75790 332784 75818
rect 333400 75804 333428 79138
rect 334412 75804 334440 79138
rect 335516 75804 335544 86822
rect 336896 75818 336924 87162
rect 337632 86206 337660 88846
rect 338080 87152 338132 87158
rect 338080 87094 338132 87100
rect 337620 86200 337672 86206
rect 337620 86142 337672 86148
rect 338092 85202 338120 87094
rect 338276 86138 338304 88846
rect 339092 86200 339144 86206
rect 339092 86142 339144 86148
rect 338264 86132 338316 86138
rect 338264 86074 338316 86080
rect 339000 86132 339052 86138
rect 339000 86074 339052 86080
rect 338092 85174 338304 85202
rect 338276 79066 338304 85174
rect 339012 79134 339040 86074
rect 339000 79128 339052 79134
rect 339000 79070 339052 79076
rect 337528 79060 337580 79066
rect 337528 79002 337580 79008
rect 338264 79060 338316 79066
rect 338264 79002 338316 79008
rect 336542 75790 336924 75818
rect 337540 75804 337568 79002
rect 339104 78726 339132 86142
rect 339564 79202 339592 88846
rect 339644 87084 339696 87090
rect 339644 87026 339696 87032
rect 339552 79196 339604 79202
rect 339552 79138 339604 79144
rect 339092 78720 339144 78726
rect 339092 78662 339144 78668
rect 338540 78652 338592 78658
rect 338540 78594 338592 78600
rect 338552 75804 338580 78594
rect 339656 75804 339684 87026
rect 340116 86138 340144 88846
rect 340944 87294 340972 88846
rect 340932 87288 340984 87294
rect 340932 87230 340984 87236
rect 341024 87016 341076 87022
rect 341024 86958 341076 86964
rect 340104 86132 340156 86138
rect 340104 86074 340156 86080
rect 341036 75818 341064 86958
rect 341680 86206 341708 88846
rect 341668 86200 341720 86206
rect 341668 86142 341720 86148
rect 342416 86138 342444 88846
rect 343520 87362 343548 88846
rect 343508 87356 343560 87362
rect 343508 87298 343560 87304
rect 344348 86682 344376 88846
rect 344336 86676 344388 86682
rect 344336 86618 344388 86624
rect 345084 86546 345112 88846
rect 345360 88846 345696 88874
rect 346188 88846 346524 88874
rect 347016 88846 347352 88874
rect 348028 88846 348272 88874
rect 348764 88846 349100 88874
rect 349592 88846 349928 88874
rect 350420 88846 350756 88874
rect 351248 88846 351584 88874
rect 352168 88846 352412 88874
rect 345256 87288 345308 87294
rect 345256 87230 345308 87236
rect 345072 86540 345124 86546
rect 345072 86482 345124 86488
rect 344612 86200 344664 86206
rect 344612 86142 344664 86148
rect 341760 86132 341812 86138
rect 341760 86074 341812 86080
rect 342404 86132 342456 86138
rect 342404 86074 342456 86080
rect 344520 86132 344572 86138
rect 344520 86074 344572 86080
rect 341772 79066 341800 86074
rect 344532 79202 344560 86074
rect 343784 79196 343836 79202
rect 343784 79138 343836 79144
rect 344520 79196 344572 79202
rect 344520 79138 344572 79144
rect 342680 79128 342732 79134
rect 342680 79070 342732 79076
rect 341760 79060 341812 79066
rect 341760 79002 341812 79008
rect 341668 78720 341720 78726
rect 341668 78662 341720 78668
rect 340682 75790 341064 75818
rect 341680 75804 341708 78662
rect 342692 75804 342720 79070
rect 343796 75804 343824 79138
rect 344624 79134 344652 86142
rect 344612 79128 344664 79134
rect 344612 79070 344664 79076
rect 344796 79060 344848 79066
rect 344796 79002 344848 79008
rect 344808 75804 344836 79002
rect 345268 75682 345296 87230
rect 345360 86818 345388 88846
rect 346188 86954 346216 88846
rect 346176 86948 346228 86954
rect 346176 86890 346228 86896
rect 345348 86812 345400 86818
rect 345348 86754 345400 86760
rect 347016 86750 347044 88846
rect 348028 86886 348056 88846
rect 348200 87356 348252 87362
rect 348200 87298 348252 87304
rect 348016 86880 348068 86886
rect 348016 86822 348068 86828
rect 347004 86744 347056 86750
rect 347004 86686 347056 86692
rect 347280 86676 347332 86682
rect 347280 86618 347332 86624
rect 345900 86132 345952 86138
rect 345900 86074 345952 86080
rect 345912 78658 345940 86074
rect 347292 79202 347320 86618
rect 347280 79196 347332 79202
rect 347280 79138 347332 79144
rect 346820 79128 346872 79134
rect 346820 79070 346872 79076
rect 347924 79128 347976 79134
rect 347924 79070 347976 79076
rect 345900 78652 345952 78658
rect 345900 78594 345952 78600
rect 346832 75804 346860 79070
rect 347936 75804 347964 79070
rect 348212 75954 348240 87298
rect 348764 87226 348792 88846
rect 348752 87220 348804 87226
rect 348752 87162 348804 87168
rect 349592 87158 349620 88846
rect 349580 87152 349632 87158
rect 349580 87094 349632 87100
rect 350420 86138 350448 88846
rect 351248 87090 351276 88846
rect 351236 87084 351288 87090
rect 351236 87026 351288 87032
rect 352168 87022 352196 88846
rect 352156 87016 352208 87022
rect 352156 86958 352208 86964
rect 350408 86132 350460 86138
rect 350408 86074 350460 86080
rect 349948 79196 350000 79202
rect 349948 79138 350000 79144
rect 348212 75926 348424 75954
rect 348396 75818 348424 75926
rect 348396 75790 348962 75818
rect 349960 75804 349988 79138
rect 350958 77872 351014 77881
rect 350958 77807 351014 77816
rect 352062 77872 352118 77881
rect 352062 77807 352118 77816
rect 350972 75804 351000 77807
rect 352076 75804 352104 77807
rect 352720 75818 352748 101918
rect 352798 97864 352854 97873
rect 352798 97799 352800 97808
rect 352852 97799 352854 97808
rect 352800 97770 352852 97776
rect 352800 92320 352852 92326
rect 352800 92262 352852 92268
rect 352812 90121 352840 92262
rect 352798 90112 352854 90121
rect 352798 90047 352854 90056
rect 352720 75790 353102 75818
rect 353548 75682 353576 107426
rect 354928 84098 354956 117082
rect 355020 112998 355048 141886
rect 355848 132446 355876 141886
rect 355836 132440 355888 132446
rect 355836 132382 355888 132388
rect 356202 126288 356258 126297
rect 356202 126223 356258 126232
rect 356216 126122 356244 126223
rect 356204 126116 356256 126122
rect 356204 126058 356256 126064
rect 356308 122654 356336 141886
rect 357688 126802 357716 141886
rect 357676 126796 357728 126802
rect 357676 126738 357728 126744
rect 356296 122648 356348 122654
rect 356296 122590 356348 122596
rect 356202 121256 356258 121265
rect 356202 121191 356258 121200
rect 356216 120614 356244 121191
rect 356204 120608 356256 120614
rect 356204 120550 356256 120556
rect 356202 116224 356258 116233
rect 356202 116159 356258 116168
rect 356216 115106 356244 116159
rect 356204 115100 356256 115106
rect 356204 115042 356256 115048
rect 355008 112992 355060 112998
rect 355008 112934 355060 112940
rect 354916 84092 354968 84098
rect 354916 84034 354968 84040
rect 355020 75818 355048 112934
rect 356202 111328 356258 111337
rect 356202 111263 356258 111272
rect 356216 110958 356244 111263
rect 356204 110952 356256 110958
rect 356204 110894 356256 110900
rect 356202 106296 356258 106305
rect 356202 106231 356258 106240
rect 356216 105450 356244 106231
rect 356204 105444 356256 105450
rect 356204 105386 356256 105392
rect 356202 101264 356258 101273
rect 356202 101199 356258 101208
rect 356216 100622 356244 101199
rect 356204 100616 356256 100622
rect 356204 100558 356256 100564
rect 356202 96232 356258 96241
rect 356202 96167 356258 96176
rect 356216 95794 356244 96167
rect 356204 95788 356256 95794
rect 356204 95730 356256 95736
rect 356202 91336 356258 91345
rect 356202 91271 356258 91280
rect 356216 90218 356244 91271
rect 356204 90212 356256 90218
rect 356204 90154 356256 90160
rect 355836 84092 355888 84098
rect 355836 84034 355888 84040
rect 355848 75818 355876 84034
rect 355020 75790 355126 75818
rect 355848 75790 356230 75818
rect 356308 75682 356336 122590
rect 357688 75682 357716 126738
rect 358516 124801 358544 144062
rect 359068 135778 359096 168247
rect 360434 165184 360490 165193
rect 360434 165119 360490 165128
rect 359056 135772 359108 135778
rect 359056 135714 359108 135720
rect 360448 132514 360476 165119
rect 360528 162700 360580 162706
rect 360528 162642 360580 162648
rect 360540 162065 360568 162642
rect 360526 162056 360582 162065
rect 360526 161991 360582 162000
rect 360436 132508 360488 132514
rect 360436 132450 360488 132456
rect 360540 130474 360568 161991
rect 360618 158928 360674 158937
rect 360618 158863 360674 158872
rect 360344 130468 360396 130474
rect 360344 130410 360396 130416
rect 360528 130468 360580 130474
rect 360528 130410 360580 130416
rect 360356 130354 360384 130410
rect 360632 130354 360660 158863
rect 360710 155800 360766 155809
rect 360710 155735 360766 155744
rect 360724 133738 360752 155735
rect 360802 152672 360858 152681
rect 360802 152607 360858 152616
rect 360816 135098 360844 152607
rect 360986 149544 361042 149553
rect 360986 149479 361042 149488
rect 360894 146416 360950 146425
rect 360894 146351 360950 146360
rect 360804 135092 360856 135098
rect 360804 135034 360856 135040
rect 360712 133732 360764 133738
rect 360712 133674 360764 133680
rect 360908 130950 360936 146351
rect 361000 132378 361028 149479
rect 361092 143433 361120 221462
rect 361184 181338 361212 224182
rect 361276 214250 361304 237335
rect 362472 233630 362500 371742
rect 429436 366224 429488 366230
rect 429436 366166 429488 366172
rect 429448 365521 429476 366166
rect 429434 365512 429490 365521
rect 429434 365447 429490 365456
rect 430078 353000 430134 353009
rect 430078 352935 430134 352944
rect 429434 340488 429490 340497
rect 429434 340423 429490 340432
rect 429448 340118 429476 340423
rect 374144 340112 374196 340118
rect 374144 340054 374196 340060
rect 429436 340112 429488 340118
rect 429436 340054 429488 340060
rect 365220 326988 365272 326994
rect 365220 326930 365272 326936
rect 364484 239404 364536 239410
rect 364484 239346 364536 239352
rect 362460 233624 362512 233630
rect 362460 233566 362512 233572
rect 362460 222948 362512 222954
rect 362460 222890 362512 222896
rect 361264 214244 361316 214250
rect 361264 214186 361316 214192
rect 361172 181332 361224 181338
rect 361172 181274 361224 181280
rect 361184 155809 361212 181274
rect 361264 165488 361316 165494
rect 361264 165430 361316 165436
rect 361276 165193 361304 165430
rect 361262 165184 361318 165193
rect 361262 165119 361318 165128
rect 361262 158928 361318 158937
rect 361262 158863 361318 158872
rect 361276 158558 361304 158863
rect 361264 158552 361316 158558
rect 361264 158494 361316 158500
rect 361170 155800 361226 155809
rect 361170 155735 361226 155744
rect 361078 143424 361134 143433
rect 361078 143359 361134 143368
rect 360988 132372 361040 132378
rect 360988 132314 361040 132320
rect 360896 130944 360948 130950
rect 360896 130886 360948 130892
rect 360356 130326 360660 130354
rect 361080 130332 361132 130338
rect 358318 124792 358374 124801
rect 358318 124727 358374 124736
rect 358502 124792 358558 124801
rect 358502 124727 358558 124736
rect 358332 108238 358360 124727
rect 358320 108232 358372 108238
rect 358320 108174 358372 108180
rect 358320 108096 358372 108102
rect 358320 108038 358372 108044
rect 358332 105382 358360 108038
rect 358320 105376 358372 105382
rect 358320 105318 358372 105324
rect 358320 95856 358372 95862
rect 358320 95798 358372 95804
rect 358332 88926 358360 95798
rect 358320 88920 358372 88926
rect 358320 88862 358372 88868
rect 358412 88716 358464 88722
rect 358412 88658 358464 88664
rect 358424 86070 358452 88658
rect 360356 87430 360384 130326
rect 361080 130274 361132 130280
rect 361092 87498 361120 130274
rect 361080 87492 361132 87498
rect 361080 87434 361132 87440
rect 359700 87424 359752 87430
rect 359700 87366 359752 87372
rect 360344 87424 360396 87430
rect 360344 87366 360396 87372
rect 358412 86064 358464 86070
rect 358412 86006 358464 86012
rect 358504 76476 358556 76482
rect 358504 76418 358556 76424
rect 330824 75654 331390 75682
rect 345268 75654 345834 75682
rect 353548 75654 354114 75682
rect 356308 75654 357242 75682
rect 357688 75654 358254 75682
rect 328418 75288 328474 75297
rect 328418 75223 328474 75232
rect 328326 74200 328382 74209
rect 328326 74135 328382 74144
rect 328340 73762 328368 74135
rect 328328 73756 328380 73762
rect 328328 73698 328380 73704
rect 327222 72568 327278 72577
rect 327222 72503 327278 72512
rect 327038 71480 327094 71489
rect 327038 71415 327094 71424
rect 327052 67098 327080 71415
rect 327130 69576 327186 69585
rect 327130 69511 327186 69520
rect 327040 67092 327092 67098
rect 327040 67034 327092 67040
rect 326946 66992 327002 67001
rect 326946 66927 327002 66936
rect 326960 63698 326988 66927
rect 327144 66010 327172 69511
rect 327236 69138 327264 72503
rect 328510 71072 328566 71081
rect 328510 71007 328566 71016
rect 328524 70974 328552 71007
rect 328512 70968 328564 70974
rect 328512 70910 328564 70916
rect 358516 69682 358544 76418
rect 358504 69676 358556 69682
rect 358504 69618 358556 69624
rect 358412 69540 358464 69546
rect 358412 69482 358464 69488
rect 327224 69132 327276 69138
rect 327224 69074 327276 69080
rect 327222 68352 327278 68361
rect 327222 68287 327278 68296
rect 327132 66004 327184 66010
rect 327132 65946 327184 65952
rect 327130 65496 327186 65505
rect 327130 65431 327186 65440
rect 326948 63692 327000 63698
rect 326948 63634 327000 63640
rect 327144 62610 327172 65431
rect 327236 64650 327264 68287
rect 328234 67264 328290 67273
rect 328234 67199 328290 67208
rect 327224 64644 327276 64650
rect 327224 64586 327276 64592
rect 327314 64544 327370 64553
rect 327314 64479 327370 64488
rect 327222 62776 327278 62785
rect 327222 62711 327278 62720
rect 327132 62604 327184 62610
rect 327132 62546 327184 62552
rect 327236 58734 327264 62711
rect 327328 61590 327356 64479
rect 328248 64174 328276 67199
rect 328236 64168 328288 64174
rect 328236 64110 328288 64116
rect 328418 63184 328474 63193
rect 328418 63119 328474 63128
rect 327316 61584 327368 61590
rect 327316 61526 327368 61532
rect 328326 61416 328382 61425
rect 328326 61351 328382 61360
rect 327224 58728 327276 58734
rect 327224 58670 327276 58676
rect 327498 58696 327554 58705
rect 327498 58631 327554 58640
rect 327512 56558 327540 58631
rect 328340 58598 328368 61351
rect 328432 60298 328460 63119
rect 328420 60292 328472 60298
rect 328420 60234 328472 60240
rect 328418 60056 328474 60065
rect 328418 59991 328474 60000
rect 328328 58592 328380 58598
rect 328328 58534 328380 58540
rect 328432 57850 328460 59991
rect 358424 59890 358452 69482
rect 358412 59884 358464 59890
rect 358412 59826 358464 59832
rect 358596 59884 358648 59890
rect 358596 59826 358648 59832
rect 328602 58968 328658 58977
rect 328602 58903 328658 58912
rect 328420 57844 328472 57850
rect 328420 57786 328472 57792
rect 328418 57200 328474 57209
rect 328418 57135 328474 57144
rect 327500 56552 327552 56558
rect 327500 56494 327552 56500
rect 327498 55976 327554 55985
rect 327498 55911 327554 55920
rect 327512 54246 327540 55911
rect 328432 55674 328460 57135
rect 328616 56354 328644 58903
rect 328604 56348 328656 56354
rect 328604 56290 328656 56296
rect 328420 55668 328472 55674
rect 328420 55610 328472 55616
rect 328510 55296 328566 55305
rect 328510 55231 328566 55240
rect 328524 55062 328552 55231
rect 328512 55056 328564 55062
rect 328512 54998 328564 55004
rect 328418 54480 328474 54489
rect 328418 54415 328420 54424
rect 328472 54415 328474 54424
rect 328420 54386 328472 54392
rect 327500 54240 327552 54246
rect 327500 54182 327552 54188
rect 328420 53696 328472 53702
rect 328420 53638 328472 53644
rect 328432 53537 328460 53638
rect 328418 53528 328474 53537
rect 328418 53463 328474 53472
rect 328512 52948 328564 52954
rect 328512 52890 328564 52896
rect 328524 52449 328552 52890
rect 328510 52440 328566 52449
rect 328510 52375 328566 52384
rect 323820 51588 323872 51594
rect 323820 51530 323872 51536
rect 327682 50944 327738 50953
rect 327682 50879 327738 50888
rect 327696 50370 327724 50879
rect 358608 50409 358636 59826
rect 328418 50400 328474 50409
rect 327684 50364 327736 50370
rect 328418 50335 328474 50344
rect 358594 50400 358650 50409
rect 358594 50335 358650 50344
rect 327684 50306 327736 50312
rect 328432 50302 328460 50335
rect 328420 50296 328472 50302
rect 328420 50238 328472 50244
rect 328418 49312 328474 49321
rect 328418 49247 328474 49256
rect 328432 48942 328460 49247
rect 328420 48936 328472 48942
rect 328420 48878 328472 48884
rect 327866 47952 327922 47961
rect 327866 47887 327922 47896
rect 327880 47514 327908 47887
rect 327868 47508 327920 47514
rect 327868 47450 327920 47456
rect 332664 45950 332692 47924
rect 322532 45944 322584 45950
rect 322532 45886 322584 45892
rect 332652 45944 332704 45950
rect 332652 45886 332704 45892
rect 336160 45814 336188 47924
rect 338356 47372 338408 47378
rect 338356 47314 338408 47320
rect 338368 46698 338396 47314
rect 339656 46698 339684 47924
rect 338356 46692 338408 46698
rect 338356 46634 338408 46640
rect 339644 46692 339696 46698
rect 339644 46634 339696 46640
rect 336148 45808 336200 45814
rect 336148 45750 336200 45756
rect 324556 45400 324608 45406
rect 324556 45342 324608 45348
rect 317472 44856 317524 44862
rect 317472 44798 317524 44804
rect 317104 37852 317156 37858
rect 317104 37794 317156 37800
rect 314068 37172 314120 37178
rect 314068 37114 314120 37120
rect 314804 37172 314856 37178
rect 314804 37114 314856 37120
rect 312780 36764 312832 36770
rect 312780 36706 312832 36712
rect 314080 34732 314108 37114
rect 317116 35154 317144 37794
rect 317024 35126 317144 35154
rect 317024 34746 317052 35126
rect 316578 34718 317052 34746
rect 299098 34582 299664 34610
rect 276164 33092 276216 33098
rect 276164 33034 276216 33040
rect 276070 26056 276126 26065
rect 276070 25991 276126 26000
rect 275518 23336 275574 23345
rect 275518 23271 275574 23280
rect 276176 20761 276204 33034
rect 276162 20752 276218 20761
rect 276162 20687 276218 20696
rect 273956 16704 274008 16710
rect 273956 16646 274008 16652
rect 265860 12352 265912 12358
rect 265860 12294 265912 12300
rect 273968 9304 273996 16646
rect 280408 12426 280436 18956
rect 285376 16778 285404 18956
rect 290068 18942 290358 18970
rect 285364 16772 285416 16778
rect 285364 16714 285416 16720
rect 290068 12494 290096 18942
rect 295404 16710 295432 18956
rect 299716 16772 299768 16778
rect 299716 16714 299768 16720
rect 295392 16704 295444 16710
rect 295392 16646 295444 16652
rect 286836 12488 286888 12494
rect 286836 12430 286888 12436
rect 290056 12488 290108 12494
rect 290056 12430 290108 12436
rect 280396 12420 280448 12426
rect 280396 12362 280448 12368
rect 286848 9304 286876 12430
rect 299728 9304 299756 16714
rect 300372 16642 300400 18956
rect 300360 16636 300412 16642
rect 300360 16578 300412 16584
rect 305340 16574 305368 18956
rect 305328 16568 305380 16574
rect 305328 16510 305380 16516
rect 310400 16506 310428 18956
rect 310388 16500 310440 16506
rect 310388 16442 310440 16448
rect 315368 16438 315396 18956
rect 315356 16432 315408 16438
rect 315356 16374 315408 16380
rect 312596 12420 312648 12426
rect 312596 12362 312648 12368
rect 312608 9304 312636 12362
rect 324568 9434 324596 45342
rect 324556 9428 324608 9434
rect 324556 9370 324608 9376
rect 325476 9428 325528 9434
rect 325476 9370 325528 9376
rect 325488 9304 325516 9370
rect 338368 9304 338396 46634
rect 343152 46057 343180 47924
rect 343138 46048 343194 46057
rect 343138 45983 343194 45992
rect 346648 45406 346676 47924
rect 350144 46086 350172 47924
rect 353640 47446 353668 47924
rect 353628 47440 353680 47446
rect 353628 47382 353680 47388
rect 350132 46080 350184 46086
rect 350132 46022 350184 46028
rect 357136 45882 357164 47924
rect 358502 47544 358558 47553
rect 358502 47479 358558 47488
rect 358516 47394 358544 47479
rect 358424 47366 358544 47394
rect 357124 45876 357176 45882
rect 357124 45818 357176 45824
rect 347924 45808 347976 45814
rect 347924 45750 347976 45756
rect 347936 45406 347964 45750
rect 357136 45406 357164 45818
rect 346636 45400 346688 45406
rect 346636 45342 346688 45348
rect 347924 45400 347976 45406
rect 347924 45342 347976 45348
rect 357124 45400 357176 45406
rect 357124 45342 357176 45348
rect 358424 40646 358452 47366
rect 359712 45814 359740 87366
rect 361092 46086 361120 87434
rect 362472 86546 362500 222890
rect 362460 86540 362512 86546
rect 362460 86482 362512 86488
rect 361080 46080 361132 46086
rect 361080 46022 361132 46028
rect 359700 45808 359752 45814
rect 359700 45750 359752 45756
rect 358412 40640 358464 40646
rect 358412 40582 358464 40588
rect 358412 37852 358464 37858
rect 358412 37794 358464 37800
rect 358424 30938 358452 37794
rect 358240 30910 358452 30938
rect 358240 28134 358268 30910
rect 358228 28128 358280 28134
rect 358228 28070 358280 28076
rect 358320 18540 358372 18546
rect 358320 18482 358372 18488
rect 358332 12970 358360 18482
rect 351236 12964 351288 12970
rect 351236 12906 351288 12912
rect 358320 12964 358372 12970
rect 358320 12906 358372 12912
rect 351248 9304 351276 12906
rect 364496 9450 364524 239346
rect 365232 233426 365260 326930
rect 367980 274492 368032 274498
rect 367980 274434 368032 274440
rect 369912 274492 369964 274498
rect 369912 274434 369964 274440
rect 365220 233420 365272 233426
rect 365220 233362 365272 233368
rect 365220 218732 365272 218738
rect 365220 218674 365272 218680
rect 365232 138770 365260 218674
rect 367992 213337 368020 274434
rect 369544 263408 369596 263414
rect 369544 263350 369596 263356
rect 369174 236584 369230 236593
rect 369174 236519 369230 236528
rect 368716 235120 368768 235126
rect 368716 235062 368768 235068
rect 368728 234145 368756 235062
rect 368714 234136 368770 234145
rect 368714 234071 368770 234080
rect 368716 233760 368768 233766
rect 368714 233728 368716 233737
rect 368768 233728 368770 233737
rect 368714 233663 368770 233672
rect 368808 233624 368860 233630
rect 368808 233566 368860 233572
rect 368820 233465 368848 233566
rect 368806 233456 368862 233465
rect 368716 233420 368768 233426
rect 368806 233391 368862 233400
rect 368716 233362 368768 233368
rect 368728 233057 368756 233362
rect 368714 233048 368770 233057
rect 368714 232983 368770 232992
rect 368900 232400 368952 232406
rect 368900 232342 368952 232348
rect 368716 232332 368768 232338
rect 368716 232274 368768 232280
rect 368728 232241 368756 232274
rect 368808 232264 368860 232270
rect 368714 232232 368770 232241
rect 368808 232206 368860 232212
rect 368714 232167 368770 232176
rect 368820 231833 368848 232206
rect 368806 231824 368862 231833
rect 368806 231759 368862 231768
rect 368912 231425 368940 232342
rect 368898 231416 368954 231425
rect 368898 231351 368954 231360
rect 368806 231008 368862 231017
rect 368806 230943 368862 230952
rect 368900 230972 368952 230978
rect 368716 230904 368768 230910
rect 368716 230846 368768 230852
rect 368728 230609 368756 230846
rect 368820 230842 368848 230943
rect 368900 230914 368952 230920
rect 368808 230836 368860 230842
rect 368808 230778 368860 230784
rect 368714 230600 368770 230609
rect 368714 230535 368770 230544
rect 368912 230201 368940 230914
rect 368898 230192 368954 230201
rect 368898 230127 368954 230136
rect 368716 229612 368768 229618
rect 368716 229554 368768 229560
rect 368728 229521 368756 229554
rect 368714 229512 368770 229521
rect 368714 229447 368770 229456
rect 368806 229104 368862 229113
rect 368806 229039 368862 229048
rect 368714 228696 368770 228705
rect 368714 228631 368770 228640
rect 368728 228462 368756 228631
rect 368716 228456 368768 228462
rect 368716 228398 368768 228404
rect 368820 228394 368848 229039
rect 368808 228388 368860 228394
rect 368808 228330 368860 228336
rect 368716 228320 368768 228326
rect 368714 228288 368716 228297
rect 368768 228288 368770 228297
rect 368714 228223 368770 228232
rect 368806 227472 368862 227481
rect 368806 227407 368862 227416
rect 368714 227064 368770 227073
rect 368714 226999 368770 227008
rect 368728 226898 368756 226999
rect 368820 226966 368848 227407
rect 368808 226960 368860 226966
rect 368808 226902 368860 226908
rect 368716 226892 368768 226898
rect 368716 226834 368768 226840
rect 369082 226520 369138 226529
rect 369082 226455 369138 226464
rect 368898 226384 368954 226393
rect 368898 226319 368954 226328
rect 368806 225976 368862 225985
rect 368806 225911 368862 225920
rect 368820 225674 368848 225911
rect 368808 225668 368860 225674
rect 368808 225610 368860 225616
rect 368716 225600 368768 225606
rect 368714 225568 368716 225577
rect 368768 225568 368770 225577
rect 368912 225538 368940 226319
rect 368714 225503 368770 225512
rect 368900 225532 368952 225538
rect 368900 225474 368952 225480
rect 368716 225396 368768 225402
rect 368716 225338 368768 225344
rect 368728 224761 368756 225338
rect 368992 225328 369044 225334
rect 368992 225270 369044 225276
rect 368806 225160 368862 225169
rect 368806 225095 368862 225104
rect 368714 224752 368770 224761
rect 368714 224687 368770 224696
rect 368820 224178 368848 225095
rect 368898 224344 368954 224353
rect 368898 224279 368954 224288
rect 368808 224172 368860 224178
rect 368808 224114 368860 224120
rect 368912 224058 368940 224279
rect 368728 224030 368940 224058
rect 368728 223378 368756 224030
rect 368806 223936 368862 223945
rect 368806 223871 368862 223880
rect 368636 223350 368756 223378
rect 368636 222698 368664 223350
rect 368714 223256 368770 223265
rect 368714 223191 368770 223200
rect 368728 222886 368756 223191
rect 368716 222880 368768 222886
rect 368716 222822 368768 222828
rect 368820 222818 368848 223871
rect 368808 222812 368860 222818
rect 368808 222754 368860 222760
rect 368636 222670 368756 222698
rect 368728 221746 368756 222670
rect 368806 222440 368862 222449
rect 368806 222375 368862 222384
rect 368636 221718 368756 221746
rect 368636 214810 368664 221718
rect 368714 221624 368770 221633
rect 368714 221559 368770 221568
rect 368728 221390 368756 221559
rect 368820 221458 368848 222375
rect 368808 221452 368860 221458
rect 368808 221394 368860 221400
rect 368716 221384 368768 221390
rect 368716 221326 368768 221332
rect 369004 221338 369032 225270
rect 369096 224042 369124 226455
rect 369188 224178 369216 236519
rect 369450 236176 369506 236185
rect 369450 236111 369506 236120
rect 369268 227572 369320 227578
rect 369268 227514 369320 227520
rect 369176 224172 369228 224178
rect 369176 224114 369228 224120
rect 369280 224058 369308 227514
rect 369084 224036 369136 224042
rect 369084 223978 369136 223984
rect 369188 224030 369308 224058
rect 369360 224036 369412 224042
rect 369084 222948 369136 222954
rect 369084 222890 369136 222896
rect 369096 222857 369124 222890
rect 369082 222848 369138 222857
rect 369082 222783 369138 222792
rect 369082 222032 369138 222041
rect 369082 221967 369138 221976
rect 369096 221526 369124 221967
rect 369084 221520 369136 221526
rect 369084 221462 369136 221468
rect 369004 221310 369124 221338
rect 368990 221216 369046 221225
rect 368990 221151 369046 221160
rect 368806 220808 368862 220817
rect 368806 220743 368862 220752
rect 368820 220574 368848 220743
rect 368808 220568 368860 220574
rect 368808 220510 368860 220516
rect 368716 220500 368768 220506
rect 368716 220442 368768 220448
rect 368728 220409 368756 220442
rect 368714 220400 368770 220409
rect 368714 220335 368770 220344
rect 369004 220098 369032 221151
rect 368992 220092 369044 220098
rect 368992 220034 369044 220040
rect 368714 219720 368770 219729
rect 368714 219655 368770 219664
rect 368728 218670 368756 219655
rect 368990 219312 369046 219321
rect 368990 219247 369046 219256
rect 368806 218904 368862 218913
rect 368806 218839 368862 218848
rect 368820 218738 368848 218839
rect 368808 218732 368860 218738
rect 368808 218674 368860 218680
rect 368716 218664 368768 218670
rect 368716 218606 368768 218612
rect 368808 218596 368860 218602
rect 368808 218538 368860 218544
rect 368714 218088 368770 218097
rect 368714 218023 368770 218032
rect 368728 217242 368756 218023
rect 368820 217281 368848 218538
rect 368806 217272 368862 217281
rect 368716 217236 368768 217242
rect 368806 217207 368862 217216
rect 368716 217178 368768 217184
rect 368716 217100 368768 217106
rect 368716 217042 368768 217048
rect 368728 216193 368756 217042
rect 369004 216601 369032 219247
rect 369096 217689 369124 221310
rect 369082 217680 369138 217689
rect 369082 217615 369138 217624
rect 369082 217544 369138 217553
rect 369082 217479 369138 217488
rect 368990 216592 369046 216601
rect 368990 216527 369046 216536
rect 368992 216488 369044 216494
rect 368992 216430 369044 216436
rect 368714 216184 368770 216193
rect 368714 216119 368770 216128
rect 368716 215808 368768 215814
rect 368714 215776 368716 215785
rect 368768 215776 368770 215785
rect 368714 215711 368770 215720
rect 368808 215740 368860 215746
rect 368808 215682 368860 215688
rect 368716 215672 368768 215678
rect 368716 215614 368768 215620
rect 368728 214969 368756 215614
rect 368714 214960 368770 214969
rect 368714 214895 368770 214904
rect 368636 214782 368756 214810
rect 368728 214402 368756 214782
rect 368820 214561 368848 215682
rect 368806 214552 368862 214561
rect 369004 214522 369032 216430
rect 368806 214487 368862 214496
rect 368992 214516 369044 214522
rect 368992 214458 369044 214464
rect 368728 214374 368848 214402
rect 368716 214312 368768 214318
rect 368716 214254 368768 214260
rect 368728 213745 368756 214254
rect 368714 213736 368770 213745
rect 368714 213671 368770 213680
rect 367978 213328 368034 213337
rect 367978 213263 368034 213272
rect 368716 213088 368768 213094
rect 368714 213056 368716 213065
rect 368768 213056 368770 213065
rect 368714 212991 368770 213000
rect 368820 195278 368848 214374
rect 368900 214244 368952 214250
rect 368900 214186 368952 214192
rect 368912 214153 368940 214186
rect 368898 214144 368954 214153
rect 368898 214079 368954 214088
rect 369096 207330 369124 217479
rect 369188 215377 369216 224030
rect 369360 223978 369412 223984
rect 369266 219992 369322 220001
rect 369266 219927 369322 219936
rect 369174 215368 369230 215377
rect 369174 215303 369230 215312
rect 369176 214516 369228 214522
rect 369176 214458 369228 214464
rect 369004 207302 369124 207330
rect 369004 204730 369032 207302
rect 369188 207194 369216 214458
rect 369096 207166 369216 207194
rect 368992 204724 369044 204730
rect 368992 204666 369044 204672
rect 368808 195272 368860 195278
rect 368808 195214 368860 195220
rect 369096 195210 369124 207166
rect 369176 204724 369228 204730
rect 369176 204666 369228 204672
rect 369084 195204 369136 195210
rect 369084 195146 369136 195152
rect 368716 192416 368768 192422
rect 368716 192358 368768 192364
rect 368728 185554 368756 192358
rect 368992 190308 369044 190314
rect 368992 190250 369044 190256
rect 368716 185548 368768 185554
rect 368716 185490 368768 185496
rect 368808 185412 368860 185418
rect 368808 185354 368860 185360
rect 368820 182714 368848 185354
rect 368728 182686 368848 182714
rect 368728 177938 368756 182686
rect 369004 179978 369032 190250
rect 368992 179972 369044 179978
rect 368992 179914 369044 179920
rect 369188 179858 369216 204666
rect 369004 179830 369216 179858
rect 368532 177932 368584 177938
rect 368532 177874 368584 177880
rect 368716 177932 368768 177938
rect 368716 177874 368768 177880
rect 368544 173081 368572 177874
rect 368530 173072 368586 173081
rect 368530 173007 368586 173016
rect 368714 173072 368770 173081
rect 368714 173007 368770 173016
rect 368728 168214 368756 173007
rect 369004 168554 369032 179830
rect 369280 168622 369308 219927
rect 369372 216873 369400 223978
rect 369358 216864 369414 216873
rect 369358 216799 369414 216808
rect 369360 195204 369412 195210
rect 369360 195146 369412 195152
rect 369372 190314 369400 195146
rect 369360 190308 369412 190314
rect 369360 190250 369412 190256
rect 369360 179972 369412 179978
rect 369360 179914 369412 179920
rect 369268 168616 369320 168622
rect 369268 168558 369320 168564
rect 368992 168548 369044 168554
rect 368992 168490 369044 168496
rect 368716 168208 368768 168214
rect 368716 168150 368768 168156
rect 368992 168208 369044 168214
rect 368992 168150 369044 168156
rect 369004 153866 369032 168150
rect 368532 153860 368584 153866
rect 368532 153802 368584 153808
rect 368992 153860 369044 153866
rect 368992 153802 369044 153808
rect 368544 152370 368572 153802
rect 368532 152364 368584 152370
rect 368532 152306 368584 152312
rect 368716 152364 368768 152370
rect 368716 152306 368768 152312
rect 365220 138764 365272 138770
rect 365220 138706 365272 138712
rect 368728 137018 368756 152306
rect 368728 136990 368940 137018
rect 368912 132310 368940 136990
rect 368900 132304 368952 132310
rect 368900 132246 368952 132252
rect 369176 54308 369228 54314
rect 369176 54250 369228 54256
rect 369188 45746 369216 54250
rect 369176 45740 369228 45746
rect 369176 45682 369228 45688
rect 369372 35018 369400 179914
rect 369188 34990 369400 35018
rect 369188 32962 369216 34990
rect 369464 33030 369492 236111
rect 369556 229929 369584 263350
rect 369728 262660 369780 262666
rect 369728 262602 369780 262608
rect 369634 235768 369690 235777
rect 369634 235703 369690 235712
rect 369542 229920 369598 229929
rect 369542 229855 369598 229864
rect 369542 227880 369598 227889
rect 369542 227815 369598 227824
rect 369556 209694 369584 227815
rect 369544 209688 369596 209694
rect 369544 209630 369596 209636
rect 369544 199964 369596 199970
rect 369544 199906 369596 199912
rect 369556 190314 369584 199906
rect 369544 190308 369596 190314
rect 369544 190250 369596 190256
rect 369544 179972 369596 179978
rect 369544 179914 369596 179920
rect 369556 54314 369584 179914
rect 369544 54308 369596 54314
rect 369544 54250 369596 54256
rect 369648 33098 369676 235703
rect 369740 232649 369768 262602
rect 369818 235360 369874 235369
rect 369818 235295 369874 235304
rect 369726 232640 369782 232649
rect 369726 232575 369782 232584
rect 369832 228938 369860 235295
rect 369924 234553 369952 274434
rect 374156 236706 374184 340054
rect 429436 319984 429488 319990
rect 429436 319926 429488 319932
rect 405976 315904 406028 315910
rect 405974 315872 405976 315881
rect 406028 315872 406030 315881
rect 405974 315807 406030 315816
rect 429448 315473 429476 319926
rect 429434 315464 429490 315473
rect 429434 315399 429490 315408
rect 427318 313832 427374 313841
rect 405976 313796 406028 313802
rect 427318 313767 427374 313776
rect 405976 313738 406028 313744
rect 405988 313705 406016 313738
rect 405974 313696 406030 313705
rect 405974 313631 406030 313640
rect 405974 310432 406030 310441
rect 405974 310367 406030 310376
rect 405988 310334 406016 310367
rect 405976 310328 406028 310334
rect 405976 310270 406028 310276
rect 405976 308288 406028 308294
rect 405974 308256 405976 308265
rect 406028 308256 406030 308265
rect 405974 308191 406030 308200
rect 406068 306248 406120 306254
rect 406066 306216 406068 306225
rect 406120 306216 406122 306225
rect 406066 306151 406122 306160
rect 405976 304140 406028 304146
rect 405976 304082 406028 304088
rect 405988 303641 406016 304082
rect 405974 303632 406030 303641
rect 405974 303567 406030 303576
rect 405976 300672 406028 300678
rect 405976 300614 406028 300620
rect 405988 300513 406016 300614
rect 405974 300504 406030 300513
rect 405974 300439 406030 300448
rect 405976 298632 406028 298638
rect 405976 298574 406028 298580
rect 405988 298337 406016 298574
rect 405974 298328 406030 298337
rect 405974 298263 406030 298272
rect 405974 295472 406030 295481
rect 405974 295407 406030 295416
rect 405988 295170 406016 295407
rect 405976 295164 406028 295170
rect 405976 295106 406028 295112
rect 405976 293804 406028 293810
rect 405976 293746 406028 293752
rect 405988 293713 406016 293746
rect 405974 293704 406030 293713
rect 405974 293639 406030 293648
rect 405976 291016 406028 291022
rect 405976 290958 406028 290964
rect 405988 290721 406016 290958
rect 405974 290712 406030 290721
rect 405974 290647 406030 290656
rect 427226 289080 427282 289089
rect 427226 289015 427228 289024
rect 427280 289015 427282 289024
rect 427228 288986 427280 288992
rect 406068 288976 406120 288982
rect 406068 288918 406120 288924
rect 406080 288681 406108 288918
rect 406066 288672 406122 288681
rect 406066 288607 406122 288616
rect 405974 285544 406030 285553
rect 405974 285479 405976 285488
rect 406028 285479 406030 285488
rect 405976 285450 406028 285456
rect 405976 283468 406028 283474
rect 405976 283410 406028 283416
rect 405988 283377 406016 283410
rect 405974 283368 406030 283377
rect 405974 283303 406030 283312
rect 405976 279320 406028 279326
rect 405976 279262 406028 279268
rect 405988 278753 406016 279262
rect 405974 278744 406030 278753
rect 405974 278679 406030 278688
rect 410220 274498 410248 276948
rect 410208 274492 410260 274498
rect 410208 274434 410260 274440
rect 385276 262592 385328 262598
rect 385276 262534 385328 262540
rect 377824 239404 377876 239410
rect 377824 239346 377876 239352
rect 373894 236678 374184 236706
rect 377836 236692 377864 239346
rect 381872 239336 381924 239342
rect 381872 239278 381924 239284
rect 381884 236692 381912 239278
rect 385288 236842 385316 262534
rect 412888 249610 412916 276948
rect 414268 276934 415570 276962
rect 417028 276934 418238 276962
rect 419788 276934 420906 276962
rect 422548 276934 423574 276962
rect 414268 253078 414296 276934
rect 417028 256546 417056 276934
rect 419788 259334 419816 276934
rect 422548 262054 422576 276934
rect 422536 262048 422588 262054
rect 422536 261990 422588 261996
rect 419776 259328 419828 259334
rect 419776 259270 419828 259276
rect 417016 256540 417068 256546
rect 417016 256482 417068 256488
rect 414256 253072 414308 253078
rect 414256 253014 414308 253020
rect 412876 249604 412928 249610
rect 412876 249546 412928 249552
rect 389876 240016 389928 240022
rect 389876 239958 389928 239964
rect 385288 236814 385592 236842
rect 385564 236706 385592 236814
rect 385564 236678 385854 236706
rect 389888 236692 389916 239958
rect 393832 239948 393884 239954
rect 393832 239890 393884 239896
rect 393844 236692 393872 239890
rect 370002 234952 370058 234961
rect 370002 234887 370058 234896
rect 369910 234544 369966 234553
rect 369910 234479 369966 234488
rect 370016 229074 370044 234887
rect 370004 229068 370056 229074
rect 370004 229010 370056 229016
rect 369820 228932 369872 228938
rect 369820 228874 369872 228880
rect 370004 228932 370056 228938
rect 370004 228874 370056 228880
rect 369726 226656 369782 226665
rect 369726 226591 369782 226600
rect 369740 46018 369768 226591
rect 369818 223528 369874 223537
rect 369818 223463 369874 223472
rect 369728 46012 369780 46018
rect 369728 45954 369780 45960
rect 369832 45950 369860 223463
rect 369912 221384 369964 221390
rect 369912 221326 369964 221332
rect 369924 211666 369952 221326
rect 369912 211660 369964 211666
rect 369912 211602 369964 211608
rect 369912 209688 369964 209694
rect 369912 209630 369964 209636
rect 369924 199970 369952 209630
rect 369912 199964 369964 199970
rect 369912 199906 369964 199912
rect 369912 190308 369964 190314
rect 369912 190250 369964 190256
rect 369924 179978 369952 190250
rect 369912 179972 369964 179978
rect 369912 179914 369964 179920
rect 370016 87362 370044 228874
rect 406618 221624 406674 221633
rect 406618 221559 406674 221568
rect 405974 218768 406030 218777
rect 405974 218703 406030 218712
rect 405988 218670 406016 218703
rect 394844 218664 394896 218670
rect 394844 218606 394896 218612
rect 405976 218664 406028 218670
rect 405976 218606 406028 218612
rect 370094 218496 370150 218505
rect 370094 218431 370150 218440
rect 370108 217553 370136 218431
rect 370094 217544 370150 217553
rect 370094 217479 370150 217488
rect 394856 213978 394884 218606
rect 405974 214144 406030 214153
rect 405974 214079 405976 214088
rect 406028 214079 406030 214088
rect 405976 214050 406028 214056
rect 406632 214046 406660 221559
rect 427332 215814 427360 313767
rect 428698 308664 428754 308673
rect 428698 308599 428754 308608
rect 427410 304176 427466 304185
rect 427410 304111 427466 304120
rect 427424 240634 427452 304111
rect 427502 298736 427558 298745
rect 427502 298671 427558 298680
rect 427516 253078 427544 298671
rect 427594 293704 427650 293713
rect 427594 293639 427650 293648
rect 427608 265522 427636 293639
rect 427688 290404 427740 290410
rect 427688 290346 427740 290352
rect 427700 284329 427728 290346
rect 427686 284320 427742 284329
rect 427686 284255 427742 284264
rect 427872 280680 427924 280686
rect 427872 280622 427924 280628
rect 427884 279433 427912 280622
rect 427870 279424 427926 279433
rect 427870 279359 427926 279368
rect 427596 265516 427648 265522
rect 427596 265458 427648 265464
rect 427504 253072 427556 253078
rect 427504 253014 427556 253020
rect 427412 240628 427464 240634
rect 427412 240570 427464 240576
rect 428712 227889 428740 308599
rect 429434 290440 429490 290449
rect 429434 290375 429436 290384
rect 429488 290375 429490 290384
rect 429436 290346 429488 290352
rect 430092 269670 430120 352935
rect 430170 327976 430226 327985
rect 430170 327911 430226 327920
rect 430184 314482 430212 327911
rect 430172 314476 430224 314482
rect 430172 314418 430224 314424
rect 430170 302952 430226 302961
rect 430170 302887 430226 302896
rect 430184 280686 430212 302887
rect 430264 289044 430316 289050
rect 430264 288986 430316 288992
rect 430172 280680 430224 280686
rect 430172 280622 430224 280628
rect 430276 277937 430304 288986
rect 430262 277928 430318 277937
rect 430262 277863 430318 277872
rect 430080 269664 430132 269670
rect 430080 269606 430132 269612
rect 429436 265516 429488 265522
rect 429436 265458 429488 265464
rect 429448 265425 429476 265458
rect 429434 265416 429490 265425
rect 429434 265351 429490 265360
rect 429436 253072 429488 253078
rect 429436 253014 429488 253020
rect 429448 252913 429476 253014
rect 429434 252904 429490 252913
rect 429434 252839 429490 252848
rect 429528 240628 429580 240634
rect 429528 240570 429580 240576
rect 429540 240401 429568 240570
rect 429526 240392 429582 240401
rect 429526 240327 429582 240336
rect 428698 227880 428754 227889
rect 428698 227815 428754 227824
rect 427410 220264 427466 220273
rect 427410 220199 427466 220208
rect 427320 215808 427372 215814
rect 427320 215750 427372 215756
rect 406620 214040 406672 214046
rect 406620 213982 406672 213988
rect 394844 213972 394896 213978
rect 394844 213914 394896 213920
rect 370740 211660 370792 211666
rect 370740 211602 370792 211608
rect 370752 181270 370780 211602
rect 383908 210918 383936 212892
rect 405974 211016 406030 211025
rect 405974 210951 405976 210960
rect 406028 210951 406030 210960
rect 405976 210922 406028 210928
rect 383896 210912 383948 210918
rect 383896 210854 383948 210860
rect 385184 210912 385236 210918
rect 385184 210854 385236 210860
rect 370740 181264 370792 181270
rect 370740 181206 370792 181212
rect 370004 87356 370056 87362
rect 370004 87298 370056 87304
rect 369820 45944 369872 45950
rect 369820 45886 369872 45892
rect 376996 45400 377048 45406
rect 376996 45342 377048 45348
rect 369636 33092 369688 33098
rect 369636 33034 369688 33040
rect 369452 33024 369504 33030
rect 369452 32966 369504 32972
rect 369176 32956 369228 32962
rect 369176 32898 369228 32904
rect 364128 9422 364524 9450
rect 364128 9304 364156 9422
rect 377008 9304 377036 45342
rect 385196 12154 385224 210854
rect 427318 210200 427374 210209
rect 427318 210135 427374 210144
rect 405976 209620 406028 209626
rect 405976 209562 406028 209568
rect 405988 209529 406016 209562
rect 405974 209520 406030 209529
rect 405974 209455 406030 209464
rect 405976 206832 406028 206838
rect 405974 206800 405976 206809
rect 406028 206800 406030 206809
rect 405974 206735 406030 206744
rect 406068 204792 406120 204798
rect 406068 204734 406120 204740
rect 406080 204633 406108 204734
rect 406066 204624 406122 204633
rect 406066 204559 406122 204568
rect 405974 201360 406030 201369
rect 405974 201295 405976 201304
rect 406028 201295 406030 201304
rect 405976 201266 406028 201272
rect 427134 200272 427190 200281
rect 427134 200207 427190 200216
rect 427148 199766 427176 200207
rect 427136 199760 427188 199766
rect 427136 199702 427188 199708
rect 405976 199284 406028 199290
rect 405976 199226 406028 199232
rect 405988 199193 406016 199226
rect 405974 199184 406030 199193
rect 405974 199119 406030 199128
rect 405974 195920 406030 195929
rect 405974 195855 406030 195864
rect 405988 195822 406016 195855
rect 405976 195816 406028 195822
rect 405976 195758 406028 195764
rect 406068 195136 406120 195142
rect 406068 195078 406120 195084
rect 406080 194569 406108 195078
rect 406066 194560 406122 194569
rect 406066 194495 406122 194504
rect 405974 191704 406030 191713
rect 405974 191639 405976 191648
rect 406028 191639 406030 191648
rect 405976 191610 406028 191616
rect 405976 189628 406028 189634
rect 405976 189570 406028 189576
rect 405988 189537 406016 189570
rect 405974 189528 406030 189537
rect 405974 189463 406030 189472
rect 405974 186264 406030 186273
rect 405974 186199 406030 186208
rect 405988 186166 406016 186199
rect 405976 186160 406028 186166
rect 405976 186102 406028 186108
rect 427228 185480 427280 185486
rect 427226 185448 427228 185457
rect 427280 185448 427282 185457
rect 427226 185383 427282 185392
rect 405976 184052 406028 184058
rect 405976 183994 406028 184000
rect 405988 183961 406016 183994
rect 405974 183952 406030 183961
rect 405974 183887 406030 183896
rect 410220 181270 410248 182836
rect 412888 181338 412916 182836
rect 412876 181332 412928 181338
rect 412876 181274 412928 181280
rect 410208 181264 410260 181270
rect 410208 181206 410260 181212
rect 415556 158558 415584 182836
rect 418224 162706 418252 182836
rect 420892 165494 420920 182836
rect 423574 182822 423680 182850
rect 423652 168894 423680 182822
rect 423640 168888 423692 168894
rect 423640 168830 423692 168836
rect 420880 165488 420932 165494
rect 420880 165430 420932 165436
rect 418212 162700 418264 162706
rect 418212 162642 418264 162648
rect 415544 158552 415596 158558
rect 415544 158494 415596 158500
rect 427332 140810 427360 210135
rect 427320 140804 427372 140810
rect 427320 140746 427372 140752
rect 405974 126968 406030 126977
rect 405974 126903 406030 126912
rect 405988 126802 406016 126903
rect 405976 126796 406028 126802
rect 405976 126738 406028 126744
rect 427318 126288 427374 126297
rect 427318 126223 427374 126232
rect 405976 126116 406028 126122
rect 405976 126058 406028 126064
rect 405988 125617 406016 126058
rect 405974 125608 406030 125617
rect 405974 125543 406030 125552
rect 405976 122648 406028 122654
rect 405974 122616 405976 122625
rect 406028 122616 406030 122625
rect 405974 122551 406030 122560
rect 405976 120608 406028 120614
rect 405974 120576 405976 120585
rect 406028 120576 406030 120585
rect 405974 120511 406030 120520
rect 405974 117448 406030 117457
rect 405974 117383 406030 117392
rect 405988 117146 406016 117383
rect 405976 117140 406028 117146
rect 405976 117082 406028 117088
rect 405976 115100 406028 115106
rect 405976 115042 406028 115048
rect 405988 114873 406016 115042
rect 405974 114864 406030 114873
rect 405974 114799 406030 114808
rect 405976 112992 406028 112998
rect 405976 112934 406028 112940
rect 405988 112697 406016 112934
rect 405974 112688 406030 112697
rect 405974 112623 406030 112632
rect 406068 110952 406120 110958
rect 406068 110894 406120 110900
rect 406080 110657 406108 110894
rect 406066 110648 406122 110657
rect 406066 110583 406122 110592
rect 405974 107656 406030 107665
rect 405974 107591 406030 107600
rect 405988 107490 406016 107591
rect 405976 107484 406028 107490
rect 405976 107426 406028 107432
rect 405976 105444 406028 105450
rect 405976 105386 406028 105392
rect 405988 105353 406016 105386
rect 405974 105344 406030 105353
rect 405974 105279 406030 105288
rect 405974 102216 406030 102225
rect 405974 102151 406030 102160
rect 405988 101982 406016 102151
rect 405976 101976 406028 101982
rect 405976 101918 406028 101924
rect 405976 100616 406028 100622
rect 405974 100584 405976 100593
rect 406028 100584 406030 100593
rect 405974 100519 406030 100528
rect 405976 97828 406028 97834
rect 405976 97770 406028 97776
rect 405988 97737 406016 97770
rect 405974 97728 406030 97737
rect 405974 97663 406030 97672
rect 427226 96232 427282 96241
rect 427226 96167 427282 96176
rect 427240 95862 427268 96167
rect 427228 95856 427280 95862
rect 427228 95798 427280 95804
rect 405976 95788 406028 95794
rect 405976 95730 406028 95736
rect 405988 95561 406016 95730
rect 405974 95552 406030 95561
rect 405974 95487 406030 95496
rect 405974 92424 406030 92433
rect 405974 92359 406030 92368
rect 405988 92326 406016 92359
rect 405976 92320 406028 92326
rect 405976 92262 406028 92268
rect 405974 90248 406030 90257
rect 405974 90183 405976 90192
rect 406028 90183 406030 90192
rect 405976 90154 406028 90160
rect 410220 87362 410248 88860
rect 410208 87356 410260 87362
rect 410208 87298 410260 87304
rect 412888 86721 412916 88860
rect 415556 87430 415584 88860
rect 418224 87498 418252 88860
rect 419788 88846 420906 88874
rect 422548 88846 423574 88874
rect 418212 87492 418264 87498
rect 418212 87434 418264 87440
rect 415544 87424 415596 87430
rect 415544 87366 415596 87372
rect 412874 86712 412930 86721
rect 412874 86647 412930 86656
rect 419788 47446 419816 88846
rect 419776 47440 419828 47446
rect 419776 47382 419828 47388
rect 422548 45406 422576 88846
rect 422536 45400 422588 45406
rect 422536 45342 422588 45348
rect 427332 15486 427360 126223
rect 427424 116466 427452 220199
rect 429712 215808 429764 215814
rect 429712 215750 429764 215756
rect 429724 215377 429752 215750
rect 429710 215368 429766 215377
rect 429710 215303 429766 215312
rect 428698 215232 428754 215241
rect 428698 215167 428754 215176
rect 427502 205304 427558 205313
rect 427502 205239 427558 205248
rect 427516 153730 427544 205239
rect 427594 195240 427650 195249
rect 427594 195175 427650 195184
rect 427608 178550 427636 195175
rect 427596 178544 427648 178550
rect 427596 178486 427648 178492
rect 427504 153724 427556 153730
rect 427504 153666 427556 153672
rect 428712 127793 428740 215167
rect 430078 202856 430134 202865
rect 430078 202791 430134 202800
rect 428792 199760 428844 199766
rect 428792 199702 428844 199708
rect 428804 165329 428832 199702
rect 430092 185486 430120 202791
rect 430080 185480 430132 185486
rect 430080 185422 430132 185428
rect 429896 178544 429948 178550
rect 429896 178486 429948 178492
rect 429908 177841 429936 178486
rect 429894 177832 429950 177841
rect 429894 177767 429950 177776
rect 428790 165320 428846 165329
rect 428790 165255 428846 165264
rect 429436 153724 429488 153730
rect 429436 153666 429488 153672
rect 429448 152817 429476 153666
rect 429434 152808 429490 152817
rect 429434 152743 429490 152752
rect 429528 140804 429580 140810
rect 429528 140746 429580 140752
rect 429540 140305 429568 140746
rect 429526 140296 429582 140305
rect 429526 140231 429582 140240
rect 428698 127784 428754 127793
rect 428698 127719 428754 127728
rect 427502 121256 427558 121265
rect 427502 121191 427558 121200
rect 427412 116460 427464 116466
rect 427412 116402 427464 116408
rect 427410 101264 427466 101273
rect 427410 101199 427466 101208
rect 427424 77842 427452 101199
rect 427412 77836 427464 77842
rect 427412 77778 427464 77784
rect 427516 28134 427544 121191
rect 429436 116460 429488 116466
rect 429436 116402 429488 116408
rect 428698 116224 428754 116233
rect 428698 116159 428754 116168
rect 427594 111328 427650 111337
rect 427594 111263 427650 111272
rect 427608 111026 427636 111263
rect 427596 111020 427648 111026
rect 427596 110962 427648 110968
rect 427594 106296 427650 106305
rect 427594 106231 427650 106240
rect 427608 105518 427636 106231
rect 427596 105512 427648 105518
rect 427596 105454 427648 105460
rect 427596 102724 427648 102730
rect 427596 102666 427648 102672
rect 427608 91617 427636 102666
rect 427594 91608 427650 91617
rect 427594 91543 427650 91552
rect 428056 81304 428108 81310
rect 428056 81246 428108 81252
rect 427504 28128 427556 28134
rect 427504 28070 427556 28076
rect 427320 15480 427372 15486
rect 427320 15422 427372 15428
rect 402756 12352 402808 12358
rect 402756 12294 402808 12300
rect 385184 12148 385236 12154
rect 385184 12090 385236 12096
rect 389876 12148 389928 12154
rect 389876 12090 389928 12096
rect 389888 9304 389916 12090
rect 402768 9304 402796 12294
rect 415636 12284 415688 12290
rect 415636 12226 415688 12232
rect 415648 9304 415676 12226
rect 428068 9434 428096 81246
rect 428712 40209 428740 116159
rect 429448 115281 429476 116402
rect 429434 115272 429490 115281
rect 429434 115207 429490 115216
rect 428792 111020 428844 111026
rect 428792 110962 428844 110968
rect 428804 52721 428832 110962
rect 430080 105512 430132 105518
rect 430080 105454 430132 105460
rect 429434 102760 429490 102769
rect 429434 102695 429436 102704
rect 429488 102695 429490 102704
rect 429436 102666 429488 102672
rect 429528 77836 429580 77842
rect 429528 77778 429580 77784
rect 429540 77745 429568 77778
rect 429526 77736 429582 77745
rect 429526 77671 429582 77680
rect 430092 65233 430120 105454
rect 430172 95856 430224 95862
rect 430172 95798 430224 95804
rect 430184 90257 430212 95798
rect 430170 90248 430226 90257
rect 430170 90183 430226 90192
rect 430078 65224 430134 65233
rect 430078 65159 430134 65168
rect 428790 52712 428846 52721
rect 428790 52647 428846 52656
rect 428698 40200 428754 40209
rect 428698 40135 428754 40144
rect 429804 28128 429856 28134
rect 429804 28070 429856 28076
rect 429816 27697 429844 28070
rect 429802 27688 429858 27697
rect 429802 27623 429858 27632
rect 429436 15480 429488 15486
rect 429436 15422 429488 15428
rect 429448 15185 429476 15422
rect 429434 15176 429490 15185
rect 429434 15111 429490 15120
rect 428056 9428 428108 9434
rect 428056 9370 428108 9376
rect 428516 9428 428568 9434
rect 428516 9370 428568 9376
rect 428528 9304 428556 9370
rect 16354 8824 16410 9304
rect 29234 8824 29290 9304
rect 42114 8824 42170 9304
rect 54994 8824 55050 9304
rect 67874 8824 67930 9304
rect 80754 8824 80810 9304
rect 93634 8824 93690 9304
rect 106514 8824 106570 9304
rect 119394 8824 119450 9304
rect 132274 8824 132330 9304
rect 145154 8824 145210 9304
rect 158034 8824 158090 9304
rect 170914 8824 170970 9304
rect 183794 8824 183850 9304
rect 196674 8824 196730 9304
rect 209554 8824 209610 9304
rect 222434 8824 222490 9304
rect 235314 8824 235370 9304
rect 248194 8824 248250 9304
rect 261074 8824 261130 9304
rect 273954 8824 274010 9304
rect 286834 8824 286890 9304
rect 299714 8824 299770 9304
rect 312594 8824 312650 9304
rect 325474 8824 325530 9304
rect 338354 8824 338410 9304
rect 351234 8824 351290 9304
rect 364114 8824 364170 9304
rect 376994 8824 377050 9304
rect 389874 8824 389930 9304
rect 402754 8824 402810 9304
rect 415634 8824 415690 9304
rect 428514 8824 428570 9304
<< via2 >>
rect 13318 390072 13374 390128
rect 12674 283040 12730 283096
rect 12858 269712 12914 269768
rect 13594 376744 13650 376800
rect 13502 363280 13558 363336
rect 13410 349952 13466 350008
rect 13410 336624 13466 336680
rect 76062 353896 76118 353952
rect 76430 353896 76486 353952
rect 13962 323160 14018 323216
rect 16078 313776 16134 313832
rect 13962 309832 14018 309888
rect 13686 296368 13742 296424
rect 12858 256248 12914 256304
rect 13134 242920 13190 242976
rect 13042 229612 13098 229648
rect 16170 308336 16226 308392
rect 16262 304120 16318 304176
rect 38802 315544 38858 315600
rect 38434 313096 38490 313152
rect 38802 310376 38858 310432
rect 16446 298680 16502 298736
rect 38802 308064 38858 308120
rect 38802 305616 38858 305672
rect 38618 303032 38674 303088
rect 38802 300620 38804 300640
rect 38804 300620 38856 300640
rect 38856 300620 38858 300640
rect 38802 300584 38858 300620
rect 38250 298136 38306 298192
rect 38802 295416 38858 295472
rect 17458 293784 17514 293840
rect 38434 293104 38490 293160
rect 38618 290520 38674 290576
rect 16722 289024 16778 289080
rect 38802 288072 38858 288128
rect 38802 285508 38858 285544
rect 38802 285488 38804 285508
rect 38804 285488 38856 285508
rect 38856 285488 38858 285508
rect 16538 283448 16594 283504
rect 38066 283040 38122 283096
rect 38066 280320 38122 280376
rect 51222 313796 51278 313832
rect 51222 313776 51224 313796
rect 51224 313776 51276 313796
rect 51276 313776 51278 313796
rect 51222 308608 51278 308664
rect 50302 300620 50304 300640
rect 50304 300620 50356 300640
rect 50356 300620 50358 300640
rect 50302 300584 50358 300620
rect 53062 327376 53118 327432
rect 54074 327376 54130 327432
rect 56098 327376 56154 327432
rect 54074 317856 54130 317912
rect 52694 315852 52696 315872
rect 52696 315852 52748 315872
rect 52748 315852 52750 315872
rect 52694 315816 52750 315852
rect 54074 310376 54130 310432
rect 73394 307112 73450 307168
rect 54442 306196 54444 306216
rect 54444 306196 54496 306216
rect 54496 306196 54498 306216
rect 54442 306160 54498 306196
rect 73394 305616 73450 305672
rect 51406 304140 51462 304176
rect 51406 304120 51408 304140
rect 51408 304120 51460 304140
rect 51460 304120 51462 304140
rect 51406 298816 51462 298872
rect 51314 293804 51370 293840
rect 51314 293784 51316 293804
rect 51316 293784 51368 293804
rect 51368 293784 51370 293804
rect 51314 289024 51370 289080
rect 74222 314456 74278 314512
rect 74130 311056 74186 311112
rect 74038 290112 74094 290168
rect 16722 279368 16778 279424
rect 38618 278144 38674 278200
rect 47082 271616 47138 271672
rect 46622 259104 46678 259160
rect 46530 255976 46586 256032
rect 51498 283720 51554 283776
rect 75510 303984 75566 304040
rect 75418 299904 75474 299960
rect 74222 296912 74278 296968
rect 51498 279368 51554 279424
rect 74038 278144 74094 278200
rect 55546 266584 55602 266640
rect 53522 265496 53578 265552
rect 54534 265496 54590 265552
rect 56558 265496 56614 265552
rect 75970 296912 76026 296968
rect 75878 292968 75934 293024
rect 74222 271616 74278 271672
rect 74222 271072 74278 271128
rect 73946 263476 74002 263512
rect 73946 263456 73948 263476
rect 73948 263456 74000 263476
rect 74000 263456 74002 263476
rect 49198 262676 49200 262696
rect 49200 262676 49252 262696
rect 49252 262676 49254 262696
rect 49198 262640 49254 262676
rect 47082 252848 47138 252904
rect 46438 249720 46494 249776
rect 47082 237344 47138 237400
rect 13042 229592 13044 229612
rect 13044 229592 13096 229612
rect 13096 229592 13098 229612
rect 16170 219936 16226 219992
rect 13318 216128 13374 216184
rect 16078 214496 16134 214552
rect 13962 202800 14018 202856
rect 13318 189372 13320 189392
rect 13320 189372 13372 189392
rect 13372 189372 13374 189392
rect 13318 189336 13374 189372
rect 13410 176008 13466 176064
rect 12858 162680 12914 162736
rect 12858 149216 12914 149272
rect 12858 135888 12914 135944
rect 16078 126096 16134 126152
rect 12674 122560 12730 122616
rect 13410 109096 13466 109152
rect 13134 95804 13136 95824
rect 13136 95804 13188 95824
rect 13188 95804 13190 95824
rect 13134 95768 13190 95804
rect 13502 82304 13558 82360
rect 13318 68976 13374 69032
rect 13134 55684 13136 55704
rect 13136 55684 13188 55704
rect 13188 55684 13190 55704
rect 13134 55648 13190 55684
rect 12858 42184 12914 42240
rect 12674 28856 12730 28912
rect 17550 209600 17606 209656
rect 16262 208920 16318 208976
rect 17550 208920 17606 208976
rect 38526 221704 38582 221760
rect 38066 219392 38122 219448
rect 38526 216808 38582 216864
rect 38526 214224 38582 214280
rect 16354 204840 16410 204896
rect 17642 199672 17698 199728
rect 17458 195320 17514 195376
rect 16446 189608 16502 189664
rect 17458 185428 17460 185448
rect 17460 185428 17512 185448
rect 17512 185428 17514 185448
rect 17458 185392 17514 185428
rect 38710 211504 38766 211560
rect 38526 209192 38582 209248
rect 38526 206608 38582 206664
rect 38526 204432 38582 204488
rect 38526 201440 38582 201496
rect 38526 199128 38582 199184
rect 38526 196408 38582 196464
rect 38802 194504 38858 194560
rect 38802 191512 38858 191568
rect 38066 189200 38122 189256
rect 38066 186480 38122 186536
rect 38802 184052 38858 184088
rect 38802 184032 38804 184052
rect 38804 184032 38856 184052
rect 38856 184032 38858 184052
rect 16170 120656 16226 120712
rect 16262 115080 16318 115136
rect 16354 111000 16410 111056
rect 18102 106240 18158 106296
rect 17458 101208 17514 101264
rect 18102 96176 18158 96232
rect 18102 91280 18158 91336
rect 45794 175872 45850 175928
rect 46898 176416 46954 176472
rect 46898 175872 46954 175928
rect 46898 165128 46954 165184
rect 46622 162000 46678 162056
rect 46530 158872 46586 158928
rect 46438 155744 46494 155800
rect 50578 222012 50580 222032
rect 50580 222012 50632 222032
rect 50632 222012 50634 222032
rect 50578 221976 50634 222012
rect 51222 200216 51278 200272
rect 51406 215176 51462 215232
rect 51406 210144 51462 210200
rect 51406 206780 51408 206800
rect 51408 206780 51460 206800
rect 51460 206780 51462 206800
rect 51406 206744 51462 206780
rect 51406 205248 51462 205304
rect 53522 232448 53578 232504
rect 54534 232448 54590 232504
rect 55546 232448 55602 232504
rect 55546 226872 55602 226928
rect 74130 233672 74186 233728
rect 74682 235032 74738 235088
rect 73946 224288 74002 224344
rect 73946 223880 74002 223936
rect 53246 221296 53302 221352
rect 52050 220208 52106 220264
rect 54074 210980 54130 211016
rect 54074 210960 54076 210980
rect 54076 210960 54128 210980
rect 54128 210960 54130 210980
rect 70818 209464 70874 209520
rect 73854 204976 73910 205032
rect 70818 204704 70874 204760
rect 73854 204704 73910 204760
rect 51314 195204 51370 195240
rect 51314 195184 51316 195204
rect 51316 195184 51368 195204
rect 51368 195184 51370 195204
rect 51222 190152 51278 190208
rect 51406 185256 51462 185312
rect 73946 185528 74002 185584
rect 73946 185392 74002 185448
rect 74222 220344 74278 220400
rect 74130 206472 74186 206528
rect 74130 204840 74186 204896
rect 74130 203480 74186 203536
rect 76062 235068 76064 235088
rect 76064 235068 76116 235088
rect 76116 235068 76118 235088
rect 76062 235032 76118 235068
rect 80202 357568 80258 357624
rect 80202 356344 80258 356400
rect 80202 354984 80258 355040
rect 79282 354576 79338 354632
rect 78914 353352 78970 353408
rect 80202 352128 80258 352184
rect 87194 351312 87250 351368
rect 80202 350632 80258 350688
rect 79098 350360 79154 350416
rect 97498 367224 97554 367280
rect 97314 352012 97370 352048
rect 97314 351992 97316 352012
rect 97316 351992 97368 352012
rect 97368 351992 97370 352012
rect 131354 384768 131410 384824
rect 225194 384768 225250 384824
rect 87470 350360 87526 350416
rect 87286 349544 87342 349600
rect 80202 349272 80258 349328
rect 80202 348048 80258 348104
rect 87102 347776 87158 347832
rect 80202 346688 80258 346744
rect 79282 346280 79338 346336
rect 80202 344804 80258 344840
rect 87378 348592 87434 348648
rect 87194 346824 87250 346880
rect 88114 346008 88170 346064
rect 87378 345056 87434 345112
rect 80202 344784 80204 344804
rect 80204 344784 80256 344804
rect 80256 344784 80258 344804
rect 79650 343968 79706 344024
rect 80202 342764 80258 342800
rect 80202 342744 80204 342764
rect 80204 342744 80256 342764
rect 80256 342744 80258 342764
rect 87286 343288 87342 343344
rect 80202 341792 80258 341848
rect 87194 341520 87250 341576
rect 80202 340976 80258 341032
rect 80202 339752 80258 339808
rect 80202 338392 80258 338448
rect 80110 337984 80166 338040
rect 79834 336760 79890 336816
rect 80202 335672 80258 335728
rect 80110 334040 80166 334096
rect 88482 344240 88538 344296
rect 87562 342336 87618 342392
rect 87378 340568 87434 340624
rect 87286 339752 87342 339808
rect 87194 337984 87250 338040
rect 87194 336216 87250 336272
rect 80202 333632 80258 333688
rect 80202 332680 80258 332736
rect 80202 330912 80258 330968
rect 87470 338800 87526 338856
rect 87562 337032 87618 337088
rect 82318 329688 82374 329744
rect 95198 333768 95254 333824
rect 131446 382048 131502 382104
rect 131538 380144 131594 380200
rect 131630 377424 131686 377480
rect 131722 374704 131778 374760
rect 131814 372120 131870 372176
rect 131814 351312 131870 351368
rect 131814 350360 131870 350416
rect 131906 349544 131962 349600
rect 131814 348592 131870 348648
rect 132182 347776 132238 347832
rect 131906 346824 131962 346880
rect 131814 346008 131870 346064
rect 132366 345056 132422 345112
rect 131814 344260 131870 344296
rect 131814 344240 131816 344260
rect 131816 344240 131868 344260
rect 131868 344240 131870 344260
rect 131814 343288 131870 343344
rect 131906 342336 131962 342392
rect 131814 341520 131870 341576
rect 131814 340568 131870 340624
rect 131906 339752 131962 339808
rect 131814 338800 131870 338856
rect 131814 337984 131870 338040
rect 131906 337032 131962 337088
rect 131814 336216 131870 336272
rect 81674 313540 81676 313560
rect 81676 313540 81728 313560
rect 81728 313540 81730 313560
rect 81674 313504 81730 313540
rect 76890 305616 76946 305672
rect 81674 296776 81730 296832
rect 81674 280184 81730 280240
rect 78914 263592 78970 263648
rect 78914 261688 78970 261744
rect 78914 260328 78970 260384
rect 78914 258832 78970 258888
rect 78914 257472 78970 257528
rect 78914 256112 78970 256168
rect 78914 254616 78970 254672
rect 87194 258016 87250 258072
rect 131354 257336 131410 257392
rect 87194 256828 87196 256848
rect 87196 256828 87248 256848
rect 87248 256828 87250 256848
rect 87194 256792 87250 256828
rect 87286 255568 87342 255624
rect 87194 255296 87250 255352
rect 131354 254636 131410 254672
rect 131354 254616 131356 254636
rect 131356 254616 131408 254636
rect 131408 254616 131410 254636
rect 78914 253256 78970 253312
rect 87194 254380 87196 254400
rect 87196 254380 87248 254400
rect 87248 254380 87250 254400
rect 87194 254344 87250 254380
rect 131354 253800 131410 253856
rect 87194 252884 87196 252904
rect 87196 252884 87248 252904
rect 87248 252884 87250 252904
rect 87194 252848 87250 252884
rect 131354 252848 131410 252904
rect 87286 252712 87342 252768
rect 78914 251896 78970 251952
rect 87194 251488 87250 251544
rect 79742 250536 79798 250592
rect 87194 250300 87196 250320
rect 87196 250300 87248 250320
rect 87248 250300 87250 250320
rect 87194 250264 87250 250300
rect 131998 255568 132054 255624
rect 131998 250264 132054 250320
rect 131814 249992 131870 250048
rect 78914 249312 78970 249368
rect 87194 249312 87250 249368
rect 132366 256384 132422 256440
rect 132182 251080 132238 251136
rect 132090 248904 132146 248960
rect 87194 248360 87250 248416
rect 78914 247952 78970 248008
rect 88482 247564 88538 247600
rect 88482 247544 88484 247564
rect 88484 247544 88536 247564
rect 88536 247544 88538 247564
rect 78914 246864 78970 246920
rect 87194 246592 87250 246648
rect 87194 245776 87250 245832
rect 78914 245504 78970 245560
rect 87102 244824 87158 244880
rect 78914 244144 78970 244200
rect 87010 244008 87066 244064
rect 78914 242512 78970 242568
rect 78914 240608 78970 240664
rect 79006 239248 79062 239304
rect 131354 245504 131410 245560
rect 87286 243056 87342 243112
rect 87194 242240 87250 242296
rect 98924 241696 98980 241752
rect 95198 239656 95254 239712
rect 91702 239384 91758 239440
rect 79098 238568 79154 238624
rect 102466 237888 102522 237944
rect 78914 236564 78916 236584
rect 78916 236564 78968 236584
rect 78968 236564 78970 236584
rect 78914 236528 78970 236564
rect 106146 235712 106202 235768
rect 117094 235848 117150 235904
rect 132458 248224 132514 248280
rect 132366 247000 132422 247056
rect 132274 246048 132330 246104
rect 133378 252032 133434 252088
rect 132550 244688 132606 244744
rect 132550 243056 132606 243112
rect 132642 242784 132698 242840
rect 139634 357704 139690 357760
rect 174042 357160 174098 357216
rect 139634 356516 139636 356536
rect 139636 356516 139688 356536
rect 139688 356516 139690 356536
rect 139634 356480 139690 356516
rect 173490 356072 173546 356128
rect 139634 355156 139636 355176
rect 139636 355156 139688 355176
rect 139688 355156 139690 355176
rect 139634 355120 139690 355156
rect 174042 355156 174044 355176
rect 174044 355156 174096 355176
rect 174096 355156 174098 355176
rect 174042 355120 174098 355156
rect 139726 354576 139782 354632
rect 173766 354032 173822 354088
rect 139634 353488 139690 353544
rect 174042 352944 174098 353000
rect 139634 352264 139690 352320
rect 174042 351992 174098 352048
rect 180850 351584 180906 351640
rect 139726 350904 139782 350960
rect 139634 350496 139690 350552
rect 174042 350940 174044 350960
rect 174044 350940 174096 350960
rect 174096 350940 174098 350960
rect 174042 350904 174098 350940
rect 173766 349816 173822 349872
rect 139634 349544 139690 349600
rect 180942 349952 180998 350008
rect 173030 348864 173086 348920
rect 139634 348220 139636 348240
rect 139636 348220 139688 348240
rect 139688 348220 139690 348240
rect 139634 348184 139690 348220
rect 182322 349544 182378 349600
rect 182138 348592 182194 348648
rect 172938 347776 172994 347832
rect 180942 347232 180998 347288
rect 139634 346860 139636 346880
rect 139636 346860 139688 346880
rect 139688 346860 139690 346880
rect 139634 346824 139690 346860
rect 139726 346280 139782 346336
rect 174042 346860 174044 346880
rect 174044 346860 174096 346880
rect 174096 346860 174098 346880
rect 174042 346824 174098 346860
rect 173766 345736 173822 345792
rect 139818 345328 139874 345384
rect 172754 344648 172810 344704
rect 139634 344104 139690 344160
rect 139634 342608 139690 342664
rect 139726 342200 139782 342256
rect 172846 343696 172902 343752
rect 181586 346824 181642 346880
rect 182322 346008 182378 346064
rect 180942 344648 180998 344704
rect 172938 342608 172994 342664
rect 172754 341520 172810 341576
rect 139818 341248 139874 341304
rect 173122 340568 173178 340624
rect 139634 339888 139690 339944
rect 139542 336760 139598 336816
rect 136874 332136 136930 332192
rect 137058 331456 137114 331512
rect 136874 307792 136930 307848
rect 139726 338564 139728 338584
rect 139728 338564 139780 338584
rect 139780 338564 139782 338584
rect 139726 338528 139782 338564
rect 139818 337984 139874 338040
rect 139634 335808 139690 335864
rect 139634 334312 139690 334368
rect 139634 333904 139690 333960
rect 137058 314048 137114 314104
rect 137518 310920 137574 310976
rect 136966 304120 137022 304176
rect 137518 304120 137574 304176
rect 136874 301536 136930 301592
rect 136874 284808 136930 284864
rect 136874 279368 136930 279424
rect 139634 332952 139690 333008
rect 172846 332272 172902 332328
rect 139818 331592 139874 331648
rect 173766 337440 173822 337496
rect 173490 335400 173546 335456
rect 182322 344240 182378 344296
rect 181402 343288 181458 343344
rect 181402 342336 181458 342392
rect 182322 341540 182378 341576
rect 182322 341520 182324 341540
rect 182324 341520 182376 341540
rect 182376 341520 182378 341540
rect 173950 339480 174006 339536
rect 181402 340568 181458 340624
rect 181586 339752 181642 339808
rect 180298 339344 180354 339400
rect 174042 338528 174098 338584
rect 173858 336352 173914 336408
rect 181770 337984 181826 338040
rect 181586 337032 181642 337088
rect 181770 336216 181826 336272
rect 174042 334348 174044 334368
rect 174044 334348 174096 334368
rect 174096 334348 174098 334368
rect 174042 334312 174098 334348
rect 173674 333224 173730 333280
rect 172938 331184 172994 331240
rect 140554 330232 140610 330288
rect 173398 330232 173454 330288
rect 159598 330096 159654 330152
rect 137702 317176 137758 317232
rect 137610 298544 137666 298600
rect 137610 285216 137666 285272
rect 137518 273792 137574 273848
rect 136874 235848 136930 235904
rect 137058 235712 137114 235768
rect 136874 235032 136930 235088
rect 75418 217352 75474 217408
rect 74682 210144 74738 210200
rect 74406 204840 74462 204896
rect 74406 204704 74462 204760
rect 74222 195184 74278 195240
rect 74498 195184 74554 195240
rect 74222 195048 74278 195104
rect 74498 195048 74554 195104
rect 74130 187976 74186 188032
rect 74314 185664 74370 185720
rect 74222 185528 74278 185584
rect 74038 184984 74094 185040
rect 53522 172880 53578 172936
rect 54534 172880 54590 172936
rect 55546 172880 55602 172936
rect 56558 172744 56614 172800
rect 74314 173696 74370 173752
rect 71646 169480 71702 169536
rect 49198 168836 49200 168856
rect 49200 168836 49252 168856
rect 49252 168836 49254 168856
rect 49198 168800 49254 168836
rect 47082 143368 47138 143424
rect 73946 142144 74002 142200
rect 75418 142144 75474 142200
rect 38802 127456 38858 127512
rect 48462 127184 48518 127240
rect 38250 125552 38306 125608
rect 38802 122696 38858 122752
rect 38802 120248 38858 120304
rect 38250 117528 38306 117584
rect 38802 114944 38858 115000
rect 38802 112768 38858 112824
rect 38250 110456 38306 110512
rect 38802 107484 38858 107520
rect 38802 107464 38804 107484
rect 38804 107464 38856 107484
rect 38856 107464 38858 107484
rect 38802 105288 38858 105344
rect 38618 102432 38674 102488
rect 38802 100256 38858 100312
rect 38802 97828 38858 97864
rect 38802 97808 38804 97828
rect 38804 97808 38856 97828
rect 38856 97808 38858 97828
rect 38066 95360 38122 95416
rect 37606 92504 37662 92560
rect 53522 139560 53578 139616
rect 54534 139560 54590 139616
rect 55546 134392 55602 134448
rect 56098 132352 56154 132408
rect 52602 126232 52658 126288
rect 54074 122016 54130 122072
rect 52602 121200 52658 121256
rect 73394 120520 73450 120576
rect 73394 119704 73450 119760
rect 54074 117140 54130 117176
rect 54074 117120 54076 117140
rect 54076 117120 54128 117140
rect 54128 117120 54130 117140
rect 52142 116168 52198 116224
rect 51866 113040 51922 113096
rect 52602 111272 52658 111328
rect 52602 106240 52658 106296
rect 38802 90056 38858 90112
rect 52602 101208 52658 101264
rect 52602 96176 52658 96232
rect 73486 115080 73542 115136
rect 52602 91280 52658 91336
rect 73394 91144 73450 91200
rect 54074 77952 54130 78008
rect 53062 77816 53118 77872
rect 55086 77816 55142 77872
rect 56098 77816 56154 77872
rect 72014 87492 72070 87528
rect 72014 87472 72016 87492
rect 72016 87472 72068 87492
rect 72068 87472 72070 87492
rect 73578 112768 73634 112824
rect 73670 109504 73726 109560
rect 73670 108824 73726 108880
rect 76062 142044 76064 142064
rect 76064 142044 76116 142064
rect 76116 142044 76118 142064
rect 76062 142008 76118 142044
rect 74222 139424 74278 139480
rect 75142 139424 75198 139480
rect 76062 137112 76118 137168
rect 74314 126368 74370 126424
rect 74222 120520 74278 120576
rect 74130 116168 74186 116224
rect 74130 115080 74186 115136
rect 75418 122696 75474 122752
rect 74038 105152 74094 105208
rect 81674 219548 81730 219584
rect 81674 219528 81676 219548
rect 81676 219528 81728 219548
rect 81728 219528 81730 219548
rect 81674 202800 81730 202856
rect 81674 186208 81730 186264
rect 79742 169072 79798 169128
rect 77258 167644 77314 167700
rect 77258 166284 77314 166340
rect 79742 164876 79798 164912
rect 79742 164856 79744 164876
rect 79744 164856 79796 164876
rect 79796 164856 79798 164876
rect 77258 163428 77314 163484
rect 77166 162068 77222 162124
rect 87194 164040 87250 164096
rect 87194 163088 87250 163144
rect 87286 161900 87288 161920
rect 87288 161900 87340 161920
rect 87340 161900 87342 161920
rect 87286 161864 87342 161900
rect 87194 161320 87250 161376
rect 87194 160368 87250 160424
rect 81674 159960 81730 160016
rect 79282 159300 79338 159336
rect 79282 159280 79284 159300
rect 79284 159280 79336 159300
rect 79336 159280 79338 159300
rect 87194 158872 87250 158928
rect 87286 158600 87342 158656
rect 79742 157940 79798 157976
rect 79742 157920 79744 157940
rect 79744 157920 79796 157940
rect 79796 157920 79798 157940
rect 87194 157784 87250 157840
rect 77258 156512 77314 156548
rect 77258 156492 77260 156512
rect 77260 156492 77312 156512
rect 77312 156492 77314 156512
rect 87194 156288 87250 156344
rect 87194 155336 87250 155392
rect 79742 155084 79798 155120
rect 79742 155064 79744 155084
rect 79744 155064 79796 155084
rect 79796 155064 79798 155084
rect 87194 154404 87250 154440
rect 87194 154384 87196 154404
rect 87196 154384 87248 154404
rect 87248 154384 87250 154404
rect 79742 153704 79798 153760
rect 87194 153568 87250 153624
rect 87194 152616 87250 152672
rect 79742 152344 79798 152400
rect 77258 150780 77314 150836
rect 87470 151800 87526 151856
rect 78914 148944 78970 149000
rect 76982 148536 77038 148592
rect 76890 145816 76946 145872
rect 78914 147856 78970 147912
rect 87010 150848 87066 150904
rect 87194 150032 87250 150088
rect 87194 149080 87250 149136
rect 87102 148264 87158 148320
rect 80110 146632 80166 146688
rect 79374 145272 79430 145328
rect 76982 144048 77038 144104
rect 78914 143504 78970 143560
rect 88574 142824 88630 142880
rect 78914 141872 78970 141928
rect 98878 144184 98934 144240
rect 95290 144048 95346 144104
rect 109734 143232 109790 143288
rect 106146 141872 106202 141928
rect 131354 163396 131356 163416
rect 131356 163396 131408 163416
rect 131408 163396 131410 163416
rect 131354 163360 131410 163396
rect 131998 162408 132054 162464
rect 131538 161592 131594 161648
rect 131354 160676 131356 160696
rect 131356 160676 131408 160696
rect 131408 160676 131410 160696
rect 131354 160640 131410 160676
rect 131354 158872 131410 158928
rect 131354 149080 131410 149136
rect 131814 159824 131870 159880
rect 131722 150440 131778 150496
rect 131998 155064 132054 155120
rect 132274 158056 132330 158112
rect 132182 156016 132238 156072
rect 132090 153568 132146 153624
rect 131906 150848 131962 150904
rect 131630 148808 131686 148864
rect 132458 157104 132514 157160
rect 132366 156288 132422 156344
rect 132550 153296 132606 153352
rect 132642 152208 132698 152264
rect 84710 127476 84766 127512
rect 84710 127456 84712 127476
rect 84712 127456 84764 127476
rect 84764 127456 84766 127476
rect 82686 125452 82688 125472
rect 82688 125452 82740 125472
rect 82740 125452 82742 125472
rect 82686 125416 82742 125452
rect 74038 89784 74094 89840
rect 73578 86248 73634 86304
rect 73854 86384 73910 86440
rect 73486 86112 73542 86168
rect 73670 86112 73726 86168
rect 84710 109796 84766 109832
rect 84710 109776 84712 109796
rect 84712 109776 84764 109796
rect 84764 109776 84766 109796
rect 82594 108824 82650 108880
rect 84802 93476 84858 93512
rect 84802 93456 84804 93476
rect 84804 93456 84856 93476
rect 84856 93456 84858 93476
rect 82686 92232 82742 92288
rect 79466 75776 79522 75832
rect 80202 73872 80258 73928
rect 79834 72784 79890 72840
rect 78914 71560 78970 71616
rect 80202 71152 80258 71208
rect 80202 69792 80258 69848
rect 79282 68568 79338 68624
rect 79466 64508 79522 64544
rect 79466 64488 79468 64508
rect 79468 64488 79520 64508
rect 79520 64488 79522 64508
rect 78914 56056 78970 56112
rect 80202 67344 80258 67400
rect 80202 66820 80258 66856
rect 80202 66800 80204 66820
rect 80204 66800 80256 66820
rect 80256 66800 80258 66820
rect 80202 65576 80258 65632
rect 87194 66700 87196 66720
rect 87196 66700 87248 66720
rect 87248 66700 87250 66720
rect 87194 66664 87250 66700
rect 87930 69384 87986 69440
rect 87654 68432 87710 68488
rect 87838 67616 87894 67672
rect 87286 65848 87342 65904
rect 80202 63264 80258 63320
rect 80202 62856 80258 62912
rect 87194 64080 87250 64136
rect 80202 61380 80258 61416
rect 80202 61360 80204 61380
rect 80204 61360 80256 61380
rect 80256 61360 80258 61380
rect 80202 60156 80258 60192
rect 80202 60136 80204 60156
rect 80204 60136 80256 60156
rect 80256 60136 80258 60156
rect 79650 59048 79706 59104
rect 80202 58540 80204 58560
rect 80204 58540 80256 58560
rect 80256 58540 80258 58560
rect 80202 58504 80258 58540
rect 131354 69384 131410 69440
rect 131814 68432 131870 68488
rect 132366 67616 132422 67672
rect 87470 64896 87526 64952
rect 87378 63128 87434 63184
rect 87286 62312 87342 62368
rect 87194 61360 87250 61416
rect 87194 60408 87250 60464
rect 87838 59592 87894 59648
rect 87194 58640 87250 58696
rect 80202 57164 80258 57200
rect 80202 57144 80204 57164
rect 80204 57144 80256 57164
rect 80256 57144 80258 57164
rect 87194 57824 87250 57880
rect 87194 56872 87250 56928
rect 87286 56056 87342 56112
rect 79558 55648 79614 55704
rect 80202 54560 80258 54616
rect 87194 55104 87250 55160
rect 87194 54308 87250 54344
rect 87194 54288 87196 54308
rect 87196 54288 87248 54308
rect 87248 54288 87250 54308
rect 80202 53644 80204 53664
rect 80204 53644 80256 53664
rect 80256 53644 80258 53664
rect 80202 53608 80258 53644
rect 80202 52656 80258 52712
rect 132550 66664 132606 66720
rect 132366 65848 132422 65904
rect 131354 64896 131410 64952
rect 132182 64080 132238 64136
rect 132366 63128 132422 63184
rect 131354 62312 131410 62368
rect 131722 61360 131778 61416
rect 131354 60408 131410 60464
rect 131354 59592 131410 59648
rect 131446 58640 131502 58696
rect 131354 57824 131410 57880
rect 131354 56872 131410 56928
rect 132182 56056 132238 56112
rect 131354 55104 131410 55160
rect 78914 50752 78970 50808
rect 80202 50244 80204 50264
rect 80204 50244 80256 50264
rect 80256 50244 80258 50264
rect 80202 50208 80258 50244
rect 88390 49256 88446 49312
rect 80202 49120 80258 49176
rect 88298 48576 88354 48632
rect 67874 48032 67930 48088
rect 74314 48032 74370 48088
rect 71462 47352 71518 47408
rect 73118 47352 73174 47408
rect 80202 48032 80258 48088
rect 88298 48032 88354 48088
rect 74222 46148 74278 46184
rect 74222 46128 74224 46148
rect 74224 46128 74276 46148
rect 74276 46128 74278 46148
rect 64194 45856 64250 45912
rect 88114 33616 88170 33672
rect 88206 30760 88262 30816
rect 88298 28040 88354 28096
rect 93634 50616 93690 50672
rect 102374 51296 102430 51352
rect 105134 49256 105190 49312
rect 105134 48032 105190 48088
rect 107526 50208 107582 50264
rect 106606 47352 106662 47408
rect 109458 50208 109514 50264
rect 109458 47216 109514 47272
rect 113966 53064 114022 53120
rect 118658 53064 118714 53120
rect 113598 43272 113654 43328
rect 118658 46128 118714 46184
rect 131354 54324 131356 54344
rect 131356 54324 131408 54344
rect 131408 54324 131410 54344
rect 131354 54288 131410 54324
rect 136966 234896 137022 234952
rect 136874 213816 136930 213872
rect 137334 234216 137390 234272
rect 137242 226328 137298 226384
rect 137886 320304 137942 320360
rect 137794 301536 137850 301592
rect 137702 279640 137758 279696
rect 137794 276512 137850 276568
rect 153250 326288 153306 326344
rect 161714 329416 161770 329472
rect 158126 327376 158182 327432
rect 198790 332136 198846 332192
rect 205598 331592 205654 331648
rect 226482 382764 226484 382784
rect 226484 382764 226536 382784
rect 226536 382764 226538 382784
rect 226482 382728 226538 382764
rect 225286 380144 225342 380200
rect 212314 333496 212370 333552
rect 225378 377424 225434 377480
rect 226482 374704 226538 374760
rect 225838 372120 225894 372176
rect 226298 351332 226354 351368
rect 226298 351312 226300 351332
rect 226300 351312 226352 351332
rect 226352 351312 226354 351332
rect 226390 350360 226446 350416
rect 226482 349544 226538 349600
rect 226390 348592 226446 348648
rect 226390 347776 226446 347832
rect 226298 346824 226354 346880
rect 226390 346008 226446 346064
rect 226482 345056 226538 345112
rect 226390 344240 226446 344296
rect 226390 343288 226446 343344
rect 226482 342336 226538 342392
rect 226390 341520 226446 341576
rect 226390 340568 226446 340624
rect 226482 339752 226538 339808
rect 226390 338800 226446 338856
rect 226390 337984 226446 338040
rect 226390 337032 226446 337088
rect 226574 336216 226630 336272
rect 225286 331592 225342 331648
rect 165118 315816 165174 315872
rect 175514 313504 175570 313560
rect 145522 310104 145578 310160
rect 145430 296776 145486 296832
rect 145154 283484 145156 283504
rect 145156 283484 145208 283504
rect 145208 283484 145210 283504
rect 145154 283448 145210 283484
rect 138162 282496 138218 282552
rect 138438 279232 138494 279288
rect 137886 273384 137942 273440
rect 138438 269848 138494 269904
rect 157758 274744 157814 274800
rect 157206 274472 157262 274528
rect 156562 274336 156618 274392
rect 154722 273792 154778 273848
rect 159046 274880 159102 274936
rect 158402 274608 158458 274664
rect 167878 306160 167934 306216
rect 175514 296776 175570 296832
rect 168062 286304 168118 286360
rect 175422 280184 175478 280240
rect 182966 269440 183022 269496
rect 139818 263048 139874 263104
rect 138806 259920 138862 259976
rect 138806 250536 138862 250592
rect 138438 245504 138494 245560
rect 138438 240880 138494 240936
rect 139818 253256 139874 253312
rect 139726 248360 139782 248416
rect 140094 244008 140150 244064
rect 138990 242784 139046 242840
rect 138898 238568 138954 238624
rect 140370 261688 140426 261744
rect 140370 260328 140426 260384
rect 140554 258832 140610 258888
rect 140554 257472 140610 257528
rect 140462 256112 140518 256168
rect 140554 254616 140610 254672
rect 140554 251896 140610 251952
rect 140738 250536 140794 250592
rect 140646 249720 140702 249776
rect 140646 246728 140702 246784
rect 140370 245504 140426 245560
rect 140278 237208 140334 237264
rect 140554 240628 140610 240664
rect 140554 240608 140556 240628
rect 140556 240608 140608 240628
rect 140608 240608 140610 240628
rect 140554 239268 140610 239304
rect 140554 239248 140556 239268
rect 140556 239248 140608 239268
rect 140608 239248 140610 239268
rect 148742 235984 148798 236040
rect 137334 223200 137390 223256
rect 137150 220072 137206 220128
rect 137058 216944 137114 217000
rect 136966 210688 137022 210744
rect 136874 204740 136876 204760
rect 136876 204740 136928 204760
rect 136928 204740 136930 204760
rect 136874 204704 136930 204740
rect 137334 185664 137390 185720
rect 137150 143232 137206 143288
rect 136874 141872 136930 141928
rect 136874 132896 136930 132952
rect 137334 141056 137390 141112
rect 137242 140240 137298 140296
rect 137242 129768 137298 129824
rect 137058 125960 137114 126016
rect 136966 123240 137022 123296
rect 136874 120384 136930 120440
rect 136874 113176 136930 113232
rect 136874 110728 136930 110784
rect 137610 191920 137666 191976
rect 138162 208240 138218 208296
rect 137794 188520 137850 188576
rect 145154 235324 145210 235360
rect 145154 235304 145156 235324
rect 145156 235304 145208 235324
rect 145208 235304 145210 235324
rect 145154 216128 145210 216184
rect 147270 235848 147326 235904
rect 167970 235984 168026 236040
rect 148190 234896 148246 234952
rect 152008 235576 152064 235632
rect 150674 233672 150730 233728
rect 167694 235712 167750 235768
rect 164382 226600 164438 226656
rect 164382 226192 164438 226248
rect 145154 202800 145210 202856
rect 145614 189472 145670 189528
rect 137610 182536 137666 182592
rect 138898 179408 138954 179464
rect 154722 181992 154778 182048
rect 155274 181176 155330 181232
rect 157206 180768 157262 180824
rect 157758 180632 157814 180688
rect 155918 180496 155974 180552
rect 156562 180496 156618 180552
rect 159046 181040 159102 181096
rect 158402 180904 158458 180960
rect 167878 212728 167934 212784
rect 167970 192736 168026 192792
rect 173490 263048 173546 263104
rect 173398 261688 173454 261744
rect 173306 256112 173362 256168
rect 173306 254616 173362 254672
rect 173306 249040 173362 249096
rect 173766 260328 173822 260384
rect 173674 257472 173730 257528
rect 173582 250536 173638 250592
rect 173490 247680 173546 247736
rect 173306 246320 173362 246376
rect 172754 244824 172810 244880
rect 173122 243464 173178 243520
rect 218018 268352 218074 268408
rect 173858 258832 173914 258888
rect 181034 257336 181090 257392
rect 181034 256384 181090 256440
rect 173950 253256 174006 253312
rect 174042 251916 174098 251952
rect 174042 251896 174044 251916
rect 174044 251896 174096 251916
rect 174096 251896 174098 251916
rect 181586 255568 181642 255624
rect 181034 254616 181090 254672
rect 181034 253800 181090 253856
rect 225930 255568 225986 255624
rect 225746 253800 225802 253856
rect 181586 252848 181642 252904
rect 181678 252032 181734 252088
rect 181494 249720 181550 249776
rect 181586 245368 181642 245424
rect 182322 251080 182378 251136
rect 181770 250264 181826 250320
rect 181954 248632 182010 248688
rect 181862 248224 181918 248280
rect 182322 247136 182378 247192
rect 182322 245776 182378 245832
rect 182322 244552 182378 244608
rect 225838 250264 225894 250320
rect 225746 249312 225802 249368
rect 226022 251080 226078 251136
rect 225930 248360 225986 248416
rect 225562 244824 225618 244880
rect 225562 244008 225618 244064
rect 181034 243364 181036 243384
rect 181036 243364 181088 243384
rect 181088 243364 181090 243384
rect 181034 243328 181090 243364
rect 181218 242784 181274 242840
rect 174042 242104 174098 242160
rect 173582 240628 173638 240664
rect 173582 240608 173584 240628
rect 173584 240608 173636 240628
rect 173636 240608 173638 240628
rect 173306 239248 173362 239304
rect 189222 239656 189278 239712
rect 196490 240336 196546 240392
rect 192902 239384 192958 239440
rect 173398 237888 173454 237944
rect 172938 236528 172994 236584
rect 200170 238432 200226 238488
rect 203114 236256 203170 236312
rect 210014 234488 210070 234544
rect 207254 234352 207310 234408
rect 225746 242240 225802 242296
rect 222434 240608 222490 240664
rect 222802 240608 222858 240664
rect 219766 237752 219822 237808
rect 226206 247544 226262 247600
rect 226482 257356 226538 257392
rect 226482 257336 226484 257356
rect 226484 257336 226536 257356
rect 226536 257336 226538 257356
rect 226482 256384 226538 256440
rect 226390 254616 226446 254672
rect 226298 246592 226354 246648
rect 226482 252848 226538 252904
rect 226114 245776 226170 245832
rect 227218 252032 227274 252088
rect 226482 243092 226484 243112
rect 226484 243092 226536 243112
rect 226536 243092 226538 243112
rect 226482 243056 226538 243092
rect 139634 164856 139690 164912
rect 139634 163516 139690 163552
rect 139634 163496 139636 163516
rect 139636 163496 139688 163516
rect 139688 163496 139690 163516
rect 139634 162136 139690 162192
rect 139634 160660 139690 160696
rect 139634 160640 139636 160660
rect 139636 160640 139688 160660
rect 139688 160640 139690 160660
rect 139634 159300 139690 159336
rect 139634 159280 139636 159300
rect 139636 159280 139688 159300
rect 139688 159280 139690 159300
rect 139634 157940 139690 157976
rect 139634 157920 139636 157940
rect 139636 157920 139688 157940
rect 139688 157920 139690 157940
rect 139726 153704 139782 153760
rect 139634 152344 139690 152400
rect 139634 149524 139636 149544
rect 139636 149524 139688 149544
rect 139688 149524 139690 149544
rect 139634 149488 139690 149524
rect 138898 148128 138954 148184
rect 140554 169072 140610 169128
rect 140554 167712 140610 167768
rect 140554 166352 140610 166408
rect 140370 156560 140426 156616
rect 140278 142552 140334 142608
rect 140554 155064 140610 155120
rect 140462 150848 140518 150904
rect 140554 146632 140610 146688
rect 140554 145272 140610 145328
rect 140554 143912 140610 143968
rect 147914 142144 147970 142200
rect 150674 142144 150730 142200
rect 167970 142180 167972 142200
rect 167972 142180 168024 142200
rect 168024 142180 168026 142200
rect 167970 142144 168026 142180
rect 146810 142008 146866 142064
rect 137518 98488 137574 98544
rect 137610 92232 137666 92288
rect 138162 94544 138218 94600
rect 144234 122288 144290 122344
rect 149110 141056 149166 141112
rect 152054 140376 152110 140432
rect 147454 139832 147510 139888
rect 148190 139832 148246 139888
rect 152698 139832 152754 139888
rect 168522 141736 168578 141792
rect 167878 118752 167934 118808
rect 146626 113176 146682 113232
rect 143958 108824 144014 108880
rect 164934 99984 164990 100040
rect 167878 98760 167934 98816
rect 164934 98624 164990 98680
rect 137702 88696 137758 88752
rect 137886 85704 137942 85760
rect 145798 90056 145854 90112
rect 155458 88832 155514 88888
rect 155734 88832 155790 88888
rect 156102 87472 156158 87528
rect 155274 87336 155330 87392
rect 156562 86792 156618 86848
rect 157758 87200 157814 87256
rect 157206 86656 157262 86712
rect 159046 87064 159102 87120
rect 158402 86928 158458 86984
rect 178918 219528 178974 219584
rect 178918 202800 178974 202856
rect 178918 186208 178974 186264
rect 178274 178184 178330 178240
rect 182138 178184 182194 178240
rect 182874 175772 182876 175792
rect 182876 175772 182928 175792
rect 182928 175772 182930 175792
rect 182874 175736 182930 175772
rect 173582 169072 173638 169128
rect 173398 167712 173454 167768
rect 173306 164856 173362 164912
rect 172846 156560 172902 156616
rect 172938 153704 172994 153760
rect 173490 166352 173546 166408
rect 174042 163496 174098 163552
rect 173674 162136 173730 162192
rect 173214 152344 173270 152400
rect 173950 160660 174006 160696
rect 173950 160640 173952 160660
rect 173952 160640 174004 160660
rect 174004 160640 174006 160660
rect 173950 159316 173952 159336
rect 173952 159316 174004 159336
rect 174004 159316 174006 159336
rect 173950 159280 174006 159316
rect 173766 157940 173822 157976
rect 173766 157920 173768 157940
rect 173768 157920 173820 157940
rect 173820 157920 173822 157940
rect 173858 146632 173914 146688
rect 173766 145272 173822 145328
rect 174042 155084 174098 155120
rect 174042 155064 174044 155084
rect 174044 155064 174096 155084
rect 174096 155064 174098 155084
rect 174042 150848 174098 150904
rect 174042 149508 174098 149544
rect 174042 149488 174044 149508
rect 174044 149488 174096 149508
rect 174096 149488 174098 149508
rect 174042 148164 174044 148184
rect 174044 148164 174096 148184
rect 174096 148164 174098 148184
rect 174042 148128 174098 148164
rect 173950 143912 174006 143968
rect 173582 142552 173638 142608
rect 175514 125436 175570 125472
rect 175514 125416 175516 125436
rect 175516 125416 175568 125436
rect 175568 125416 175570 125436
rect 175514 92232 175570 92288
rect 218018 175464 218074 175520
rect 182322 163396 182324 163416
rect 182324 163396 182376 163416
rect 182376 163396 182378 163416
rect 182322 163360 182378 163396
rect 181770 162408 181826 162464
rect 182322 161592 182378 161648
rect 181678 160640 181734 160696
rect 180298 158328 180354 158384
rect 181126 154656 181182 154712
rect 181402 153160 181458 153216
rect 182322 159824 182378 159880
rect 182322 158056 182378 158112
rect 181770 157104 181826 157160
rect 182230 156288 182286 156344
rect 182322 156016 182378 156072
rect 181954 153604 181956 153624
rect 181956 153604 182008 153624
rect 182008 153604 182010 153624
rect 181954 153568 182010 153604
rect 182322 152072 182378 152128
rect 182322 150884 182324 150904
rect 182324 150884 182376 150904
rect 182376 150884 182378 150904
rect 182322 150848 182378 150884
rect 182230 150576 182286 150632
rect 180390 148536 180446 148592
rect 182322 148264 182378 148320
rect 192902 144592 192958 144648
rect 196490 144048 196546 144104
rect 196858 144048 196914 144104
rect 197686 143912 197742 143968
rect 203758 144456 203814 144512
rect 200170 141872 200226 141928
rect 225654 160640 225710 160696
rect 211026 143096 211082 143152
rect 207254 141056 207310 141112
rect 219674 142028 219730 142064
rect 219674 142008 219676 142028
rect 219676 142008 219728 142028
rect 219728 142008 219730 142028
rect 197686 135072 197742 135128
rect 225838 155336 225894 155392
rect 226022 154384 226078 154440
rect 225930 153568 225986 153624
rect 225746 152616 225802 152672
rect 226298 163360 226354 163416
rect 226298 162428 226354 162464
rect 226298 162408 226300 162428
rect 226300 162408 226352 162428
rect 226352 162408 226354 162428
rect 226390 161592 226446 161648
rect 226298 159824 226354 159880
rect 226390 158872 226446 158928
rect 226298 158056 226354 158112
rect 226114 151800 226170 151856
rect 226206 150848 226262 150904
rect 225562 150032 225618 150088
rect 225286 149080 225342 149136
rect 225194 148264 225250 148320
rect 226390 157104 226446 157160
rect 226482 156288 226538 156344
rect 176250 108824 176306 108880
rect 178734 84208 178790 84264
rect 182322 84208 182378 84264
rect 139634 75232 139690 75288
rect 173858 75232 173914 75288
rect 174042 74144 174098 74200
rect 139726 73736 139782 73792
rect 139542 72512 139598 72568
rect 139634 71016 139690 71072
rect 172938 73192 172994 73248
rect 173306 72104 173362 72160
rect 139910 71424 139966 71480
rect 139818 69520 139874 69576
rect 139634 68296 139690 68352
rect 139726 67344 139782 67400
rect 139634 67072 139690 67128
rect 174042 71036 174098 71072
rect 174042 71016 174044 71036
rect 174044 71016 174096 71036
rect 174096 71016 174098 71036
rect 174042 70064 174098 70120
rect 172938 68976 172994 69032
rect 173858 67888 173914 67944
rect 139910 65440 139966 65496
rect 139634 64216 139690 64272
rect 139726 63128 139782 63184
rect 139634 61360 139690 61416
rect 139818 62720 139874 62776
rect 139726 60000 139782 60056
rect 173122 61768 173178 61824
rect 173122 60680 173178 60736
rect 173030 59592 173086 59648
rect 140462 58912 140518 58968
rect 140370 58640 140426 58696
rect 140278 57144 140334 57200
rect 173306 57552 173362 57608
rect 140462 56192 140518 56248
rect 174042 66956 174098 66992
rect 174042 66936 174044 66956
rect 174044 66936 174096 66956
rect 174096 66936 174098 66956
rect 181034 69384 181090 69440
rect 226482 69384 226538 69440
rect 180942 68432 180998 68488
rect 225930 68432 225986 68488
rect 173858 65848 173914 65904
rect 173490 64916 173546 64952
rect 173490 64896 173492 64916
rect 173492 64896 173544 64916
rect 173544 64896 173546 64916
rect 173490 63808 173546 63864
rect 174042 62740 174098 62776
rect 174042 62720 174044 62740
rect 174044 62720 174096 62740
rect 174096 62720 174098 62740
rect 173582 58660 173638 58696
rect 173582 58640 173584 58660
rect 173584 58640 173636 58660
rect 173636 58640 173638 58660
rect 173490 56600 173546 56656
rect 181402 67616 181458 67672
rect 226298 67616 226354 67672
rect 180942 64352 180998 64408
rect 181954 66392 182010 66448
rect 182138 65848 182194 65904
rect 181770 64080 181826 64136
rect 182322 63128 182378 63184
rect 182322 62312 182378 62368
rect 181586 61360 181642 61416
rect 181218 60408 181274 60464
rect 181034 59592 181090 59648
rect 181126 58640 181182 58696
rect 181034 57824 181090 57880
rect 181034 56600 181090 56656
rect 181126 56056 181182 56112
rect 173398 55512 173454 55568
rect 140646 55240 140702 55296
rect 140370 54444 140426 54480
rect 140370 54424 140372 54444
rect 140372 54424 140424 54444
rect 140424 54424 140426 54444
rect 173582 54444 173638 54480
rect 173582 54424 173584 54444
rect 173584 54424 173636 54444
rect 173636 54424 173638 54444
rect 181034 55104 181090 55160
rect 226298 66684 226354 66720
rect 226298 66664 226300 66684
rect 226300 66664 226352 66684
rect 226352 66664 226354 66684
rect 226390 65848 226446 65904
rect 226206 64896 226262 64952
rect 225930 64080 225986 64136
rect 225746 63128 225802 63184
rect 226298 62312 226354 62368
rect 226298 61396 226300 61416
rect 226300 61396 226352 61416
rect 226352 61396 226354 61416
rect 226298 61360 226354 61396
rect 225746 60408 225802 60464
rect 226298 59592 226354 59648
rect 225746 58640 225802 58696
rect 225562 57824 225618 57880
rect 226298 56872 226354 56928
rect 225654 56056 225710 56112
rect 226390 55104 226446 55160
rect 181034 54288 181090 54344
rect 140554 53472 140610 53528
rect 173582 53472 173638 53528
rect 140002 52384 140058 52440
rect 171834 52384 171890 52440
rect 173306 51296 173362 51352
rect 142854 51024 142910 51080
rect 140646 50752 140702 50808
rect 140370 50344 140426 50400
rect 140554 48984 140610 49040
rect 140002 48032 140058 48088
rect 147730 48032 147786 48088
rect 153986 48032 154042 48088
rect 160058 47896 160114 47952
rect 163002 46536 163058 46592
rect 168890 47896 168946 47952
rect 166406 47760 166462 47816
rect 167234 47760 167290 47816
rect 167694 47508 167750 47544
rect 167694 47488 167696 47508
rect 167696 47488 167748 47508
rect 167748 47488 167750 47508
rect 169534 45992 169590 46048
rect 169718 46028 169720 46048
rect 169720 46028 169772 46048
rect 169772 46028 169774 46048
rect 169718 45992 169774 46028
rect 165946 45856 166002 45912
rect 163002 45720 163058 45776
rect 170546 50616 170602 50672
rect 173582 50344 173638 50400
rect 172938 49256 172994 49312
rect 173306 48304 173362 48360
rect 181862 47896 181918 47952
rect 182138 49256 182194 49312
rect 182138 46672 182194 46728
rect 88390 26000 88446 26056
rect 88022 23280 88078 23336
rect 181954 45348 181956 45368
rect 181956 45348 182008 45368
rect 182008 45348 182010 45368
rect 181954 45312 182010 45348
rect 181954 33616 182010 33672
rect 182046 30760 182102 30816
rect 182138 28040 182194 28096
rect 191982 51568 192038 51624
rect 187290 50616 187346 50672
rect 199066 46672 199122 46728
rect 203758 51568 203814 51624
rect 207898 51296 207954 51352
rect 212498 53064 212554 53120
rect 212590 47352 212646 47408
rect 207530 37696 207586 37752
rect 226482 54288 226538 54344
rect 182230 26000 182286 26056
rect 181862 23280 181918 23336
rect 88482 20696 88538 20752
rect 182322 20696 182378 20752
rect 13042 15564 13044 15584
rect 13044 15564 13096 15584
rect 13096 15564 13098 15584
rect 13042 15528 13098 15564
rect 284350 393744 284406 393800
rect 233474 357704 233530 357760
rect 233474 356516 233476 356536
rect 233476 356516 233528 356536
rect 233528 356516 233530 356536
rect 233474 356480 233530 356516
rect 233474 355156 233476 355176
rect 233476 355156 233528 355176
rect 233528 355156 233530 355176
rect 233474 355120 233530 355156
rect 233566 354576 233622 354632
rect 233474 353488 233530 353544
rect 233474 352264 233530 352320
rect 233474 350940 233476 350960
rect 233476 350940 233528 350960
rect 233528 350940 233530 350960
rect 233474 350904 233530 350940
rect 233566 350360 233622 350416
rect 233474 349544 233530 349600
rect 233474 348220 233476 348240
rect 233476 348220 233528 348240
rect 233528 348220 233530 348240
rect 233474 348184 233530 348220
rect 233382 346824 233438 346880
rect 233290 346416 233346 346472
rect 233474 345192 233530 345248
rect 233474 343968 233530 344024
rect 234578 342608 234634 342664
rect 234486 342200 234542 342256
rect 234394 341248 234450 341304
rect 233474 339888 233530 339944
rect 233474 338564 233476 338584
rect 233476 338564 233528 338584
rect 233528 338564 233530 338584
rect 233474 338528 233530 338564
rect 233658 338120 233714 338176
rect 233566 337032 233622 337088
rect 233474 335844 233476 335864
rect 233476 335844 233528 335864
rect 233528 335844 233530 335864
rect 233474 335808 233530 335844
rect 234118 334312 234174 334368
rect 234302 333904 234358 333960
rect 231818 333532 231820 333552
rect 231820 333532 231872 333552
rect 231872 333532 231874 333552
rect 230898 332136 230954 332192
rect 230806 331456 230862 331512
rect 231818 333496 231874 333532
rect 233934 332952 233990 333008
rect 231358 332136 231414 332192
rect 231450 331456 231506 331512
rect 233474 331456 233530 331512
rect 233474 330232 233530 330288
rect 252610 330096 252666 330152
rect 251966 329960 252022 330016
rect 230990 320304 231046 320360
rect 231450 317176 231506 317232
rect 231358 314048 231414 314104
rect 230898 310920 230954 310976
rect 230806 307792 230862 307848
rect 230714 298408 230770 298464
rect 230806 294600 230862 294656
rect 230714 234352 230770 234408
rect 230714 234080 230770 234136
rect 230714 223200 230770 223256
rect 231082 289024 231138 289080
rect 230898 237888 230954 237944
rect 230990 220072 231046 220128
rect 230898 216944 230954 217000
rect 230806 200624 230862 200680
rect 230714 197496 230770 197552
rect 231358 285216 231414 285272
rect 231174 234896 231230 234952
rect 231174 234488 231230 234544
rect 231174 226328 231230 226384
rect 232002 304664 232058 304720
rect 232002 301536 232058 301592
rect 231450 279640 231506 279696
rect 231634 282788 231690 282824
rect 231634 282768 231636 282788
rect 231636 282768 231688 282788
rect 231688 282768 231690 282788
rect 231542 276512 231598 276568
rect 256014 327512 256070 327568
rect 240650 310104 240706 310160
rect 240926 296776 240982 296832
rect 240374 283484 240376 283504
rect 240376 283484 240428 283504
rect 240428 283484 240430 283504
rect 240374 283448 240430 283484
rect 232738 274336 232794 274392
rect 231634 273384 231690 273440
rect 233474 263048 233530 263104
rect 233474 261688 233530 261744
rect 233474 260328 233530 260384
rect 233474 258832 233530 258888
rect 233474 257472 233530 257528
rect 232738 254616 232794 254672
rect 233474 256112 233530 256168
rect 233474 253256 233530 253312
rect 233566 251896 233622 251952
rect 233474 250980 233476 251000
rect 233476 250980 233528 251000
rect 233528 250980 233530 251000
rect 233474 250944 233530 250980
rect 232830 249720 232886 249776
rect 233474 248360 233530 248416
rect 233474 245504 233530 245560
rect 233474 242784 233530 242840
rect 233474 240628 233530 240664
rect 233474 240608 233476 240628
rect 233476 240608 233528 240628
rect 233528 240608 233530 240628
rect 233474 239268 233530 239304
rect 233474 239248 233476 239268
rect 233476 239248 233528 239268
rect 233528 239248 233530 239268
rect 234578 246864 234634 246920
rect 234210 244144 234266 244200
rect 234118 238568 234174 238624
rect 233474 237072 233530 237128
rect 247274 274336 247330 274392
rect 247826 273964 247828 273984
rect 247828 273964 247880 273984
rect 247880 273964 247882 273984
rect 247826 273928 247882 273964
rect 250862 274336 250918 274392
rect 252702 274608 252758 274664
rect 252058 274472 252114 274528
rect 250954 273792 251010 273848
rect 253162 274744 253218 274800
rect 261718 306160 261774 306216
rect 261258 286324 261314 286360
rect 261258 286304 261260 286324
rect 261260 286304 261312 286324
rect 261312 286304 261314 286324
rect 244238 236120 244294 236176
rect 230898 194912 230954 194968
rect 231082 194912 231138 194968
rect 230806 107872 230862 107928
rect 230714 104336 230770 104392
rect 231542 216536 231598 216592
rect 231450 207696 231506 207752
rect 231358 185664 231414 185720
rect 231726 213816 231782 213872
rect 231634 210688 231690 210744
rect 231634 204296 231690 204352
rect 231542 191920 231598 191976
rect 232002 188812 232058 188848
rect 241478 233400 241534 233456
rect 242490 235848 242546 235904
rect 246032 235576 246088 235632
rect 246630 234896 246686 234952
rect 243042 233672 243098 233728
rect 239914 232448 239970 232504
rect 246630 233264 246686 233320
rect 262546 235712 262602 235768
rect 240926 216128 240982 216184
rect 242214 207696 242270 207752
rect 242214 204568 242270 204624
rect 237522 204296 237578 204352
rect 240374 202800 240430 202856
rect 242582 201984 242638 202040
rect 242582 192464 242638 192520
rect 240374 189472 240430 189528
rect 232002 188792 232004 188812
rect 232004 188792 232056 188812
rect 232056 188792 232058 188812
rect 231450 182536 231506 182592
rect 230990 179408 231046 179464
rect 248930 183080 248986 183136
rect 249022 182128 249078 182184
rect 251414 180632 251470 180688
rect 251322 180496 251378 180552
rect 250218 180088 250274 180144
rect 249574 179952 249630 180008
rect 252702 180632 252758 180688
rect 253346 180768 253402 180824
rect 261718 212728 261774 212784
rect 262362 192736 262418 192792
rect 233474 169072 233530 169128
rect 233474 167712 233530 167768
rect 236878 167032 236934 167088
rect 233474 166352 233530 166408
rect 233474 164856 233530 164912
rect 233474 163496 233530 163552
rect 233474 162136 233530 162192
rect 232830 155064 232886 155120
rect 233474 160660 233530 160696
rect 233474 160640 233476 160660
rect 233476 160640 233528 160660
rect 233528 160640 233530 160660
rect 233474 159300 233530 159336
rect 233474 159280 233476 159300
rect 233476 159280 233528 159300
rect 233528 159280 233530 159300
rect 233474 157940 233530 157976
rect 233474 157920 233476 157940
rect 233476 157920 233528 157940
rect 233528 157920 233530 157940
rect 233474 156560 233530 156616
rect 234026 153704 234082 153760
rect 232922 152344 232978 152400
rect 233474 150884 233476 150904
rect 233476 150884 233528 150904
rect 233528 150884 233530 150904
rect 233474 150848 233530 150884
rect 232738 149488 232794 149544
rect 233474 148164 233476 148184
rect 233476 148164 233528 148184
rect 233528 148164 233530 148184
rect 233474 148128 233530 148164
rect 233474 146632 233530 146688
rect 233474 145272 233530 145328
rect 233474 143912 233530 143968
rect 233474 142028 233530 142064
rect 233474 142008 233476 142028
rect 233476 142008 233528 142028
rect 233528 142008 233530 142028
rect 230990 139968 231046 140024
rect 231450 139696 231506 139752
rect 231358 132896 231414 132952
rect 231082 129768 231138 129824
rect 230990 123240 231046 123296
rect 230898 99984 230954 100040
rect 231450 125960 231506 126016
rect 231358 98488 231414 98544
rect 232002 109912 232058 109968
rect 231450 92232 231506 92288
rect 232002 94988 232004 95008
rect 232004 94988 232056 95008
rect 232056 94988 232058 95008
rect 232002 94952 232058 94988
rect 231542 88832 231598 88888
rect 231082 85740 231084 85760
rect 231084 85740 231136 85760
rect 231136 85740 231138 85760
rect 231082 85704 231138 85740
rect 242030 142144 242086 142200
rect 241754 139732 241756 139752
rect 241756 139732 241808 139752
rect 241808 139732 241810 139752
rect 241754 139696 241810 139732
rect 261902 142180 261904 142200
rect 261904 142180 261956 142200
rect 261956 142180 261958 142200
rect 261902 142144 261958 142180
rect 243226 141736 243282 141792
rect 244054 139832 244110 139888
rect 242030 129496 242086 129552
rect 246354 139696 246410 139752
rect 246446 130212 246448 130232
rect 246448 130212 246500 130232
rect 246500 130212 246502 130232
rect 246446 130176 246502 130212
rect 249666 138336 249722 138392
rect 249114 135752 249170 135808
rect 249114 134392 249170 134448
rect 252242 138472 252298 138528
rect 242030 124736 242086 124792
rect 240374 122152 240430 122208
rect 240098 109776 240154 109832
rect 240834 108824 240890 108880
rect 242030 100664 242086 100720
rect 242030 95768 242086 95824
rect 240374 95496 240430 95552
rect 248930 89104 248986 89160
rect 250218 88968 250274 89024
rect 249666 88832 249722 88888
rect 251736 88560 251792 88616
rect 251322 86656 251378 86712
rect 252058 86248 252114 86304
rect 249574 86112 249630 86168
rect 253346 86792 253402 86848
rect 262362 118752 262418 118808
rect 261166 98760 261222 98816
rect 233474 75232 233530 75288
rect 233474 73756 233530 73792
rect 233474 73736 233476 73756
rect 233476 73736 233528 73756
rect 233528 73736 233530 73756
rect 233474 72512 233530 72568
rect 233474 71424 233530 71480
rect 233566 71016 233622 71072
rect 233566 69520 233622 69576
rect 233474 67208 233530 67264
rect 233658 68296 233714 68352
rect 234210 66936 234266 66992
rect 233474 64488 233530 64544
rect 234394 65440 234450 65496
rect 233474 63128 233530 63184
rect 233566 62720 233622 62776
rect 233474 61360 233530 61416
rect 233474 60000 233530 60056
rect 233658 58912 233714 58968
rect 233474 58640 233530 58696
rect 233566 57144 233622 57200
rect 233474 56056 233530 56112
rect 233474 55240 233530 55296
rect 233474 54444 233530 54480
rect 233474 54424 233476 54444
rect 233476 54424 233528 54444
rect 233528 54424 233530 54444
rect 233474 53472 233530 53528
rect 233474 52384 233530 52440
rect 233566 50752 233622 50808
rect 233474 50344 233530 50400
rect 233474 48984 233530 49040
rect 238626 48032 238682 48088
rect 233474 47760 233530 47816
rect 250494 47896 250550 47952
rect 248010 47216 248066 47272
rect 244882 45992 244938 46048
rect 260430 48032 260486 48088
rect 262822 48032 262878 48088
rect 257302 47896 257358 47952
rect 262546 45992 262602 46048
rect 262822 45856 262878 45912
rect 319770 393744 319826 393800
rect 302106 393064 302162 393120
rect 319126 384768 319182 384824
rect 319034 382048 319090 382104
rect 267330 357160 267386 357216
rect 267882 356072 267938 356128
rect 267882 355156 267884 355176
rect 267884 355156 267936 355176
rect 267936 355156 267938 355176
rect 267882 355120 267938 355156
rect 267422 354032 267478 354088
rect 267882 352944 267938 353000
rect 267882 351992 267938 352048
rect 274782 351312 274838 351368
rect 267698 350904 267754 350960
rect 267514 349816 267570 349872
rect 285270 367224 285326 367280
rect 284994 351604 285050 351640
rect 284994 351584 284996 351604
rect 284996 351584 285048 351604
rect 285048 351584 285050 351604
rect 274966 350360 275022 350416
rect 274874 349544 274930 349600
rect 267882 348864 267938 348920
rect 267882 347776 267938 347832
rect 275058 348592 275114 348648
rect 267882 346860 267884 346880
rect 267884 346860 267936 346880
rect 267936 346860 267938 346880
rect 267882 346824 267938 346860
rect 274966 346824 275022 346880
rect 275150 347776 275206 347832
rect 274874 346008 274930 346064
rect 267422 345736 267478 345792
rect 267882 344648 267938 344704
rect 266962 344104 267018 344160
rect 267146 344104 267202 344160
rect 266686 343696 266742 343752
rect 274874 345056 274930 345112
rect 275058 344240 275114 344296
rect 267882 342644 267884 342664
rect 267884 342644 267936 342664
rect 267936 342644 267938 342664
rect 267882 342608 267938 342644
rect 267606 341520 267662 341576
rect 274966 341520 275022 341576
rect 267882 340568 267938 340624
rect 274874 340568 274930 340624
rect 267882 339480 267938 339536
rect 267514 337440 267570 337496
rect 267330 336352 267386 336408
rect 267882 338548 267938 338584
rect 267882 338528 267884 338548
rect 267884 338528 267936 338548
rect 267936 338528 267938 338548
rect 267882 335400 267938 335456
rect 267790 334312 267846 334368
rect 267330 333224 267386 333280
rect 274874 338800 274930 338856
rect 275150 343288 275206 343344
rect 275242 342336 275298 342392
rect 275058 339752 275114 339808
rect 274874 337984 274930 338040
rect 274966 337032 275022 337088
rect 274874 336216 274930 336272
rect 267146 332272 267202 332328
rect 266778 331184 266834 331240
rect 267882 330232 267938 330288
rect 282878 333088 282934 333144
rect 296218 333088 296274 333144
rect 296218 332136 296274 332192
rect 292906 331592 292962 331648
rect 306246 333496 306302 333552
rect 319218 380144 319274 380200
rect 319310 377424 319366 377480
rect 319402 374704 319458 374760
rect 319310 333088 319366 333144
rect 320322 372120 320378 372176
rect 328418 357432 328474 357488
rect 328326 356072 328382 356128
rect 328418 355156 328420 355176
rect 328420 355156 328472 355176
rect 328472 355156 328474 355176
rect 328418 355120 328474 355156
rect 328510 354576 328566 354632
rect 328050 353352 328106 353408
rect 328510 352264 328566 352320
rect 320598 351312 320654 351368
rect 321610 350360 321666 350416
rect 320690 349544 320746 349600
rect 321610 348592 321666 348648
rect 321058 347776 321114 347832
rect 320506 346824 320562 346880
rect 321610 346008 321666 346064
rect 327498 350904 327554 350960
rect 327866 350360 327922 350416
rect 327222 349544 327278 349600
rect 327130 348184 327186 348240
rect 327222 346824 327278 346880
rect 327038 346416 327094 346472
rect 320966 345056 321022 345112
rect 321610 344260 321666 344296
rect 321610 344240 321612 344260
rect 321612 344240 321664 344260
rect 321664 344240 321666 344260
rect 321610 343288 321666 343344
rect 328050 345056 328106 345112
rect 326946 342608 327002 342664
rect 321058 342336 321114 342392
rect 321610 341520 321666 341576
rect 320598 340568 320654 340624
rect 320506 339752 320562 339808
rect 320414 338820 320470 338856
rect 320414 338800 320416 338820
rect 320416 338800 320468 338820
rect 320468 338800 320470 338820
rect 320414 337984 320470 338040
rect 320414 337032 320470 337088
rect 320506 336216 320562 336272
rect 319862 333088 319918 333144
rect 328510 343968 328566 344024
rect 328050 342064 328106 342120
rect 327406 341248 327462 341304
rect 327222 339888 327278 339944
rect 327130 338528 327186 338584
rect 327038 338120 327094 338176
rect 326578 334312 326634 334368
rect 327866 337032 327922 337088
rect 327222 335808 327278 335864
rect 326762 333904 326818 333960
rect 319402 331592 319458 331648
rect 319678 331592 319734 331648
rect 319586 330232 319642 330288
rect 270274 313504 270330 313560
rect 270366 296776 270422 296832
rect 269262 280184 269318 280240
rect 266594 256112 266650 256168
rect 266594 254616 266650 254672
rect 266594 253256 266650 253312
rect 266594 251896 266650 251952
rect 266594 249040 266650 249096
rect 266594 247680 266650 247736
rect 266594 244824 266650 244880
rect 266594 243464 266650 243520
rect 266778 239248 266834 239304
rect 267422 263048 267478 263104
rect 267330 258832 267386 258888
rect 267330 250536 267386 250592
rect 267514 261688 267570 261744
rect 267606 260328 267662 260384
rect 267790 257472 267846 257528
rect 267882 246320 267938 246376
rect 267882 242140 267884 242160
rect 267884 242140 267936 242160
rect 267936 242140 267938 242160
rect 267882 242104 267938 242140
rect 267882 240628 267938 240664
rect 267882 240608 267884 240628
rect 267884 240608 267936 240628
rect 267936 240608 267938 240628
rect 267606 237888 267662 237944
rect 267238 236528 267294 236584
rect 276162 257336 276218 257392
rect 321058 257336 321114 257392
rect 274966 256384 275022 256440
rect 274874 255568 274930 255624
rect 274874 252848 274930 252904
rect 274874 249992 274930 250048
rect 275794 254616 275850 254672
rect 275610 252032 275666 252088
rect 275518 251080 275574 251136
rect 274874 248804 274876 248824
rect 274876 248804 274928 248824
rect 274928 248804 274930 248824
rect 274874 248768 274930 248804
rect 274966 248224 275022 248280
rect 274874 247272 274930 247328
rect 274874 246048 274930 246104
rect 274966 245504 275022 245560
rect 274874 244552 274930 244608
rect 275426 243364 275428 243384
rect 275428 243364 275480 243384
rect 275480 243364 275482 243384
rect 275426 243328 275482 243364
rect 275702 250264 275758 250320
rect 275886 253800 275942 253856
rect 321058 256384 321114 256440
rect 321610 255568 321666 255624
rect 320598 254616 320654 254672
rect 321610 253800 321666 253856
rect 320506 252848 320562 252904
rect 321610 252032 321666 252088
rect 321610 251080 321666 251136
rect 321058 250264 321114 250320
rect 321610 249312 321666 249368
rect 321610 248360 321666 248416
rect 321794 247564 321850 247600
rect 321794 247544 321796 247564
rect 321796 247544 321848 247564
rect 321848 247544 321850 247564
rect 321426 246592 321482 246648
rect 321610 245776 321666 245832
rect 321702 244860 321704 244880
rect 321704 244860 321756 244880
rect 321756 244860 321758 244880
rect 321702 244824 321758 244860
rect 321610 244008 321666 244064
rect 321610 243056 321666 243112
rect 275978 242784 276034 242840
rect 320506 242240 320562 242296
rect 283246 239384 283302 239440
rect 294194 239792 294250 239848
rect 290054 238432 290110 238488
rect 286926 236256 286982 236312
rect 305142 240336 305198 240392
rect 301094 234896 301150 234952
rect 324554 320304 324610 320360
rect 324738 317176 324794 317232
rect 327314 332952 327370 333008
rect 328510 331456 328566 331512
rect 325198 310920 325254 310976
rect 325106 305480 325162 305536
rect 325106 298408 325162 298464
rect 324554 292152 324610 292208
rect 322990 226328 323046 226384
rect 272942 219528 272998 219584
rect 272942 202800 272998 202856
rect 273126 186208 273182 186264
rect 267146 164856 267202 164912
rect 267054 162136 267110 162192
rect 266594 160676 266596 160696
rect 266596 160676 266648 160696
rect 266648 160676 266650 160696
rect 266594 160640 266650 160676
rect 266594 159300 266650 159336
rect 266594 159280 266596 159300
rect 266596 159280 266648 159300
rect 266648 159280 266650 159300
rect 266594 157956 266596 157976
rect 266596 157956 266648 157976
rect 266648 157956 266650 157976
rect 266594 157920 266650 157956
rect 266594 155064 266650 155120
rect 266870 153704 266926 153760
rect 266962 152344 267018 152400
rect 266594 150868 266650 150904
rect 266594 150848 266596 150868
rect 266596 150848 266648 150868
rect 266648 150848 266650 150868
rect 266594 149488 266650 149544
rect 266594 148164 266596 148184
rect 266596 148164 266648 148184
rect 266648 148164 266650 148184
rect 266594 148128 266650 148164
rect 266778 145272 266834 145328
rect 267422 169072 267478 169128
rect 267330 156560 267386 156616
rect 267238 142552 267294 142608
rect 267698 167712 267754 167768
rect 267514 166352 267570 166408
rect 267882 163496 267938 163552
rect 274506 163360 274562 163416
rect 274138 158872 274194 158928
rect 274322 150576 274378 150632
rect 274230 149488 274286 149544
rect 321610 163360 321666 163416
rect 274874 162408 274930 162464
rect 320966 162408 321022 162464
rect 274874 161592 274930 161648
rect 274874 160660 274930 160696
rect 274874 160640 274876 160660
rect 274876 160640 274928 160660
rect 274928 160640 274930 160660
rect 320782 160640 320838 160696
rect 321794 161864 321850 161920
rect 275702 159824 275758 159880
rect 321702 159824 321758 159880
rect 275518 158056 275574 158112
rect 274966 156288 275022 156344
rect 274874 156016 274930 156072
rect 274874 154928 274930 154984
rect 274874 153604 274876 153624
rect 274876 153604 274928 153624
rect 274928 153604 274930 153624
rect 274874 153568 274930 153604
rect 274966 153296 275022 153352
rect 274874 152072 274930 152128
rect 274874 150884 274876 150904
rect 274876 150884 274928 150904
rect 274928 150884 274930 150904
rect 274874 150848 274930 150884
rect 274414 148808 274470 148864
rect 275610 157104 275666 157160
rect 267882 146632 267938 146688
rect 321058 158872 321114 158928
rect 321610 158056 321666 158112
rect 321610 157104 321666 157160
rect 321610 156288 321666 156344
rect 321610 155336 321666 155392
rect 320874 154384 320930 154440
rect 321610 153568 321666 153624
rect 320506 152616 320562 152672
rect 320782 151800 320838 151856
rect 321058 150848 321114 150904
rect 321610 150032 321666 150088
rect 321610 149080 321666 149136
rect 321702 148264 321758 148320
rect 267790 143912 267846 143968
rect 283154 138472 283210 138528
rect 284442 138472 284498 138528
rect 290514 144456 290570 144512
rect 294286 143096 294342 143152
rect 301094 141056 301150 141112
rect 296954 137792 297010 137848
rect 285914 135752 285970 135808
rect 286742 135752 286798 135808
rect 270366 125416 270422 125472
rect 269998 108824 270054 108880
rect 270366 92232 270422 92288
rect 266594 75232 266650 75288
rect 266594 74144 266650 74200
rect 266594 73192 266650 73248
rect 266686 72104 266742 72160
rect 266594 71036 266650 71072
rect 266594 71016 266596 71036
rect 266596 71016 266648 71036
rect 266648 71016 266650 71036
rect 266594 70064 266650 70120
rect 266594 68976 266650 69032
rect 266686 67888 266742 67944
rect 266594 66936 266650 66992
rect 266594 65848 266650 65904
rect 266594 64896 266650 64952
rect 266686 63808 266742 63864
rect 266594 62740 266650 62776
rect 266594 62720 266596 62740
rect 266596 62720 266648 62740
rect 266648 62720 266650 62740
rect 266594 61768 266650 61824
rect 266594 60680 266650 60736
rect 274690 68432 274746 68488
rect 267330 59592 267386 59648
rect 267882 58660 267938 58696
rect 267882 58640 267884 58660
rect 267884 58640 267936 58660
rect 267936 58640 267938 58660
rect 267698 57552 267754 57608
rect 267330 56600 267386 56656
rect 267238 55512 267294 55568
rect 267882 54444 267938 54480
rect 267882 54424 267884 54444
rect 267884 54424 267936 54444
rect 267936 54424 267938 54444
rect 274874 69384 274930 69440
rect 274782 67616 274838 67672
rect 274874 66700 274876 66720
rect 274876 66700 274928 66720
rect 274928 66700 274930 66720
rect 274874 66664 274930 66700
rect 321702 69384 321758 69440
rect 321610 68432 321666 68488
rect 321610 67616 321666 67672
rect 321242 66664 321298 66720
rect 274966 65848 275022 65904
rect 321610 65848 321666 65904
rect 274690 64896 274746 64952
rect 274230 63128 274286 63184
rect 321610 64896 321666 64952
rect 274874 64080 274930 64136
rect 321610 64116 321612 64136
rect 321612 64116 321664 64136
rect 321664 64116 321666 64136
rect 321610 64080 321666 64116
rect 320506 62720 320562 62776
rect 274782 62312 274838 62368
rect 318390 61768 318446 61824
rect 320690 61532 320692 61552
rect 320692 61532 320744 61552
rect 320744 61532 320746 61552
rect 320690 61496 320746 61532
rect 274966 61360 275022 61416
rect 318390 61360 318446 61416
rect 321058 61360 321114 61416
rect 274874 60408 274930 60464
rect 321058 59864 321114 59920
rect 275702 59592 275758 59648
rect 320506 59592 320562 59648
rect 275426 58640 275482 58696
rect 320414 58640 320470 58696
rect 275702 57824 275758 57880
rect 320414 57844 320470 57880
rect 320414 57824 320416 57844
rect 320416 57824 320468 57844
rect 320468 57824 320470 57844
rect 275702 56872 275758 56928
rect 275242 56056 275298 56112
rect 275426 55104 275482 55160
rect 320506 56872 320562 56928
rect 320414 56056 320470 56112
rect 320414 55104 320470 55160
rect 275702 54324 275704 54344
rect 275704 54324 275756 54344
rect 275756 54324 275758 54344
rect 275702 54288 275758 54324
rect 320414 54288 320470 54344
rect 267882 53472 267938 53528
rect 267882 52384 267938 52440
rect 267514 51296 267570 51352
rect 281314 51296 281370 51352
rect 266778 50344 266834 50400
rect 267882 49256 267938 49312
rect 267882 48304 267938 48360
rect 275794 47896 275850 47952
rect 276070 47896 276126 47952
rect 275978 46536 276034 46592
rect 275886 33616 275942 33672
rect 275978 30760 276034 30816
rect 275794 28040 275850 28096
rect 283706 48032 283762 48088
rect 284350 48032 284406 48088
rect 286006 47372 286062 47408
rect 286006 47352 286008 47372
rect 286008 47352 286060 47372
rect 286060 47352 286062 47372
rect 301646 53064 301702 53120
rect 306614 53064 306670 53120
rect 306614 47352 306670 47408
rect 301554 37696 301610 37752
rect 325290 292152 325346 292208
rect 325290 285896 325346 285952
rect 324646 234352 324702 234408
rect 324738 226348 324794 226384
rect 324738 226328 324740 226348
rect 324740 226328 324792 226348
rect 324792 226328 324794 226348
rect 324646 223200 324702 223256
rect 324922 213816 324978 213872
rect 324554 198720 324610 198776
rect 324554 188792 324610 188848
rect 324554 179408 324610 179464
rect 324646 132488 324702 132544
rect 324554 132352 324610 132408
rect 324646 125960 324702 126016
rect 325106 129768 325162 129824
rect 324738 123240 324794 123296
rect 324554 119876 324556 119896
rect 324556 119876 324608 119896
rect 324608 119876 324610 119896
rect 324554 119840 324610 119876
rect 324554 117256 324610 117312
rect 325474 305480 325530 305536
rect 325566 305344 325622 305400
rect 325842 314048 325898 314104
rect 325750 307792 325806 307848
rect 325658 301536 325714 301592
rect 325382 279640 325438 279696
rect 325474 276512 325530 276568
rect 325842 282804 325844 282824
rect 325844 282804 325896 282824
rect 325896 282804 325898 282824
rect 325842 282768 325898 282804
rect 325566 273384 325622 273440
rect 325842 239656 325898 239712
rect 325474 207560 325530 207616
rect 339182 327376 339238 327432
rect 340010 327376 340066 327432
rect 334214 309716 334270 309752
rect 334214 309696 334216 309716
rect 334216 309696 334268 309716
rect 334268 309696 334270 309716
rect 352798 297184 352854 297240
rect 353994 297184 354050 297240
rect 334214 296232 334270 296288
rect 334214 283584 334270 283640
rect 352062 266720 352118 266776
rect 350958 266584 351014 266640
rect 354270 285216 354326 285272
rect 356202 314048 356258 314104
rect 356202 308608 356258 308664
rect 356202 304140 356258 304176
rect 356202 304120 356204 304140
rect 356204 304120 356256 304140
rect 356256 304120 356258 304140
rect 356202 298816 356258 298872
rect 356202 293804 356258 293840
rect 356202 293784 356204 293804
rect 356204 293784 356256 293804
rect 356256 293784 356258 293804
rect 356202 289024 356258 289080
rect 356202 283720 356258 283776
rect 356202 279368 356258 279424
rect 328418 263456 328474 263512
rect 327682 261688 327738 261744
rect 327958 260328 328014 260384
rect 327222 258832 327278 258888
rect 327130 257472 327186 257528
rect 328510 256112 328566 256168
rect 328418 254616 328474 254672
rect 327130 253256 327186 253312
rect 327222 251896 327278 251952
rect 327222 250536 327278 250592
rect 328418 249076 328420 249096
rect 328420 249076 328472 249096
rect 328472 249076 328474 249096
rect 328418 249040 328474 249076
rect 328418 247700 328474 247736
rect 328418 247680 328420 247700
rect 328420 247680 328472 247700
rect 328472 247680 328474 247700
rect 328418 246864 328474 246920
rect 327866 245504 327922 245560
rect 327866 244008 327922 244064
rect 327866 242648 327922 242704
rect 327222 240608 327278 240664
rect 328050 239248 328106 239304
rect 327866 238568 327922 238624
rect 328418 236564 328420 236584
rect 328420 236564 328472 236584
rect 328472 236564 328474 236584
rect 328418 236528 328474 236564
rect 325750 220072 325806 220128
rect 325842 216944 325898 217000
rect 325658 210688 325714 210744
rect 325566 204432 325622 204488
rect 325382 191920 325438 191976
rect 325290 185664 325346 185720
rect 350958 232448 351014 232504
rect 352062 232448 352118 232504
rect 334214 216128 334270 216184
rect 334214 202800 334270 202856
rect 334214 189472 334270 189528
rect 325474 182536 325530 182592
rect 350958 172608 351014 172664
rect 352062 172608 352118 172664
rect 352798 191376 352854 191432
rect 352798 184032 352854 184088
rect 352890 182128 352946 182184
rect 352982 181992 353038 182048
rect 355098 220208 355154 220264
rect 356294 215856 356350 215912
rect 356202 215176 356258 215232
rect 356202 210144 356258 210200
rect 356202 205248 356258 205304
rect 356202 200216 356258 200272
rect 356202 195184 356258 195240
rect 356202 190152 356258 190208
rect 356202 185256 356258 185312
rect 358042 219936 358098 219992
rect 358226 219936 358282 219992
rect 429434 390480 429490 390536
rect 429434 377968 429490 378024
rect 360618 259104 360674 259160
rect 360526 255976 360582 256032
rect 360802 262232 360858 262288
rect 361170 255976 361226 256032
rect 360710 252848 360766 252904
rect 361170 252848 361226 252904
rect 360710 249720 360766 249776
rect 358410 211640 358466 211696
rect 358594 211640 358650 211696
rect 328418 169072 328474 169128
rect 327222 167712 327278 167768
rect 328418 166352 328474 166408
rect 328510 164856 328566 164912
rect 327222 163360 327278 163416
rect 360802 246592 360858 246648
rect 360894 243464 360950 243520
rect 360986 240336 361042 240392
rect 361262 237344 361318 237400
rect 359054 168256 359110 168312
rect 359698 168256 359754 168312
rect 328418 162136 328474 162192
rect 327314 160640 327370 160696
rect 327222 159280 327278 159336
rect 327222 157920 327278 157976
rect 327222 156560 327278 156616
rect 328418 155084 328474 155120
rect 328418 155064 328420 155084
rect 328420 155064 328472 155084
rect 328472 155064 328474 155084
rect 328418 153740 328420 153760
rect 328420 153740 328472 153760
rect 328472 153740 328474 153760
rect 328418 153704 328474 153740
rect 328418 152380 328420 152400
rect 328420 152380 328472 152400
rect 328472 152380 328474 152400
rect 328418 152344 328474 152380
rect 328418 150884 328420 150904
rect 328420 150884 328472 150904
rect 328472 150884 328474 150904
rect 328418 150848 328474 150884
rect 328418 149524 328420 149544
rect 328420 149524 328472 149544
rect 328472 149524 328474 149544
rect 328418 149488 328474 149524
rect 327222 146632 327278 146688
rect 328418 148164 328420 148184
rect 328420 148164 328472 148184
rect 328472 148164 328474 148184
rect 328418 148128 328474 148164
rect 327866 145272 327922 145328
rect 327314 143912 327370 143968
rect 327314 141872 327370 141928
rect 325198 98488 325254 98544
rect 324554 94952 324610 95008
rect 325474 113584 325530 113640
rect 325382 110864 325438 110920
rect 325290 92232 325346 92288
rect 325382 88832 325438 88888
rect 350958 139560 351014 139616
rect 352062 139560 352118 139616
rect 334214 122152 334270 122208
rect 334214 108824 334270 108880
rect 334214 95496 334270 95552
rect 326578 86656 326634 86712
rect 324554 85704 324610 85760
rect 350958 77816 351014 77872
rect 352062 77816 352118 77872
rect 352798 97828 352854 97864
rect 352798 97808 352800 97828
rect 352800 97808 352852 97828
rect 352852 97808 352854 97828
rect 352798 90056 352854 90112
rect 356202 126232 356258 126288
rect 356202 121200 356258 121256
rect 356202 116168 356258 116224
rect 356202 111272 356258 111328
rect 356202 106240 356258 106296
rect 356202 101208 356258 101264
rect 356202 96176 356258 96232
rect 356202 91280 356258 91336
rect 360434 165128 360490 165184
rect 360526 162000 360582 162056
rect 360618 158872 360674 158928
rect 360710 155744 360766 155800
rect 360802 152616 360858 152672
rect 360986 149488 361042 149544
rect 360894 146360 360950 146416
rect 429434 365456 429490 365512
rect 430078 352944 430134 353000
rect 429434 340432 429490 340488
rect 361262 165128 361318 165184
rect 361262 158872 361318 158928
rect 361170 155744 361226 155800
rect 361078 143368 361134 143424
rect 358318 124736 358374 124792
rect 358502 124736 358558 124792
rect 328418 75232 328474 75288
rect 328326 74144 328382 74200
rect 327222 72512 327278 72568
rect 327038 71424 327094 71480
rect 327130 69520 327186 69576
rect 326946 66936 327002 66992
rect 328510 71016 328566 71072
rect 327222 68296 327278 68352
rect 327130 65440 327186 65496
rect 328234 67208 328290 67264
rect 327314 64488 327370 64544
rect 327222 62720 327278 62776
rect 328418 63128 328474 63184
rect 328326 61360 328382 61416
rect 327498 58640 327554 58696
rect 328418 60000 328474 60056
rect 328602 58912 328658 58968
rect 328418 57144 328474 57200
rect 327498 55920 327554 55976
rect 328510 55240 328566 55296
rect 328418 54444 328474 54480
rect 328418 54424 328420 54444
rect 328420 54424 328472 54444
rect 328472 54424 328474 54444
rect 328418 53472 328474 53528
rect 328510 52384 328566 52440
rect 327682 50888 327738 50944
rect 328418 50344 328474 50400
rect 358594 50344 358650 50400
rect 328418 49256 328474 49312
rect 327866 47896 327922 47952
rect 276070 26000 276126 26056
rect 275518 23280 275574 23336
rect 276162 20696 276218 20752
rect 343138 45992 343194 46048
rect 358502 47488 358558 47544
rect 369174 236528 369230 236584
rect 368714 234080 368770 234136
rect 368714 233708 368716 233728
rect 368716 233708 368768 233728
rect 368768 233708 368770 233728
rect 368714 233672 368770 233708
rect 368806 233400 368862 233456
rect 368714 232992 368770 233048
rect 368714 232176 368770 232232
rect 368806 231768 368862 231824
rect 368898 231360 368954 231416
rect 368806 230952 368862 231008
rect 368714 230544 368770 230600
rect 368898 230136 368954 230192
rect 368714 229456 368770 229512
rect 368806 229048 368862 229104
rect 368714 228640 368770 228696
rect 368714 228268 368716 228288
rect 368716 228268 368768 228288
rect 368768 228268 368770 228288
rect 368714 228232 368770 228268
rect 368806 227416 368862 227472
rect 368714 227008 368770 227064
rect 369082 226464 369138 226520
rect 368898 226328 368954 226384
rect 368806 225920 368862 225976
rect 368714 225548 368716 225568
rect 368716 225548 368768 225568
rect 368768 225548 368770 225568
rect 368714 225512 368770 225548
rect 368806 225104 368862 225160
rect 368714 224696 368770 224752
rect 368898 224288 368954 224344
rect 368806 223880 368862 223936
rect 368714 223200 368770 223256
rect 368806 222384 368862 222440
rect 368714 221568 368770 221624
rect 369450 236120 369506 236176
rect 369082 222792 369138 222848
rect 369082 221976 369138 222032
rect 368990 221160 369046 221216
rect 368806 220752 368862 220808
rect 368714 220344 368770 220400
rect 368714 219664 368770 219720
rect 368990 219256 369046 219312
rect 368806 218848 368862 218904
rect 368714 218032 368770 218088
rect 368806 217216 368862 217272
rect 369082 217624 369138 217680
rect 369082 217488 369138 217544
rect 368990 216536 369046 216592
rect 368714 216128 368770 216184
rect 368714 215756 368716 215776
rect 368716 215756 368768 215776
rect 368768 215756 368770 215776
rect 368714 215720 368770 215756
rect 368714 214904 368770 214960
rect 368806 214496 368862 214552
rect 368714 213680 368770 213736
rect 367978 213272 368034 213328
rect 368714 213036 368716 213056
rect 368716 213036 368768 213056
rect 368768 213036 368770 213056
rect 368714 213000 368770 213036
rect 368898 214088 368954 214144
rect 369266 219936 369322 219992
rect 369174 215312 369230 215368
rect 368530 173016 368586 173072
rect 368714 173016 368770 173072
rect 369358 216808 369414 216864
rect 369634 235712 369690 235768
rect 369542 229864 369598 229920
rect 369542 227824 369598 227880
rect 369818 235304 369874 235360
rect 369726 232584 369782 232640
rect 405974 315852 405976 315872
rect 405976 315852 406028 315872
rect 406028 315852 406030 315872
rect 405974 315816 406030 315852
rect 429434 315408 429490 315464
rect 427318 313776 427374 313832
rect 405974 313640 406030 313696
rect 405974 310376 406030 310432
rect 405974 308236 405976 308256
rect 405976 308236 406028 308256
rect 406028 308236 406030 308256
rect 405974 308200 406030 308236
rect 406066 306196 406068 306216
rect 406068 306196 406120 306216
rect 406120 306196 406122 306216
rect 406066 306160 406122 306196
rect 405974 303576 406030 303632
rect 405974 300448 406030 300504
rect 405974 298272 406030 298328
rect 405974 295416 406030 295472
rect 405974 293648 406030 293704
rect 405974 290656 406030 290712
rect 427226 289044 427282 289080
rect 427226 289024 427228 289044
rect 427228 289024 427280 289044
rect 427280 289024 427282 289044
rect 406066 288616 406122 288672
rect 405974 285508 406030 285544
rect 405974 285488 405976 285508
rect 405976 285488 406028 285508
rect 406028 285488 406030 285508
rect 405974 283312 406030 283368
rect 405974 278688 406030 278744
rect 370002 234896 370058 234952
rect 369910 234488 369966 234544
rect 369726 226600 369782 226656
rect 369818 223472 369874 223528
rect 406618 221568 406674 221624
rect 405974 218712 406030 218768
rect 370094 218440 370150 218496
rect 370094 217488 370150 217544
rect 405974 214108 406030 214144
rect 405974 214088 405976 214108
rect 405976 214088 406028 214108
rect 406028 214088 406030 214108
rect 428698 308608 428754 308664
rect 427410 304120 427466 304176
rect 427502 298680 427558 298736
rect 427594 293648 427650 293704
rect 427686 284264 427742 284320
rect 427870 279368 427926 279424
rect 429434 290404 429490 290440
rect 429434 290384 429436 290404
rect 429436 290384 429488 290404
rect 429488 290384 429490 290404
rect 430170 327920 430226 327976
rect 430170 302896 430226 302952
rect 430262 277872 430318 277928
rect 429434 265360 429490 265416
rect 429434 252848 429490 252904
rect 429526 240336 429582 240392
rect 428698 227824 428754 227880
rect 427410 220208 427466 220264
rect 405974 210980 406030 211016
rect 405974 210960 405976 210980
rect 405976 210960 406028 210980
rect 406028 210960 406030 210980
rect 427318 210144 427374 210200
rect 405974 209464 406030 209520
rect 405974 206780 405976 206800
rect 405976 206780 406028 206800
rect 406028 206780 406030 206800
rect 405974 206744 406030 206780
rect 406066 204568 406122 204624
rect 405974 201324 406030 201360
rect 405974 201304 405976 201324
rect 405976 201304 406028 201324
rect 406028 201304 406030 201324
rect 427134 200216 427190 200272
rect 405974 199128 406030 199184
rect 405974 195864 406030 195920
rect 406066 194504 406122 194560
rect 405974 191668 406030 191704
rect 405974 191648 405976 191668
rect 405976 191648 406028 191668
rect 406028 191648 406030 191668
rect 405974 189472 406030 189528
rect 405974 186208 406030 186264
rect 427226 185428 427228 185448
rect 427228 185428 427280 185448
rect 427280 185428 427282 185448
rect 427226 185392 427282 185428
rect 405974 183896 406030 183952
rect 405974 126912 406030 126968
rect 427318 126232 427374 126288
rect 405974 125552 406030 125608
rect 405974 122596 405976 122616
rect 405976 122596 406028 122616
rect 406028 122596 406030 122616
rect 405974 122560 406030 122596
rect 405974 120556 405976 120576
rect 405976 120556 406028 120576
rect 406028 120556 406030 120576
rect 405974 120520 406030 120556
rect 405974 117392 406030 117448
rect 405974 114808 406030 114864
rect 405974 112632 406030 112688
rect 406066 110592 406122 110648
rect 405974 107600 406030 107656
rect 405974 105288 406030 105344
rect 405974 102160 406030 102216
rect 405974 100564 405976 100584
rect 405976 100564 406028 100584
rect 406028 100564 406030 100584
rect 405974 100528 406030 100564
rect 405974 97672 406030 97728
rect 427226 96176 427282 96232
rect 405974 95496 406030 95552
rect 405974 92368 406030 92424
rect 405974 90212 406030 90248
rect 405974 90192 405976 90212
rect 405976 90192 406028 90212
rect 406028 90192 406030 90212
rect 412874 86656 412930 86712
rect 429710 215312 429766 215368
rect 428698 215176 428754 215232
rect 427502 205248 427558 205304
rect 427594 195184 427650 195240
rect 430078 202800 430134 202856
rect 429894 177776 429950 177832
rect 428790 165264 428846 165320
rect 429434 152752 429490 152808
rect 429526 140240 429582 140296
rect 428698 127728 428754 127784
rect 427502 121200 427558 121256
rect 427410 101208 427466 101264
rect 428698 116168 428754 116224
rect 427594 111272 427650 111328
rect 427594 106240 427650 106296
rect 427594 91552 427650 91608
rect 429434 115216 429490 115272
rect 429434 102724 429490 102760
rect 429434 102704 429436 102724
rect 429436 102704 429488 102724
rect 429488 102704 429490 102724
rect 429526 77680 429582 77736
rect 430170 90192 430226 90248
rect 430078 65168 430134 65224
rect 428790 52656 428846 52712
rect 428698 40144 428754 40200
rect 429802 27632 429858 27688
rect 429434 15120 429490 15176
<< metal3 >>
rect 280246 393740 280252 393804
rect 280316 393802 280322 393804
rect 284345 393802 284411 393805
rect 280316 393800 284411 393802
rect 280316 393744 284350 393800
rect 284406 393744 284411 393800
rect 280316 393742 284411 393744
rect 280316 393740 280322 393742
rect 284345 393739 284411 393742
rect 319765 393802 319831 393805
rect 323118 393802 323124 393804
rect 319765 393800 323124 393802
rect 319765 393744 319770 393800
rect 319826 393744 323124 393800
rect 319765 393742 323124 393744
rect 319765 393739 319831 393742
rect 323118 393740 323124 393742
rect 323188 393740 323194 393804
rect 302101 393122 302167 393125
rect 323486 393122 323492 393124
rect 302101 393120 323492 393122
rect 302101 393064 302106 393120
rect 302162 393064 323492 393120
rect 302101 393062 323492 393064
rect 302101 393059 302167 393062
rect 323486 393060 323492 393062
rect 323556 393060 323562 393124
rect 429429 390538 429495 390541
rect 434416 390538 434896 390568
rect 429429 390536 434896 390538
rect 429429 390480 429434 390536
rect 429490 390480 434896 390536
rect 429429 390478 434896 390480
rect 429429 390475 429495 390478
rect 434416 390448 434896 390478
rect 9896 390130 10376 390160
rect 13313 390130 13379 390133
rect 9896 390128 13379 390130
rect 9896 390072 13318 390128
rect 13374 390072 13379 390128
rect 9896 390070 13379 390072
rect 9896 390040 10376 390070
rect 13313 390067 13379 390070
rect 128638 384826 128698 385408
rect 131349 384826 131415 384829
rect 128638 384824 131415 384826
rect 128638 384768 131354 384824
rect 131410 384768 131415 384824
rect 128638 384766 131415 384768
rect 222662 384826 222722 385408
rect 225189 384826 225255 384829
rect 222662 384824 225255 384826
rect 222662 384768 225194 384824
rect 225250 384768 225255 384824
rect 222662 384766 225255 384768
rect 316686 384826 316746 385408
rect 319121 384826 319187 384829
rect 316686 384824 319187 384826
rect 316686 384768 319126 384824
rect 319182 384768 319187 384824
rect 316686 384766 319187 384768
rect 131349 384763 131415 384766
rect 225189 384763 225255 384766
rect 319121 384763 319187 384766
rect 226477 382786 226543 382789
rect 222692 382784 226543 382786
rect 222692 382728 226482 382784
rect 226538 382728 226543 382784
rect 222692 382726 226543 382728
rect 226477 382723 226543 382726
rect 128638 382106 128698 382688
rect 131441 382106 131507 382109
rect 128638 382104 131507 382106
rect 128638 382048 131446 382104
rect 131502 382048 131507 382104
rect 128638 382046 131507 382048
rect 316686 382106 316746 382688
rect 319029 382106 319095 382109
rect 316686 382104 319095 382106
rect 316686 382048 319034 382104
rect 319090 382048 319095 382104
rect 316686 382046 319095 382048
rect 131441 382043 131507 382046
rect 319029 382043 319095 382046
rect 131533 380202 131599 380205
rect 225281 380202 225347 380205
rect 319213 380202 319279 380205
rect 128668 380200 131599 380202
rect 128668 380144 131538 380200
rect 131594 380144 131599 380200
rect 128668 380142 131599 380144
rect 222692 380200 225347 380202
rect 222692 380144 225286 380200
rect 225342 380144 225347 380200
rect 222692 380142 225347 380144
rect 316716 380200 319279 380202
rect 316716 380144 319218 380200
rect 319274 380144 319279 380200
rect 316716 380142 319279 380144
rect 131533 380139 131599 380142
rect 225281 380139 225347 380142
rect 319213 380139 319279 380142
rect 429429 378026 429495 378029
rect 434416 378026 434896 378056
rect 429429 378024 434896 378026
rect 429429 377968 429434 378024
rect 429490 377968 434896 378024
rect 429429 377966 434896 377968
rect 429429 377963 429495 377966
rect 434416 377936 434896 377966
rect 131625 377482 131691 377485
rect 225373 377482 225439 377485
rect 319305 377482 319371 377485
rect 128668 377480 131691 377482
rect 128668 377424 131630 377480
rect 131686 377424 131691 377480
rect 128668 377422 131691 377424
rect 222692 377480 225439 377482
rect 222692 377424 225378 377480
rect 225434 377424 225439 377480
rect 222692 377422 225439 377424
rect 316716 377480 319371 377482
rect 316716 377424 319310 377480
rect 319366 377424 319371 377480
rect 316716 377422 319371 377424
rect 131625 377419 131691 377422
rect 225373 377419 225439 377422
rect 319305 377419 319371 377422
rect 9896 376802 10376 376832
rect 13589 376802 13655 376805
rect 9896 376800 13655 376802
rect 9896 376744 13594 376800
rect 13650 376744 13655 376800
rect 9896 376742 13655 376744
rect 9896 376712 10376 376742
rect 13589 376739 13655 376742
rect 131717 374762 131783 374765
rect 226477 374762 226543 374765
rect 319397 374762 319463 374765
rect 128668 374760 131783 374762
rect 128668 374704 131722 374760
rect 131778 374704 131783 374760
rect 128668 374702 131783 374704
rect 222692 374760 226543 374762
rect 222692 374704 226482 374760
rect 226538 374704 226543 374760
rect 222692 374702 226543 374704
rect 316716 374760 319463 374762
rect 316716 374704 319402 374760
rect 319458 374704 319463 374760
rect 316716 374702 319463 374704
rect 131717 374699 131783 374702
rect 226477 374699 226543 374702
rect 319397 374699 319463 374702
rect 131809 372178 131875 372181
rect 225833 372178 225899 372181
rect 320317 372178 320383 372181
rect 128668 372176 131875 372178
rect 128668 372120 131814 372176
rect 131870 372120 131875 372176
rect 128668 372118 131875 372120
rect 222692 372176 225899 372178
rect 222692 372120 225838 372176
rect 225894 372120 225899 372176
rect 222692 372118 225899 372120
rect 316716 372176 320383 372178
rect 316716 372120 320322 372176
rect 320378 372120 320383 372176
rect 316716 372118 320383 372120
rect 131809 372115 131875 372118
rect 225833 372115 225899 372118
rect 320317 372115 320383 372118
rect 97350 367220 97356 367284
rect 97420 367282 97426 367284
rect 97493 367282 97559 367285
rect 97420 367280 97559 367282
rect 97420 367224 97498 367280
rect 97554 367224 97559 367280
rect 97420 367222 97559 367224
rect 97420 367220 97426 367222
rect 97493 367219 97559 367222
rect 285030 367220 285036 367284
rect 285100 367282 285106 367284
rect 285265 367282 285331 367285
rect 285100 367280 285331 367282
rect 285100 367224 285270 367280
rect 285326 367224 285331 367280
rect 285100 367222 285331 367224
rect 285100 367220 285106 367222
rect 285265 367219 285331 367222
rect 429429 365514 429495 365517
rect 434416 365514 434896 365544
rect 429429 365512 434896 365514
rect 429429 365456 429434 365512
rect 429490 365456 434896 365512
rect 429429 365454 434896 365456
rect 429429 365451 429495 365454
rect 434416 365424 434896 365454
rect 9896 363338 10376 363368
rect 13497 363338 13563 363341
rect 9896 363336 13563 363338
rect 9896 363280 13502 363336
rect 13558 363280 13563 363336
rect 9896 363278 13563 363280
rect 9896 363248 10376 363278
rect 13497 363275 13563 363278
rect 139629 357762 139695 357765
rect 233469 357762 233535 357765
rect 139629 357760 143050 357762
rect 139629 357704 139634 357760
rect 139690 357704 143050 357760
rect 139629 357702 143050 357704
rect 139629 357699 139695 357702
rect 80197 357626 80263 357629
rect 76382 357624 80263 357626
rect 76382 357568 80202 357624
rect 80258 357568 80263 357624
rect 76382 357566 80263 357568
rect 76382 357188 76442 357566
rect 80197 357563 80263 357566
rect 142990 357256 143050 357702
rect 233469 357760 237074 357762
rect 233469 357704 233474 357760
rect 233530 357704 237074 357760
rect 233469 357702 237074 357704
rect 233469 357699 233535 357702
rect 237014 357256 237074 357702
rect 328413 357490 328479 357493
rect 328413 357488 331098 357490
rect 328413 357432 328418 357488
rect 328474 357432 331098 357488
rect 328413 357430 331098 357432
rect 328413 357427 328479 357430
rect 331038 357256 331098 357430
rect 174037 357218 174103 357221
rect 267325 357218 267391 357221
rect 170804 357216 174103 357218
rect 170804 357160 174042 357216
rect 174098 357160 174103 357216
rect 170804 357158 174103 357160
rect 264828 357216 267391 357218
rect 264828 357160 267330 357216
rect 267386 357160 267391 357216
rect 264828 357158 267391 357160
rect 174037 357155 174103 357158
rect 267325 357155 267391 357158
rect 139629 356538 139695 356541
rect 233469 356538 233535 356541
rect 139629 356536 143050 356538
rect 139629 356480 139634 356536
rect 139690 356480 143050 356536
rect 139629 356478 143050 356480
rect 139629 356475 139695 356478
rect 80197 356402 80263 356405
rect 76382 356400 80263 356402
rect 76382 356344 80202 356400
rect 80258 356344 80263 356400
rect 76382 356342 80263 356344
rect 76382 356100 76442 356342
rect 80197 356339 80263 356342
rect 142990 356168 143050 356478
rect 233469 356536 237074 356538
rect 233469 356480 233474 356536
rect 233530 356480 237074 356536
rect 233469 356478 237074 356480
rect 233469 356475 233535 356478
rect 237014 356168 237074 356478
rect 173485 356130 173551 356133
rect 267877 356130 267943 356133
rect 170804 356128 173551 356130
rect 170804 356072 173490 356128
rect 173546 356072 173551 356128
rect 170804 356070 173551 356072
rect 264828 356128 267943 356130
rect 264828 356072 267882 356128
rect 267938 356072 267943 356128
rect 264828 356070 267943 356072
rect 173485 356067 173551 356070
rect 267877 356067 267943 356070
rect 328321 356130 328387 356133
rect 328321 356128 331068 356130
rect 328321 356072 328326 356128
rect 328382 356072 331068 356128
rect 328321 356070 331068 356072
rect 328321 356067 328387 356070
rect 139629 355178 139695 355181
rect 174037 355178 174103 355181
rect 139629 355176 143020 355178
rect 76198 355042 76258 355148
rect 139629 355120 139634 355176
rect 139690 355120 143020 355176
rect 139629 355118 143020 355120
rect 170804 355176 174103 355178
rect 170804 355120 174042 355176
rect 174098 355120 174103 355176
rect 170804 355118 174103 355120
rect 139629 355115 139695 355118
rect 174037 355115 174103 355118
rect 233469 355178 233535 355181
rect 267877 355178 267943 355181
rect 233469 355176 237044 355178
rect 233469 355120 233474 355176
rect 233530 355120 237044 355176
rect 233469 355118 237044 355120
rect 264828 355176 267943 355178
rect 264828 355120 267882 355176
rect 267938 355120 267943 355176
rect 264828 355118 267943 355120
rect 233469 355115 233535 355118
rect 267877 355115 267943 355118
rect 328413 355178 328479 355181
rect 328413 355176 331068 355178
rect 328413 355120 328418 355176
rect 328474 355120 331068 355176
rect 328413 355118 331068 355120
rect 328413 355115 328479 355118
rect 80197 355042 80263 355045
rect 76198 355040 80263 355042
rect 76198 354984 80202 355040
rect 80258 354984 80263 355040
rect 76198 354982 80263 354984
rect 80197 354979 80263 354982
rect 79277 354634 79343 354637
rect 76382 354632 79343 354634
rect 76382 354576 79282 354632
rect 79338 354576 79343 354632
rect 76382 354574 79343 354576
rect 76382 354060 76442 354574
rect 79277 354571 79343 354574
rect 139721 354634 139787 354637
rect 233561 354634 233627 354637
rect 328505 354634 328571 354637
rect 139721 354632 143050 354634
rect 139721 354576 139726 354632
rect 139782 354576 143050 354632
rect 139721 354574 143050 354576
rect 139721 354571 139787 354574
rect 142990 354128 143050 354574
rect 233561 354632 237074 354634
rect 233561 354576 233566 354632
rect 233622 354576 237074 354632
rect 233561 354574 237074 354576
rect 233561 354571 233627 354574
rect 237014 354128 237074 354574
rect 328505 354632 331098 354634
rect 328505 354576 328510 354632
rect 328566 354576 331098 354632
rect 328505 354574 331098 354576
rect 328505 354571 328571 354574
rect 331038 354128 331098 354574
rect 173761 354090 173827 354093
rect 267417 354090 267483 354093
rect 170804 354088 173827 354090
rect 170804 354032 173766 354088
rect 173822 354032 173827 354088
rect 170804 354030 173827 354032
rect 264828 354088 267483 354090
rect 264828 354032 267422 354088
rect 267478 354032 267483 354088
rect 264828 354030 267483 354032
rect 173761 354027 173827 354030
rect 267417 354027 267483 354030
rect 76057 353954 76123 353957
rect 76425 353954 76491 353957
rect 76057 353952 76491 353954
rect 76057 353896 76062 353952
rect 76118 353896 76430 353952
rect 76486 353896 76491 353952
rect 76057 353894 76491 353896
rect 76057 353891 76123 353894
rect 76425 353891 76491 353894
rect 139629 353546 139695 353549
rect 233469 353546 233535 353549
rect 139629 353544 143050 353546
rect 139629 353488 139634 353544
rect 139690 353488 143050 353544
rect 139629 353486 143050 353488
rect 139629 353483 139695 353486
rect 78909 353410 78975 353413
rect 76382 353408 78975 353410
rect 76382 353352 78914 353408
rect 78970 353352 78975 353408
rect 76382 353350 78975 353352
rect 76382 352972 76442 353350
rect 78909 353347 78975 353350
rect 142990 353040 143050 353486
rect 233469 353544 237074 353546
rect 233469 353488 233474 353544
rect 233530 353488 237074 353544
rect 233469 353486 237074 353488
rect 233469 353483 233535 353486
rect 237014 353040 237074 353486
rect 328045 353410 328111 353413
rect 328045 353408 331098 353410
rect 328045 353352 328050 353408
rect 328106 353352 331098 353408
rect 328045 353350 331098 353352
rect 328045 353347 328111 353350
rect 331038 353040 331098 353350
rect 174037 353002 174103 353005
rect 267877 353002 267943 353005
rect 170804 353000 174103 353002
rect 170804 352944 174042 353000
rect 174098 352944 174103 353000
rect 170804 352942 174103 352944
rect 264828 353000 267943 353002
rect 264828 352944 267882 353000
rect 267938 352944 267943 353000
rect 264828 352942 267943 352944
rect 174037 352939 174103 352942
rect 267877 352939 267943 352942
rect 430073 353002 430139 353005
rect 434416 353002 434896 353032
rect 430073 353000 434896 353002
rect 430073 352944 430078 353000
rect 430134 352944 434896 353000
rect 430073 352942 434896 352944
rect 430073 352939 430139 352942
rect 434416 352912 434896 352942
rect 139629 352322 139695 352325
rect 233469 352322 233535 352325
rect 328505 352322 328571 352325
rect 139629 352320 143050 352322
rect 139629 352264 139634 352320
rect 139690 352264 143050 352320
rect 139629 352262 143050 352264
rect 139629 352259 139695 352262
rect 80197 352186 80263 352189
rect 76382 352184 80263 352186
rect 76382 352128 80202 352184
rect 80258 352128 80263 352184
rect 76382 352126 80263 352128
rect 76382 352020 76442 352126
rect 80197 352123 80263 352126
rect 142990 352088 143050 352262
rect 233469 352320 237074 352322
rect 233469 352264 233474 352320
rect 233530 352264 237074 352320
rect 233469 352262 237074 352264
rect 233469 352259 233535 352262
rect 237014 352088 237074 352262
rect 328505 352320 331098 352322
rect 328505 352264 328510 352320
rect 328566 352264 331098 352320
rect 328505 352262 331098 352264
rect 328505 352259 328571 352262
rect 331038 352088 331098 352262
rect 97309 352052 97375 352053
rect 97309 352048 97356 352052
rect 97420 352050 97426 352052
rect 174037 352050 174103 352053
rect 267877 352050 267943 352053
rect 97309 351992 97314 352048
rect 97309 351988 97356 351992
rect 97420 351990 97466 352050
rect 170804 352048 174103 352050
rect 170804 351992 174042 352048
rect 174098 351992 174103 352048
rect 170804 351990 174103 351992
rect 264828 352048 267943 352050
rect 264828 351992 267882 352048
rect 267938 351992 267943 352048
rect 264828 351990 267943 351992
rect 97420 351988 97426 351990
rect 97309 351987 97375 351988
rect 174037 351987 174103 351990
rect 267877 351987 267943 351990
rect 180845 351642 180911 351645
rect 284989 351644 285055 351645
rect 180845 351640 184082 351642
rect 180845 351584 180850 351640
rect 180906 351584 184082 351640
rect 180845 351582 184082 351584
rect 180845 351579 180911 351582
rect 184022 351408 184082 351582
rect 284989 351640 285036 351644
rect 285100 351642 285106 351644
rect 284989 351584 284994 351640
rect 284989 351580 285036 351584
rect 285100 351582 285146 351642
rect 285100 351580 285106 351582
rect 284989 351579 285055 351580
rect 87189 351370 87255 351373
rect 131809 351370 131875 351373
rect 226293 351370 226359 351373
rect 87189 351368 90028 351370
rect 87189 351312 87194 351368
rect 87250 351312 90028 351368
rect 87189 351310 90028 351312
rect 129772 351368 131875 351370
rect 129772 351312 131814 351368
rect 131870 351312 131875 351368
rect 129772 351310 131875 351312
rect 223796 351368 226359 351370
rect 223796 351312 226298 351368
rect 226354 351312 226359 351368
rect 223796 351310 226359 351312
rect 87189 351307 87255 351310
rect 131809 351307 131875 351310
rect 226293 351307 226359 351310
rect 274777 351370 274843 351373
rect 320593 351370 320659 351373
rect 274777 351368 278076 351370
rect 274777 351312 274782 351368
rect 274838 351312 278076 351368
rect 274777 351310 278076 351312
rect 317820 351368 320659 351370
rect 317820 351312 320598 351368
rect 320654 351312 320659 351368
rect 317820 351310 320659 351312
rect 274777 351307 274843 351310
rect 320593 351307 320659 351310
rect 139721 350962 139787 350965
rect 174037 350962 174103 350965
rect 139721 350960 143020 350962
rect 76198 350690 76258 350932
rect 139721 350904 139726 350960
rect 139782 350904 143020 350960
rect 139721 350902 143020 350904
rect 170804 350960 174103 350962
rect 170804 350904 174042 350960
rect 174098 350904 174103 350960
rect 170804 350902 174103 350904
rect 139721 350899 139787 350902
rect 174037 350899 174103 350902
rect 233469 350962 233535 350965
rect 267693 350962 267759 350965
rect 233469 350960 237044 350962
rect 233469 350904 233474 350960
rect 233530 350904 237044 350960
rect 233469 350902 237044 350904
rect 264828 350960 267759 350962
rect 264828 350904 267698 350960
rect 267754 350904 267759 350960
rect 264828 350902 267759 350904
rect 233469 350899 233535 350902
rect 267693 350899 267759 350902
rect 327493 350962 327559 350965
rect 327493 350960 331068 350962
rect 327493 350904 327498 350960
rect 327554 350904 331068 350960
rect 327493 350902 331068 350904
rect 327493 350899 327559 350902
rect 80197 350690 80263 350693
rect 76198 350688 80263 350690
rect 76198 350632 80202 350688
rect 80258 350632 80263 350688
rect 76198 350630 80263 350632
rect 80197 350627 80263 350630
rect 139629 350554 139695 350557
rect 139629 350552 143050 350554
rect 139629 350496 139634 350552
rect 139690 350496 143050 350552
rect 139629 350494 143050 350496
rect 139629 350491 139695 350494
rect 79093 350418 79159 350421
rect 76382 350416 79159 350418
rect 76382 350360 79098 350416
rect 79154 350360 79159 350416
rect 76382 350358 79159 350360
rect 9896 350010 10376 350040
rect 13405 350010 13471 350013
rect 9896 350008 13471 350010
rect 9896 349952 13410 350008
rect 13466 349952 13471 350008
rect 9896 349950 13471 349952
rect 9896 349920 10376 349950
rect 13405 349947 13471 349950
rect 76382 349844 76442 350358
rect 79093 350355 79159 350358
rect 87465 350418 87531 350421
rect 131809 350418 131875 350421
rect 87465 350416 90028 350418
rect 87465 350360 87470 350416
rect 87526 350360 90028 350416
rect 87465 350358 90028 350360
rect 129772 350416 131875 350418
rect 129772 350360 131814 350416
rect 131870 350360 131875 350416
rect 129772 350358 131875 350360
rect 87465 350355 87531 350358
rect 131809 350355 131875 350358
rect 142990 349912 143050 350494
rect 226385 350418 226451 350421
rect 223796 350416 226451 350418
rect 180937 350010 181003 350013
rect 184022 350010 184082 350388
rect 223796 350360 226390 350416
rect 226446 350360 226451 350416
rect 223796 350358 226451 350360
rect 226385 350355 226451 350358
rect 233561 350418 233627 350421
rect 274961 350418 275027 350421
rect 321605 350418 321671 350421
rect 233561 350416 237074 350418
rect 233561 350360 233566 350416
rect 233622 350360 237074 350416
rect 233561 350358 237074 350360
rect 233561 350355 233627 350358
rect 180937 350008 184082 350010
rect 180937 349952 180942 350008
rect 180998 349952 184082 350008
rect 180937 349950 184082 349952
rect 180937 349947 181003 349950
rect 237014 349912 237074 350358
rect 274961 350416 278076 350418
rect 274961 350360 274966 350416
rect 275022 350360 278076 350416
rect 274961 350358 278076 350360
rect 317820 350416 321671 350418
rect 317820 350360 321610 350416
rect 321666 350360 321671 350416
rect 317820 350358 321671 350360
rect 274961 350355 275027 350358
rect 321605 350355 321671 350358
rect 327861 350418 327927 350421
rect 327861 350416 331098 350418
rect 327861 350360 327866 350416
rect 327922 350360 331098 350416
rect 327861 350358 331098 350360
rect 327861 350355 327927 350358
rect 331038 349912 331098 350358
rect 173761 349874 173827 349877
rect 267509 349874 267575 349877
rect 170804 349872 173827 349874
rect 170804 349816 173766 349872
rect 173822 349816 173827 349872
rect 170804 349814 173827 349816
rect 264828 349872 267575 349874
rect 264828 349816 267514 349872
rect 267570 349816 267575 349872
rect 264828 349814 267575 349816
rect 173761 349811 173827 349814
rect 267509 349811 267575 349814
rect 87281 349602 87347 349605
rect 131901 349602 131967 349605
rect 87281 349600 90028 349602
rect 87281 349544 87286 349600
rect 87342 349544 90028 349600
rect 87281 349542 90028 349544
rect 129772 349600 131967 349602
rect 129772 349544 131906 349600
rect 131962 349544 131967 349600
rect 129772 349542 131967 349544
rect 87281 349539 87347 349542
rect 131901 349539 131967 349542
rect 139629 349602 139695 349605
rect 182317 349602 182383 349605
rect 226477 349602 226543 349605
rect 139629 349600 143050 349602
rect 139629 349544 139634 349600
rect 139690 349544 143050 349600
rect 139629 349542 143050 349544
rect 139629 349539 139695 349542
rect 80197 349330 80263 349333
rect 76382 349328 80263 349330
rect 76382 349272 80202 349328
rect 80258 349272 80263 349328
rect 76382 349270 80263 349272
rect 76382 348892 76442 349270
rect 80197 349267 80263 349270
rect 142990 348960 143050 349542
rect 182317 349600 184052 349602
rect 182317 349544 182322 349600
rect 182378 349544 184052 349600
rect 182317 349542 184052 349544
rect 223796 349600 226543 349602
rect 223796 349544 226482 349600
rect 226538 349544 226543 349600
rect 223796 349542 226543 349544
rect 182317 349539 182383 349542
rect 226477 349539 226543 349542
rect 233469 349602 233535 349605
rect 274869 349602 274935 349605
rect 320685 349602 320751 349605
rect 233469 349600 237074 349602
rect 233469 349544 233474 349600
rect 233530 349544 237074 349600
rect 233469 349542 237074 349544
rect 233469 349539 233535 349542
rect 237014 348960 237074 349542
rect 274869 349600 278076 349602
rect 274869 349544 274874 349600
rect 274930 349544 278076 349600
rect 274869 349542 278076 349544
rect 317820 349600 320751 349602
rect 317820 349544 320690 349600
rect 320746 349544 320751 349600
rect 317820 349542 320751 349544
rect 274869 349539 274935 349542
rect 320685 349539 320751 349542
rect 327217 349602 327283 349605
rect 327217 349600 331098 349602
rect 327217 349544 327222 349600
rect 327278 349544 331098 349600
rect 327217 349542 331098 349544
rect 327217 349539 327283 349542
rect 331038 348960 331098 349542
rect 173025 348922 173091 348925
rect 267877 348922 267943 348925
rect 170804 348920 173091 348922
rect 170804 348864 173030 348920
rect 173086 348864 173091 348920
rect 170804 348862 173091 348864
rect 264828 348920 267943 348922
rect 264828 348864 267882 348920
rect 267938 348864 267943 348920
rect 264828 348862 267943 348864
rect 173025 348859 173091 348862
rect 267877 348859 267943 348862
rect 87373 348650 87439 348653
rect 131809 348650 131875 348653
rect 87373 348648 90028 348650
rect 87373 348592 87378 348648
rect 87434 348592 90028 348648
rect 87373 348590 90028 348592
rect 129772 348648 131875 348650
rect 129772 348592 131814 348648
rect 131870 348592 131875 348648
rect 129772 348590 131875 348592
rect 87373 348587 87439 348590
rect 131809 348587 131875 348590
rect 182133 348650 182199 348653
rect 226385 348650 226451 348653
rect 182133 348648 184052 348650
rect 182133 348592 182138 348648
rect 182194 348592 184052 348648
rect 182133 348590 184052 348592
rect 223796 348648 226451 348650
rect 223796 348592 226390 348648
rect 226446 348592 226451 348648
rect 223796 348590 226451 348592
rect 182133 348587 182199 348590
rect 226385 348587 226451 348590
rect 275053 348650 275119 348653
rect 321605 348650 321671 348653
rect 275053 348648 278076 348650
rect 275053 348592 275058 348648
rect 275114 348592 278076 348648
rect 275053 348590 278076 348592
rect 317820 348648 321671 348650
rect 317820 348592 321610 348648
rect 321666 348592 321671 348648
rect 317820 348590 321671 348592
rect 275053 348587 275119 348590
rect 321605 348587 321671 348590
rect 139629 348242 139695 348245
rect 233469 348242 233535 348245
rect 327125 348242 327191 348245
rect 139629 348240 143050 348242
rect 139629 348184 139634 348240
rect 139690 348184 143050 348240
rect 139629 348182 143050 348184
rect 139629 348179 139695 348182
rect 80197 348106 80263 348109
rect 76382 348104 80263 348106
rect 76382 348048 80202 348104
rect 80258 348048 80263 348104
rect 76382 348046 80263 348048
rect 76382 347804 76442 348046
rect 80197 348043 80263 348046
rect 142990 347872 143050 348182
rect 233469 348240 237074 348242
rect 233469 348184 233474 348240
rect 233530 348184 237074 348240
rect 233469 348182 237074 348184
rect 233469 348179 233535 348182
rect 237014 347872 237074 348182
rect 327125 348240 331098 348242
rect 327125 348184 327130 348240
rect 327186 348184 331098 348240
rect 327125 348182 331098 348184
rect 327125 348179 327191 348182
rect 331038 347872 331098 348182
rect 87097 347834 87163 347837
rect 132177 347834 132243 347837
rect 172933 347834 172999 347837
rect 226385 347834 226451 347837
rect 267877 347834 267943 347837
rect 87097 347832 90028 347834
rect 87097 347776 87102 347832
rect 87158 347776 90028 347832
rect 87097 347774 90028 347776
rect 129772 347832 132243 347834
rect 129772 347776 132182 347832
rect 132238 347776 132243 347832
rect 129772 347774 132243 347776
rect 170804 347832 172999 347834
rect 170804 347776 172938 347832
rect 172994 347776 172999 347832
rect 223796 347832 226451 347834
rect 170804 347774 172999 347776
rect 87097 347771 87163 347774
rect 132177 347771 132243 347774
rect 172933 347771 172999 347774
rect 180937 347290 181003 347293
rect 184022 347290 184082 347804
rect 223796 347776 226390 347832
rect 226446 347776 226451 347832
rect 223796 347774 226451 347776
rect 264828 347832 267943 347834
rect 264828 347776 267882 347832
rect 267938 347776 267943 347832
rect 264828 347774 267943 347776
rect 226385 347771 226451 347774
rect 267877 347771 267943 347774
rect 275145 347834 275211 347837
rect 321053 347834 321119 347837
rect 275145 347832 278076 347834
rect 275145 347776 275150 347832
rect 275206 347776 278076 347832
rect 275145 347774 278076 347776
rect 317820 347832 321119 347834
rect 317820 347776 321058 347832
rect 321114 347776 321119 347832
rect 317820 347774 321119 347776
rect 275145 347771 275211 347774
rect 321053 347771 321119 347774
rect 180937 347288 184082 347290
rect 180937 347232 180942 347288
rect 180998 347232 184082 347288
rect 180937 347230 184082 347232
rect 180937 347227 181003 347230
rect 87189 346882 87255 346885
rect 131901 346882 131967 346885
rect 87189 346880 90028 346882
rect 76198 346746 76258 346852
rect 87189 346824 87194 346880
rect 87250 346824 90028 346880
rect 87189 346822 90028 346824
rect 129772 346880 131967 346882
rect 129772 346824 131906 346880
rect 131962 346824 131967 346880
rect 129772 346822 131967 346824
rect 87189 346819 87255 346822
rect 131901 346819 131967 346822
rect 139629 346882 139695 346885
rect 174037 346882 174103 346885
rect 139629 346880 143020 346882
rect 139629 346824 139634 346880
rect 139690 346824 143020 346880
rect 139629 346822 143020 346824
rect 170804 346880 174103 346882
rect 170804 346824 174042 346880
rect 174098 346824 174103 346880
rect 170804 346822 174103 346824
rect 139629 346819 139695 346822
rect 174037 346819 174103 346822
rect 181581 346882 181647 346885
rect 226293 346882 226359 346885
rect 181581 346880 184052 346882
rect 181581 346824 181586 346880
rect 181642 346824 184052 346880
rect 181581 346822 184052 346824
rect 223796 346880 226359 346882
rect 223796 346824 226298 346880
rect 226354 346824 226359 346880
rect 223796 346822 226359 346824
rect 181581 346819 181647 346822
rect 226293 346819 226359 346822
rect 233377 346882 233443 346885
rect 267877 346882 267943 346885
rect 233377 346880 237044 346882
rect 233377 346824 233382 346880
rect 233438 346824 237044 346880
rect 233377 346822 237044 346824
rect 264828 346880 267943 346882
rect 264828 346824 267882 346880
rect 267938 346824 267943 346880
rect 264828 346822 267943 346824
rect 233377 346819 233443 346822
rect 267877 346819 267943 346822
rect 274961 346882 275027 346885
rect 320501 346882 320567 346885
rect 274961 346880 278076 346882
rect 274961 346824 274966 346880
rect 275022 346824 278076 346880
rect 274961 346822 278076 346824
rect 317820 346880 320567 346882
rect 317820 346824 320506 346880
rect 320562 346824 320567 346880
rect 317820 346822 320567 346824
rect 274961 346819 275027 346822
rect 320501 346819 320567 346822
rect 327217 346882 327283 346885
rect 327217 346880 331068 346882
rect 327217 346824 327222 346880
rect 327278 346824 331068 346880
rect 327217 346822 331068 346824
rect 327217 346819 327283 346822
rect 80197 346746 80263 346749
rect 76198 346744 80263 346746
rect 76198 346688 80202 346744
rect 80258 346688 80263 346744
rect 76198 346686 80263 346688
rect 80197 346683 80263 346686
rect 233285 346474 233351 346477
rect 327033 346474 327099 346477
rect 233285 346472 237074 346474
rect 233285 346416 233290 346472
rect 233346 346416 237074 346472
rect 233285 346414 237074 346416
rect 233285 346411 233351 346414
rect 79277 346338 79343 346341
rect 76382 346336 79343 346338
rect 76382 346280 79282 346336
rect 79338 346280 79343 346336
rect 76382 346278 79343 346280
rect 76382 345764 76442 346278
rect 79277 346275 79343 346278
rect 139721 346338 139787 346341
rect 139721 346336 143050 346338
rect 139721 346280 139726 346336
rect 139782 346280 143050 346336
rect 139721 346278 143050 346280
rect 139721 346275 139787 346278
rect 88109 346066 88175 346069
rect 131809 346066 131875 346069
rect 88109 346064 90028 346066
rect 88109 346008 88114 346064
rect 88170 346008 90028 346064
rect 88109 346006 90028 346008
rect 129772 346064 131875 346066
rect 129772 346008 131814 346064
rect 131870 346008 131875 346064
rect 129772 346006 131875 346008
rect 88109 346003 88175 346006
rect 131809 346003 131875 346006
rect 142990 345832 143050 346278
rect 182317 346066 182383 346069
rect 226385 346066 226451 346069
rect 182317 346064 184052 346066
rect 182317 346008 182322 346064
rect 182378 346008 184052 346064
rect 182317 346006 184052 346008
rect 223796 346064 226451 346066
rect 223796 346008 226390 346064
rect 226446 346008 226451 346064
rect 223796 346006 226451 346008
rect 182317 346003 182383 346006
rect 226385 346003 226451 346006
rect 237014 345832 237074 346414
rect 327033 346472 331098 346474
rect 327033 346416 327038 346472
rect 327094 346416 331098 346472
rect 327033 346414 331098 346416
rect 327033 346411 327099 346414
rect 274869 346066 274935 346069
rect 321605 346066 321671 346069
rect 274869 346064 278076 346066
rect 274869 346008 274874 346064
rect 274930 346008 278076 346064
rect 274869 346006 278076 346008
rect 317820 346064 321671 346066
rect 317820 346008 321610 346064
rect 321666 346008 321671 346064
rect 317820 346006 321671 346008
rect 274869 346003 274935 346006
rect 321605 346003 321671 346006
rect 331038 345832 331098 346414
rect 173761 345794 173827 345797
rect 267417 345794 267483 345797
rect 170804 345792 173827 345794
rect 170804 345736 173766 345792
rect 173822 345736 173827 345792
rect 170804 345734 173827 345736
rect 264828 345792 267483 345794
rect 264828 345736 267422 345792
rect 267478 345736 267483 345792
rect 264828 345734 267483 345736
rect 173761 345731 173827 345734
rect 267417 345731 267483 345734
rect 139813 345386 139879 345389
rect 139813 345384 143050 345386
rect 139813 345328 139818 345384
rect 139874 345328 143050 345384
rect 139813 345326 143050 345328
rect 139813 345323 139879 345326
rect 87373 345114 87439 345117
rect 132361 345114 132427 345117
rect 87373 345112 90028 345114
rect 87373 345056 87378 345112
rect 87434 345056 90028 345112
rect 87373 345054 90028 345056
rect 129772 345112 132427 345114
rect 129772 345056 132366 345112
rect 132422 345056 132427 345112
rect 129772 345054 132427 345056
rect 87373 345051 87439 345054
rect 132361 345051 132427 345054
rect 80197 344842 80263 344845
rect 76382 344840 80263 344842
rect 76382 344784 80202 344840
rect 80258 344784 80263 344840
rect 76382 344782 80263 344784
rect 76382 344676 76442 344782
rect 80197 344779 80263 344782
rect 142990 344744 143050 345326
rect 233469 345250 233535 345253
rect 233469 345248 237074 345250
rect 233469 345192 233474 345248
rect 233530 345192 237074 345248
rect 233469 345190 237074 345192
rect 233469 345187 233535 345190
rect 226477 345114 226543 345117
rect 223796 345112 226543 345114
rect 172749 344706 172815 344709
rect 170804 344704 172815 344706
rect 170804 344648 172754 344704
rect 172810 344648 172815 344704
rect 170804 344646 172815 344648
rect 172749 344643 172815 344646
rect 180937 344706 181003 344709
rect 184022 344706 184082 345084
rect 223796 345056 226482 345112
rect 226538 345056 226543 345112
rect 223796 345054 226543 345056
rect 226477 345051 226543 345054
rect 237014 344744 237074 345190
rect 274869 345114 274935 345117
rect 320961 345114 321027 345117
rect 274869 345112 278076 345114
rect 274869 345056 274874 345112
rect 274930 345056 278076 345112
rect 274869 345054 278076 345056
rect 317820 345112 321027 345114
rect 317820 345056 320966 345112
rect 321022 345056 321027 345112
rect 317820 345054 321027 345056
rect 274869 345051 274935 345054
rect 320961 345051 321027 345054
rect 328045 345114 328111 345117
rect 328045 345112 331098 345114
rect 328045 345056 328050 345112
rect 328106 345056 331098 345112
rect 328045 345054 331098 345056
rect 328045 345051 328111 345054
rect 331038 344744 331098 345054
rect 267877 344706 267943 344709
rect 180937 344704 184082 344706
rect 180937 344648 180942 344704
rect 180998 344648 184082 344704
rect 180937 344646 184082 344648
rect 264828 344704 267943 344706
rect 264828 344648 267882 344704
rect 267938 344648 267943 344704
rect 264828 344646 267943 344648
rect 180937 344643 181003 344646
rect 267877 344643 267943 344646
rect 88477 344298 88543 344301
rect 131809 344298 131875 344301
rect 88477 344296 90028 344298
rect 88477 344240 88482 344296
rect 88538 344240 90028 344296
rect 88477 344238 90028 344240
rect 129772 344296 131875 344298
rect 129772 344240 131814 344296
rect 131870 344240 131875 344296
rect 129772 344238 131875 344240
rect 88477 344235 88543 344238
rect 131809 344235 131875 344238
rect 182317 344298 182383 344301
rect 226385 344298 226451 344301
rect 182317 344296 184052 344298
rect 182317 344240 182322 344296
rect 182378 344240 184052 344296
rect 182317 344238 184052 344240
rect 223796 344296 226451 344298
rect 223796 344240 226390 344296
rect 226446 344240 226451 344296
rect 223796 344238 226451 344240
rect 182317 344235 182383 344238
rect 226385 344235 226451 344238
rect 275053 344298 275119 344301
rect 321605 344298 321671 344301
rect 275053 344296 278076 344298
rect 275053 344240 275058 344296
rect 275114 344240 278076 344296
rect 275053 344238 278076 344240
rect 317820 344296 321671 344298
rect 317820 344240 321610 344296
rect 321666 344240 321671 344296
rect 317820 344238 321671 344240
rect 275053 344235 275119 344238
rect 321605 344235 321671 344238
rect 139629 344162 139695 344165
rect 266957 344162 267023 344165
rect 267141 344162 267207 344165
rect 139629 344160 143050 344162
rect 139629 344104 139634 344160
rect 139690 344104 143050 344160
rect 139629 344102 143050 344104
rect 139629 344099 139695 344102
rect 79645 344026 79711 344029
rect 76382 344024 79711 344026
rect 76382 343968 79650 344024
rect 79706 343968 79711 344024
rect 76382 343966 79711 343968
rect 76382 343724 76442 343966
rect 79645 343963 79711 343966
rect 142990 343792 143050 344102
rect 266957 344160 267207 344162
rect 266957 344104 266962 344160
rect 267018 344104 267146 344160
rect 267202 344104 267207 344160
rect 266957 344102 267207 344104
rect 266957 344099 267023 344102
rect 267141 344099 267207 344102
rect 233469 344026 233535 344029
rect 328505 344026 328571 344029
rect 233469 344024 237074 344026
rect 233469 343968 233474 344024
rect 233530 343968 237074 344024
rect 233469 343966 237074 343968
rect 233469 343963 233535 343966
rect 237014 343792 237074 343966
rect 328505 344024 331098 344026
rect 328505 343968 328510 344024
rect 328566 343968 331098 344024
rect 328505 343966 331098 343968
rect 328505 343963 328571 343966
rect 331038 343792 331098 343966
rect 172841 343754 172907 343757
rect 266681 343754 266747 343757
rect 170804 343752 172907 343754
rect 170804 343696 172846 343752
rect 172902 343696 172907 343752
rect 170804 343694 172907 343696
rect 264828 343752 266747 343754
rect 264828 343696 266686 343752
rect 266742 343696 266747 343752
rect 264828 343694 266747 343696
rect 172841 343691 172907 343694
rect 266681 343691 266747 343694
rect 87281 343346 87347 343349
rect 131809 343346 131875 343349
rect 87281 343344 90028 343346
rect 87281 343288 87286 343344
rect 87342 343288 90028 343344
rect 87281 343286 90028 343288
rect 129772 343344 131875 343346
rect 129772 343288 131814 343344
rect 131870 343288 131875 343344
rect 129772 343286 131875 343288
rect 87281 343283 87347 343286
rect 131809 343283 131875 343286
rect 181397 343346 181463 343349
rect 226385 343346 226451 343349
rect 181397 343344 184052 343346
rect 181397 343288 181402 343344
rect 181458 343288 184052 343344
rect 181397 343286 184052 343288
rect 223796 343344 226451 343346
rect 223796 343288 226390 343344
rect 226446 343288 226451 343344
rect 223796 343286 226451 343288
rect 181397 343283 181463 343286
rect 226385 343283 226451 343286
rect 275145 343346 275211 343349
rect 321605 343346 321671 343349
rect 275145 343344 278076 343346
rect 275145 343288 275150 343344
rect 275206 343288 278076 343344
rect 275145 343286 278076 343288
rect 317820 343344 321671 343346
rect 317820 343288 321610 343344
rect 321666 343288 321671 343344
rect 317820 343286 321671 343288
rect 275145 343283 275211 343286
rect 321605 343283 321671 343286
rect 80197 342802 80263 342805
rect 76382 342800 80263 342802
rect 76382 342744 80202 342800
rect 80258 342744 80263 342800
rect 76382 342742 80263 342744
rect 76382 342636 76442 342742
rect 80197 342739 80263 342742
rect 139629 342666 139695 342669
rect 172933 342666 172999 342669
rect 139629 342664 143020 342666
rect 139629 342608 139634 342664
rect 139690 342608 143020 342664
rect 139629 342606 143020 342608
rect 170804 342664 172999 342666
rect 170804 342608 172938 342664
rect 172994 342608 172999 342664
rect 170804 342606 172999 342608
rect 139629 342603 139695 342606
rect 172933 342603 172999 342606
rect 234573 342666 234639 342669
rect 267877 342666 267943 342669
rect 234573 342664 237044 342666
rect 234573 342608 234578 342664
rect 234634 342608 237044 342664
rect 234573 342606 237044 342608
rect 264828 342664 267943 342666
rect 264828 342608 267882 342664
rect 267938 342608 267943 342664
rect 264828 342606 267943 342608
rect 234573 342603 234639 342606
rect 267877 342603 267943 342606
rect 326941 342666 327007 342669
rect 326941 342664 331068 342666
rect 326941 342608 326946 342664
rect 327002 342608 331068 342664
rect 326941 342606 331068 342608
rect 326941 342603 327007 342606
rect 87557 342394 87623 342397
rect 131901 342394 131967 342397
rect 87557 342392 90028 342394
rect 87557 342336 87562 342392
rect 87618 342336 90028 342392
rect 87557 342334 90028 342336
rect 129772 342392 131967 342394
rect 129772 342336 131906 342392
rect 131962 342336 131967 342392
rect 129772 342334 131967 342336
rect 87557 342331 87623 342334
rect 131901 342331 131967 342334
rect 181397 342394 181463 342397
rect 226477 342394 226543 342397
rect 181397 342392 184052 342394
rect 181397 342336 181402 342392
rect 181458 342336 184052 342392
rect 181397 342334 184052 342336
rect 223796 342392 226543 342394
rect 223796 342336 226482 342392
rect 226538 342336 226543 342392
rect 223796 342334 226543 342336
rect 181397 342331 181463 342334
rect 226477 342331 226543 342334
rect 275237 342394 275303 342397
rect 321053 342394 321119 342397
rect 275237 342392 278076 342394
rect 275237 342336 275242 342392
rect 275298 342336 278076 342392
rect 275237 342334 278076 342336
rect 317820 342392 321119 342394
rect 317820 342336 321058 342392
rect 321114 342336 321119 342392
rect 317820 342334 321119 342336
rect 275237 342331 275303 342334
rect 321053 342331 321119 342334
rect 139721 342258 139787 342261
rect 234481 342258 234547 342261
rect 139721 342256 143050 342258
rect 139721 342200 139726 342256
rect 139782 342200 143050 342256
rect 139721 342198 143050 342200
rect 139721 342195 139787 342198
rect 80197 341850 80263 341853
rect 76382 341848 80263 341850
rect 76382 341792 80202 341848
rect 80258 341792 80263 341848
rect 76382 341790 80263 341792
rect 76382 341548 76442 341790
rect 80197 341787 80263 341790
rect 142990 341616 143050 342198
rect 234481 342256 237074 342258
rect 234481 342200 234486 342256
rect 234542 342200 237074 342256
rect 234481 342198 237074 342200
rect 234481 342195 234547 342198
rect 237014 341616 237074 342198
rect 328045 342122 328111 342125
rect 328045 342120 331098 342122
rect 328045 342064 328050 342120
rect 328106 342064 331098 342120
rect 328045 342062 331098 342064
rect 328045 342059 328111 342062
rect 331038 341616 331098 342062
rect 87189 341578 87255 341581
rect 131809 341578 131875 341581
rect 172749 341578 172815 341581
rect 87189 341576 90028 341578
rect 87189 341520 87194 341576
rect 87250 341520 90028 341576
rect 87189 341518 90028 341520
rect 129772 341576 131875 341578
rect 129772 341520 131814 341576
rect 131870 341520 131875 341576
rect 129772 341518 131875 341520
rect 170804 341576 172815 341578
rect 170804 341520 172754 341576
rect 172810 341520 172815 341576
rect 170804 341518 172815 341520
rect 87189 341515 87255 341518
rect 131809 341515 131875 341518
rect 172749 341515 172815 341518
rect 182317 341578 182383 341581
rect 226385 341578 226451 341581
rect 267601 341578 267667 341581
rect 182317 341576 184052 341578
rect 182317 341520 182322 341576
rect 182378 341520 184052 341576
rect 182317 341518 184052 341520
rect 223796 341576 226451 341578
rect 223796 341520 226390 341576
rect 226446 341520 226451 341576
rect 223796 341518 226451 341520
rect 264828 341576 267667 341578
rect 264828 341520 267606 341576
rect 267662 341520 267667 341576
rect 264828 341518 267667 341520
rect 182317 341515 182383 341518
rect 226385 341515 226451 341518
rect 267601 341515 267667 341518
rect 274961 341578 275027 341581
rect 321605 341578 321671 341581
rect 274961 341576 278076 341578
rect 274961 341520 274966 341576
rect 275022 341520 278076 341576
rect 274961 341518 278076 341520
rect 317820 341576 321671 341578
rect 317820 341520 321610 341576
rect 321666 341520 321671 341576
rect 317820 341518 321671 341520
rect 274961 341515 275027 341518
rect 321605 341515 321671 341518
rect 139813 341306 139879 341309
rect 234389 341306 234455 341309
rect 327401 341306 327467 341309
rect 139813 341304 143050 341306
rect 139813 341248 139818 341304
rect 139874 341248 143050 341304
rect 139813 341246 143050 341248
rect 139813 341243 139879 341246
rect 80197 341034 80263 341037
rect 76382 341032 80263 341034
rect 76382 340976 80202 341032
rect 80258 340976 80263 341032
rect 76382 340974 80263 340976
rect 76382 340596 76442 340974
rect 80197 340971 80263 340974
rect 142990 340664 143050 341246
rect 234389 341304 237074 341306
rect 234389 341248 234394 341304
rect 234450 341248 237074 341304
rect 234389 341246 237074 341248
rect 234389 341243 234455 341246
rect 237014 340664 237074 341246
rect 327401 341304 331098 341306
rect 327401 341248 327406 341304
rect 327462 341248 331098 341304
rect 327401 341246 331098 341248
rect 327401 341243 327467 341246
rect 331038 340664 331098 341246
rect 87373 340626 87439 340629
rect 131809 340626 131875 340629
rect 173117 340626 173183 340629
rect 87373 340624 90028 340626
rect 87373 340568 87378 340624
rect 87434 340568 90028 340624
rect 87373 340566 90028 340568
rect 129772 340624 131875 340626
rect 129772 340568 131814 340624
rect 131870 340568 131875 340624
rect 129772 340566 131875 340568
rect 170804 340624 173183 340626
rect 170804 340568 173122 340624
rect 173178 340568 173183 340624
rect 170804 340566 173183 340568
rect 87373 340563 87439 340566
rect 131809 340563 131875 340566
rect 173117 340563 173183 340566
rect 181397 340626 181463 340629
rect 226385 340626 226451 340629
rect 267877 340626 267943 340629
rect 181397 340624 184052 340626
rect 181397 340568 181402 340624
rect 181458 340568 184052 340624
rect 181397 340566 184052 340568
rect 223796 340624 226451 340626
rect 223796 340568 226390 340624
rect 226446 340568 226451 340624
rect 223796 340566 226451 340568
rect 264828 340624 267943 340626
rect 264828 340568 267882 340624
rect 267938 340568 267943 340624
rect 264828 340566 267943 340568
rect 181397 340563 181463 340566
rect 226385 340563 226451 340566
rect 267877 340563 267943 340566
rect 274869 340626 274935 340629
rect 320593 340626 320659 340629
rect 274869 340624 278076 340626
rect 274869 340568 274874 340624
rect 274930 340568 278076 340624
rect 274869 340566 278076 340568
rect 317820 340624 320659 340626
rect 317820 340568 320598 340624
rect 320654 340568 320659 340624
rect 317820 340566 320659 340568
rect 274869 340563 274935 340566
rect 320593 340563 320659 340566
rect 429429 340490 429495 340493
rect 434416 340490 434896 340520
rect 429429 340488 434896 340490
rect 429429 340432 429434 340488
rect 429490 340432 434896 340488
rect 429429 340430 434896 340432
rect 429429 340427 429495 340430
rect 434416 340400 434896 340430
rect 139629 339946 139695 339949
rect 233469 339946 233535 339949
rect 327217 339946 327283 339949
rect 139629 339944 143050 339946
rect 139629 339888 139634 339944
rect 139690 339888 143050 339944
rect 139629 339886 143050 339888
rect 139629 339883 139695 339886
rect 80197 339810 80263 339813
rect 76382 339808 80263 339810
rect 76382 339752 80202 339808
rect 80258 339752 80263 339808
rect 76382 339750 80263 339752
rect 76382 339508 76442 339750
rect 80197 339747 80263 339750
rect 87281 339810 87347 339813
rect 131901 339810 131967 339813
rect 87281 339808 90028 339810
rect 87281 339752 87286 339808
rect 87342 339752 90028 339808
rect 87281 339750 90028 339752
rect 129772 339808 131967 339810
rect 129772 339752 131906 339808
rect 131962 339752 131967 339808
rect 129772 339750 131967 339752
rect 87281 339747 87347 339750
rect 131901 339747 131967 339750
rect 142990 339576 143050 339886
rect 233469 339944 237074 339946
rect 233469 339888 233474 339944
rect 233530 339888 237074 339944
rect 233469 339886 237074 339888
rect 233469 339883 233535 339886
rect 181581 339810 181647 339813
rect 226477 339810 226543 339813
rect 181581 339808 184052 339810
rect 181581 339752 181586 339808
rect 181642 339752 184052 339808
rect 181581 339750 184052 339752
rect 223796 339808 226543 339810
rect 223796 339752 226482 339808
rect 226538 339752 226543 339808
rect 223796 339750 226543 339752
rect 181581 339747 181647 339750
rect 226477 339747 226543 339750
rect 237014 339576 237074 339886
rect 327217 339944 331098 339946
rect 327217 339888 327222 339944
rect 327278 339888 331098 339944
rect 327217 339886 331098 339888
rect 327217 339883 327283 339886
rect 275053 339810 275119 339813
rect 320501 339810 320567 339813
rect 275053 339808 278076 339810
rect 275053 339752 275058 339808
rect 275114 339752 278076 339808
rect 275053 339750 278076 339752
rect 317820 339808 320567 339810
rect 317820 339752 320506 339808
rect 320562 339752 320567 339808
rect 317820 339750 320567 339752
rect 275053 339747 275119 339750
rect 320501 339747 320567 339750
rect 331038 339576 331098 339886
rect 173945 339538 174011 339541
rect 267877 339538 267943 339541
rect 170804 339536 174011 339538
rect 170804 339480 173950 339536
rect 174006 339480 174011 339536
rect 170804 339478 174011 339480
rect 264828 339536 267943 339538
rect 264828 339480 267882 339536
rect 267938 339480 267943 339536
rect 264828 339478 267943 339480
rect 173945 339475 174011 339478
rect 267877 339475 267943 339478
rect 180293 339402 180359 339405
rect 180293 339400 184082 339402
rect 180293 339344 180298 339400
rect 180354 339344 184082 339400
rect 180293 339342 184082 339344
rect 180293 339339 180359 339342
rect 184022 338896 184082 339342
rect 87465 338858 87531 338861
rect 131809 338858 131875 338861
rect 226385 338858 226451 338861
rect 87465 338856 90028 338858
rect 87465 338800 87470 338856
rect 87526 338800 90028 338856
rect 87465 338798 90028 338800
rect 129772 338856 131875 338858
rect 129772 338800 131814 338856
rect 131870 338800 131875 338856
rect 129772 338798 131875 338800
rect 223796 338856 226451 338858
rect 223796 338800 226390 338856
rect 226446 338800 226451 338856
rect 223796 338798 226451 338800
rect 87465 338795 87531 338798
rect 131809 338795 131875 338798
rect 226385 338795 226451 338798
rect 274869 338858 274935 338861
rect 320409 338858 320475 338861
rect 274869 338856 278076 338858
rect 274869 338800 274874 338856
rect 274930 338800 278076 338856
rect 274869 338798 278076 338800
rect 317820 338856 320475 338858
rect 317820 338800 320414 338856
rect 320470 338800 320475 338856
rect 317820 338798 320475 338800
rect 274869 338795 274935 338798
rect 320409 338795 320475 338798
rect 139721 338586 139787 338589
rect 174037 338586 174103 338589
rect 139721 338584 143020 338586
rect 76198 338450 76258 338556
rect 139721 338528 139726 338584
rect 139782 338528 143020 338584
rect 139721 338526 143020 338528
rect 170804 338584 174103 338586
rect 170804 338528 174042 338584
rect 174098 338528 174103 338584
rect 170804 338526 174103 338528
rect 139721 338523 139787 338526
rect 174037 338523 174103 338526
rect 233469 338586 233535 338589
rect 267877 338586 267943 338589
rect 233469 338584 237044 338586
rect 233469 338528 233474 338584
rect 233530 338528 237044 338584
rect 233469 338526 237044 338528
rect 264828 338584 267943 338586
rect 264828 338528 267882 338584
rect 267938 338528 267943 338584
rect 264828 338526 267943 338528
rect 233469 338523 233535 338526
rect 267877 338523 267943 338526
rect 327125 338586 327191 338589
rect 327125 338584 331068 338586
rect 327125 338528 327130 338584
rect 327186 338528 331068 338584
rect 327125 338526 331068 338528
rect 327125 338523 327191 338526
rect 80197 338450 80263 338453
rect 76198 338448 80263 338450
rect 76198 338392 80202 338448
rect 80258 338392 80263 338448
rect 76198 338390 80263 338392
rect 80197 338387 80263 338390
rect 233653 338178 233719 338181
rect 327033 338178 327099 338181
rect 233653 338176 237074 338178
rect 233653 338120 233658 338176
rect 233714 338120 237074 338176
rect 233653 338118 237074 338120
rect 233653 338115 233719 338118
rect 80105 338042 80171 338045
rect 76382 338040 80171 338042
rect 76382 337984 80110 338040
rect 80166 337984 80171 338040
rect 76382 337982 80171 337984
rect 76382 337468 76442 337982
rect 80105 337979 80171 337982
rect 87189 338042 87255 338045
rect 131809 338042 131875 338045
rect 87189 338040 90028 338042
rect 87189 337984 87194 338040
rect 87250 337984 90028 338040
rect 87189 337982 90028 337984
rect 129772 338040 131875 338042
rect 129772 337984 131814 338040
rect 131870 337984 131875 338040
rect 129772 337982 131875 337984
rect 87189 337979 87255 337982
rect 131809 337979 131875 337982
rect 139813 338042 139879 338045
rect 181765 338042 181831 338045
rect 226385 338042 226451 338045
rect 139813 338040 143050 338042
rect 139813 337984 139818 338040
rect 139874 337984 143050 338040
rect 139813 337982 143050 337984
rect 139813 337979 139879 337982
rect 142990 337536 143050 337982
rect 181765 338040 184052 338042
rect 181765 337984 181770 338040
rect 181826 337984 184052 338040
rect 181765 337982 184052 337984
rect 223796 338040 226451 338042
rect 223796 337984 226390 338040
rect 226446 337984 226451 338040
rect 223796 337982 226451 337984
rect 181765 337979 181831 337982
rect 226385 337979 226451 337982
rect 237014 337536 237074 338118
rect 327033 338176 331098 338178
rect 327033 338120 327038 338176
rect 327094 338120 331098 338176
rect 327033 338118 331098 338120
rect 327033 338115 327099 338118
rect 274869 338042 274935 338045
rect 320409 338042 320475 338045
rect 274869 338040 278076 338042
rect 274869 337984 274874 338040
rect 274930 337984 278076 338040
rect 274869 337982 278076 337984
rect 317820 338040 320475 338042
rect 317820 337984 320414 338040
rect 320470 337984 320475 338040
rect 317820 337982 320475 337984
rect 274869 337979 274935 337982
rect 320409 337979 320475 337982
rect 331038 337536 331098 338118
rect 173761 337498 173827 337501
rect 267509 337498 267575 337501
rect 170804 337496 173827 337498
rect 170804 337440 173766 337496
rect 173822 337440 173827 337496
rect 170804 337438 173827 337440
rect 264828 337496 267575 337498
rect 264828 337440 267514 337496
rect 267570 337440 267575 337496
rect 264828 337438 267575 337440
rect 173761 337435 173827 337438
rect 267509 337435 267575 337438
rect 87557 337090 87623 337093
rect 131901 337090 131967 337093
rect 87557 337088 90028 337090
rect 87557 337032 87562 337088
rect 87618 337032 90028 337088
rect 87557 337030 90028 337032
rect 129772 337088 131967 337090
rect 129772 337032 131906 337088
rect 131962 337032 131967 337088
rect 129772 337030 131967 337032
rect 87557 337027 87623 337030
rect 131901 337027 131967 337030
rect 181581 337090 181647 337093
rect 226385 337090 226451 337093
rect 181581 337088 184052 337090
rect 181581 337032 181586 337088
rect 181642 337032 184052 337088
rect 181581 337030 184052 337032
rect 223796 337088 226451 337090
rect 223796 337032 226390 337088
rect 226446 337032 226451 337088
rect 223796 337030 226451 337032
rect 181581 337027 181647 337030
rect 226385 337027 226451 337030
rect 233561 337090 233627 337093
rect 274961 337090 275027 337093
rect 320409 337090 320475 337093
rect 233561 337088 237074 337090
rect 233561 337032 233566 337088
rect 233622 337032 237074 337088
rect 233561 337030 237074 337032
rect 233561 337027 233627 337030
rect 79829 336818 79895 336821
rect 76382 336816 79895 336818
rect 76382 336760 79834 336816
rect 79890 336760 79895 336816
rect 76382 336758 79895 336760
rect 9896 336682 10376 336712
rect 13405 336682 13471 336685
rect 9896 336680 13471 336682
rect 9896 336624 13410 336680
rect 13466 336624 13471 336680
rect 9896 336622 13471 336624
rect 9896 336592 10376 336622
rect 13405 336619 13471 336622
rect 76382 336380 76442 336758
rect 79829 336755 79895 336758
rect 139537 336818 139603 336821
rect 139537 336816 143050 336818
rect 139537 336760 139542 336816
rect 139598 336760 143050 336816
rect 139537 336758 143050 336760
rect 139537 336755 139603 336758
rect 142990 336448 143050 336758
rect 237014 336448 237074 337030
rect 274961 337088 278076 337090
rect 274961 337032 274966 337088
rect 275022 337032 278076 337088
rect 274961 337030 278076 337032
rect 317820 337088 320475 337090
rect 317820 337032 320414 337088
rect 320470 337032 320475 337088
rect 317820 337030 320475 337032
rect 274961 337027 275027 337030
rect 320409 337027 320475 337030
rect 327861 337090 327927 337093
rect 327861 337088 331098 337090
rect 327861 337032 327866 337088
rect 327922 337032 331098 337088
rect 327861 337030 331098 337032
rect 327861 337027 327927 337030
rect 331038 336448 331098 337030
rect 173853 336410 173919 336413
rect 267325 336410 267391 336413
rect 170804 336408 173919 336410
rect 170804 336352 173858 336408
rect 173914 336352 173919 336408
rect 170804 336350 173919 336352
rect 264828 336408 267391 336410
rect 264828 336352 267330 336408
rect 267386 336352 267391 336408
rect 264828 336350 267391 336352
rect 173853 336347 173919 336350
rect 267325 336347 267391 336350
rect 87189 336274 87255 336277
rect 131809 336274 131875 336277
rect 87189 336272 90028 336274
rect 87189 336216 87194 336272
rect 87250 336216 90028 336272
rect 87189 336214 90028 336216
rect 129772 336272 131875 336274
rect 129772 336216 131814 336272
rect 131870 336216 131875 336272
rect 129772 336214 131875 336216
rect 87189 336211 87255 336214
rect 131809 336211 131875 336214
rect 181765 336274 181831 336277
rect 226569 336274 226635 336277
rect 181765 336272 184052 336274
rect 181765 336216 181770 336272
rect 181826 336216 184052 336272
rect 181765 336214 184052 336216
rect 223796 336272 226635 336274
rect 223796 336216 226574 336272
rect 226630 336216 226635 336272
rect 223796 336214 226635 336216
rect 181765 336211 181831 336214
rect 226569 336211 226635 336214
rect 274869 336274 274935 336277
rect 320501 336274 320567 336277
rect 274869 336272 278076 336274
rect 274869 336216 274874 336272
rect 274930 336216 278076 336272
rect 274869 336214 278076 336216
rect 317820 336272 320567 336274
rect 317820 336216 320506 336272
rect 320562 336216 320567 336272
rect 317820 336214 320567 336216
rect 274869 336211 274935 336214
rect 320501 336211 320567 336214
rect 139629 335866 139695 335869
rect 233469 335866 233535 335869
rect 327217 335866 327283 335869
rect 139629 335864 143050 335866
rect 139629 335808 139634 335864
rect 139690 335808 143050 335864
rect 139629 335806 143050 335808
rect 139629 335803 139695 335806
rect 80197 335730 80263 335733
rect 76382 335728 80263 335730
rect 76382 335672 80202 335728
rect 80258 335672 80263 335728
rect 76382 335670 80263 335672
rect 76382 335428 76442 335670
rect 80197 335667 80263 335670
rect 142990 335496 143050 335806
rect 233469 335864 237074 335866
rect 233469 335808 233474 335864
rect 233530 335808 237074 335864
rect 233469 335806 237074 335808
rect 233469 335803 233535 335806
rect 237014 335496 237074 335806
rect 327217 335864 331098 335866
rect 327217 335808 327222 335864
rect 327278 335808 331098 335864
rect 327217 335806 331098 335808
rect 327217 335803 327283 335806
rect 331038 335496 331098 335806
rect 173485 335458 173551 335461
rect 267877 335458 267943 335461
rect 170804 335456 173551 335458
rect 170804 335400 173490 335456
rect 173546 335400 173551 335456
rect 170804 335398 173551 335400
rect 264828 335456 267943 335458
rect 264828 335400 267882 335456
rect 267938 335400 267943 335456
rect 264828 335398 267943 335400
rect 173485 335395 173551 335398
rect 267877 335395 267943 335398
rect 139629 334370 139695 334373
rect 174037 334370 174103 334373
rect 139629 334368 143020 334370
rect 76198 334098 76258 334340
rect 139629 334312 139634 334368
rect 139690 334312 143020 334368
rect 139629 334310 143020 334312
rect 170804 334368 174103 334370
rect 170804 334312 174042 334368
rect 174098 334312 174103 334368
rect 170804 334310 174103 334312
rect 139629 334307 139695 334310
rect 174037 334307 174103 334310
rect 234113 334370 234179 334373
rect 267785 334370 267851 334373
rect 234113 334368 237044 334370
rect 234113 334312 234118 334368
rect 234174 334312 237044 334368
rect 234113 334310 237044 334312
rect 264828 334368 267851 334370
rect 264828 334312 267790 334368
rect 267846 334312 267851 334368
rect 264828 334310 267851 334312
rect 234113 334307 234179 334310
rect 267785 334307 267851 334310
rect 326573 334370 326639 334373
rect 326573 334368 331068 334370
rect 326573 334312 326578 334368
rect 326634 334312 331068 334368
rect 326573 334310 331068 334312
rect 326573 334307 326639 334310
rect 80105 334098 80171 334101
rect 76198 334096 80171 334098
rect 76198 334040 80110 334096
rect 80166 334040 80171 334096
rect 76198 334038 80171 334040
rect 80105 334035 80171 334038
rect 139629 333962 139695 333965
rect 234297 333962 234363 333965
rect 326757 333962 326823 333965
rect 139629 333960 143050 333962
rect 139629 333904 139634 333960
rect 139690 333904 143050 333960
rect 139629 333902 143050 333904
rect 139629 333899 139695 333902
rect 95193 333826 95259 333829
rect 104894 333826 104900 333828
rect 95193 333824 104900 333826
rect 95193 333768 95198 333824
rect 95254 333768 104900 333824
rect 95193 333766 104900 333768
rect 95193 333763 95259 333766
rect 104894 333764 104900 333766
rect 104964 333764 104970 333828
rect 80197 333690 80263 333693
rect 76382 333688 80263 333690
rect 76382 333632 80202 333688
rect 80258 333632 80263 333688
rect 76382 333630 80263 333632
rect 76382 333252 76442 333630
rect 80197 333627 80263 333630
rect 142990 333320 143050 333902
rect 234297 333960 237074 333962
rect 234297 333904 234302 333960
rect 234358 333904 237074 333960
rect 234297 333902 237074 333904
rect 234297 333899 234363 333902
rect 212166 333492 212172 333556
rect 212236 333554 212242 333556
rect 212309 333554 212375 333557
rect 231813 333556 231879 333557
rect 231813 333554 231860 333556
rect 212236 333552 212375 333554
rect 212236 333496 212314 333552
rect 212370 333496 212375 333552
rect 212236 333494 212375 333496
rect 231768 333552 231860 333554
rect 231768 333496 231818 333552
rect 231768 333494 231860 333496
rect 212236 333492 212242 333494
rect 212309 333491 212375 333494
rect 231813 333492 231860 333494
rect 231924 333492 231930 333556
rect 231813 333491 231879 333492
rect 237014 333320 237074 333902
rect 326757 333960 331098 333962
rect 326757 333904 326762 333960
rect 326818 333904 331098 333960
rect 326757 333902 331098 333904
rect 326757 333899 326823 333902
rect 306241 333556 306307 333557
rect 306190 333492 306196 333556
rect 306260 333554 306307 333556
rect 306260 333552 306352 333554
rect 306302 333496 306352 333552
rect 306260 333494 306352 333496
rect 306260 333492 306307 333494
rect 306241 333491 306307 333492
rect 331038 333320 331098 333902
rect 173669 333282 173735 333285
rect 267325 333282 267391 333285
rect 170804 333280 173735 333282
rect 170804 333224 173674 333280
rect 173730 333224 173735 333280
rect 170804 333222 173735 333224
rect 264828 333280 267391 333282
rect 264828 333224 267330 333280
rect 267386 333224 267391 333280
rect 264828 333222 267391 333224
rect 173669 333219 173735 333222
rect 267325 333219 267391 333222
rect 280246 333084 280252 333148
rect 280316 333146 280322 333148
rect 282873 333146 282939 333149
rect 280316 333144 282939 333146
rect 280316 333088 282878 333144
rect 282934 333088 282939 333144
rect 280316 333086 282939 333088
rect 280316 333084 280322 333086
rect 282873 333083 282939 333086
rect 296213 333146 296279 333149
rect 319305 333146 319371 333149
rect 319857 333146 319923 333149
rect 296213 333144 319923 333146
rect 296213 333088 296218 333144
rect 296274 333088 319310 333144
rect 319366 333088 319862 333144
rect 319918 333088 319923 333144
rect 296213 333086 319923 333088
rect 296213 333083 296279 333086
rect 319305 333083 319371 333086
rect 319857 333083 319923 333086
rect 139629 333010 139695 333013
rect 233929 333010 233995 333013
rect 327309 333010 327375 333013
rect 139629 333008 143050 333010
rect 139629 332952 139634 333008
rect 139690 332952 143050 333008
rect 139629 332950 143050 332952
rect 139629 332947 139695 332950
rect 80197 332738 80263 332741
rect 76382 332736 80263 332738
rect 76382 332680 80202 332736
rect 80258 332680 80263 332736
rect 76382 332678 80263 332680
rect 76382 332300 76442 332678
rect 80197 332675 80263 332678
rect 142990 332368 143050 332950
rect 233929 333008 237074 333010
rect 233929 332952 233934 333008
rect 233990 332952 237074 333008
rect 233929 332950 237074 332952
rect 233929 332947 233995 332950
rect 237014 332368 237074 332950
rect 327309 333008 331098 333010
rect 327309 332952 327314 333008
rect 327370 332952 331098 333008
rect 327309 332950 331098 332952
rect 327309 332947 327375 332950
rect 331038 332368 331098 332950
rect 172841 332330 172907 332333
rect 267141 332330 267207 332333
rect 170804 332328 172907 332330
rect 170804 332272 172846 332328
rect 172902 332272 172907 332328
rect 170804 332270 172907 332272
rect 264828 332328 267207 332330
rect 264828 332272 267146 332328
rect 267202 332272 267207 332328
rect 264828 332270 267207 332272
rect 172841 332267 172907 332270
rect 267141 332267 267207 332270
rect 136869 332194 136935 332197
rect 198785 332196 198851 332197
rect 137278 332194 137284 332196
rect 136869 332192 137284 332194
rect 136869 332136 136874 332192
rect 136930 332136 137284 332192
rect 136869 332134 137284 332136
rect 136869 332131 136935 332134
rect 137278 332132 137284 332134
rect 137348 332132 137354 332196
rect 198734 332132 198740 332196
rect 198804 332194 198851 332196
rect 230893 332194 230959 332197
rect 231353 332194 231419 332197
rect 231854 332194 231860 332196
rect 198804 332192 198896 332194
rect 198846 332136 198896 332192
rect 198804 332134 198896 332136
rect 230893 332192 231860 332194
rect 230893 332136 230898 332192
rect 230954 332136 231358 332192
rect 231414 332136 231860 332192
rect 230893 332134 231860 332136
rect 198804 332132 198851 332134
rect 198785 332131 198851 332132
rect 230893 332131 230959 332134
rect 231353 332131 231419 332134
rect 231854 332132 231860 332134
rect 231924 332132 231930 332196
rect 296070 332132 296076 332196
rect 296140 332194 296146 332196
rect 296213 332194 296279 332197
rect 296140 332192 296279 332194
rect 296140 332136 296218 332192
rect 296274 332136 296279 332192
rect 296140 332134 296279 332136
rect 296140 332132 296146 332134
rect 296213 332131 296279 332134
rect 139813 331650 139879 331653
rect 139813 331648 143050 331650
rect 139813 331592 139818 331648
rect 139874 331592 143050 331648
rect 139813 331590 143050 331592
rect 139813 331587 139879 331590
rect 137053 331514 137119 331517
rect 137278 331514 137284 331516
rect 137053 331512 137284 331514
rect 137053 331456 137058 331512
rect 137114 331456 137284 331512
rect 137053 331454 137284 331456
rect 137053 331451 137119 331454
rect 137278 331452 137284 331454
rect 137348 331452 137354 331516
rect 142990 331280 143050 331590
rect 204438 331588 204444 331652
rect 204508 331650 204514 331652
rect 205593 331650 205659 331653
rect 225281 331650 225347 331653
rect 204508 331648 225347 331650
rect 204508 331592 205598 331648
rect 205654 331592 225286 331648
rect 225342 331592 225347 331648
rect 204508 331590 225347 331592
rect 204508 331588 204514 331590
rect 205593 331587 205659 331590
rect 225281 331587 225347 331590
rect 292901 331650 292967 331653
rect 294046 331650 294052 331652
rect 292901 331648 294052 331650
rect 292901 331592 292906 331648
rect 292962 331592 294052 331648
rect 292901 331590 294052 331592
rect 292901 331587 292967 331590
rect 294046 331588 294052 331590
rect 294116 331650 294122 331652
rect 319397 331650 319463 331653
rect 319673 331650 319739 331653
rect 294116 331648 319739 331650
rect 294116 331592 319402 331648
rect 319458 331592 319678 331648
rect 319734 331592 319739 331648
rect 294116 331590 319739 331592
rect 294116 331588 294122 331590
rect 319397 331587 319463 331590
rect 319673 331587 319739 331590
rect 230801 331514 230867 331517
rect 231445 331514 231511 331517
rect 231854 331514 231860 331516
rect 230801 331512 231860 331514
rect 230801 331456 230806 331512
rect 230862 331456 231450 331512
rect 231506 331456 231860 331512
rect 230801 331454 231860 331456
rect 230801 331451 230867 331454
rect 231445 331451 231511 331454
rect 231854 331452 231860 331454
rect 231924 331452 231930 331516
rect 233469 331514 233535 331517
rect 328505 331514 328571 331517
rect 233469 331512 237074 331514
rect 233469 331456 233474 331512
rect 233530 331456 237074 331512
rect 233469 331454 237074 331456
rect 233469 331451 233535 331454
rect 237014 331280 237074 331454
rect 328505 331512 331098 331514
rect 328505 331456 328510 331512
rect 328566 331456 331098 331512
rect 328505 331454 331098 331456
rect 328505 331451 328571 331454
rect 331038 331280 331098 331454
rect 172933 331242 172999 331245
rect 266773 331242 266839 331245
rect 170804 331240 172999 331242
rect 76198 330970 76258 331212
rect 170804 331184 172938 331240
rect 172994 331184 172999 331240
rect 170804 331182 172999 331184
rect 264828 331240 266839 331242
rect 264828 331184 266778 331240
rect 266834 331184 266839 331240
rect 264828 331182 266839 331184
rect 172933 331179 172999 331182
rect 266773 331179 266839 331182
rect 80197 330970 80263 330973
rect 76198 330968 80263 330970
rect 76198 330912 80202 330968
rect 80258 330912 80263 330968
rect 76198 330910 80263 330912
rect 80197 330907 80263 330910
rect 140549 330290 140615 330293
rect 173393 330290 173459 330293
rect 140549 330288 143020 330290
rect 76198 329746 76258 330260
rect 140549 330232 140554 330288
rect 140610 330232 143020 330288
rect 140549 330230 143020 330232
rect 170804 330288 173459 330290
rect 170804 330232 173398 330288
rect 173454 330232 173459 330288
rect 170804 330230 173459 330232
rect 140549 330227 140615 330230
rect 173393 330227 173459 330230
rect 233469 330290 233535 330293
rect 267877 330290 267943 330293
rect 233469 330288 237044 330290
rect 233469 330232 233474 330288
rect 233530 330232 237044 330288
rect 233469 330230 237044 330232
rect 264828 330288 267943 330290
rect 264828 330232 267882 330288
rect 267938 330232 267943 330288
rect 264828 330230 267943 330232
rect 233469 330227 233535 330230
rect 267877 330227 267943 330230
rect 319581 330290 319647 330293
rect 319581 330288 331068 330290
rect 319581 330232 319586 330288
rect 319642 330232 331068 330288
rect 319581 330230 331068 330232
rect 319581 330227 319647 330230
rect 159593 330156 159659 330157
rect 159542 330092 159548 330156
rect 159612 330154 159659 330156
rect 159612 330152 159704 330154
rect 159654 330096 159704 330152
rect 159612 330094 159704 330096
rect 159612 330092 159659 330094
rect 252278 330092 252284 330156
rect 252348 330154 252354 330156
rect 252605 330154 252671 330157
rect 252348 330152 252671 330154
rect 252348 330096 252610 330152
rect 252666 330096 252671 330152
rect 252348 330094 252671 330096
rect 252348 330092 252354 330094
rect 159593 330091 159659 330092
rect 252605 330091 252671 330094
rect 251542 329956 251548 330020
rect 251612 330018 251618 330020
rect 251961 330018 252027 330021
rect 253014 330018 253020 330020
rect 251612 330016 253020 330018
rect 251612 329960 251966 330016
rect 252022 329960 253020 330016
rect 251612 329958 253020 329960
rect 251612 329956 251618 329958
rect 251961 329955 252027 329958
rect 253014 329956 253020 329958
rect 253084 329956 253090 330020
rect 82313 329746 82379 329749
rect 76198 329744 82379 329746
rect 76198 329688 82318 329744
rect 82374 329688 82379 329744
rect 76198 329686 82379 329688
rect 82313 329683 82379 329686
rect 161709 329476 161775 329477
rect 161709 329474 161756 329476
rect 161664 329472 161756 329474
rect 161664 329416 161714 329472
rect 161664 329414 161756 329416
rect 161709 329412 161756 329414
rect 161820 329412 161826 329476
rect 161709 329411 161775 329412
rect 430165 327978 430231 327981
rect 434416 327978 434896 328008
rect 430165 327976 434896 327978
rect 430165 327920 430170 327976
rect 430226 327920 434896 327976
rect 430165 327918 434896 327920
rect 430165 327915 430231 327918
rect 434416 327888 434896 327918
rect 256009 327570 256075 327573
rect 262398 327570 262404 327572
rect 256009 327568 262404 327570
rect 256009 327512 256014 327568
rect 256070 327512 262404 327568
rect 256009 327510 262404 327512
rect 256009 327507 256075 327510
rect 262398 327508 262404 327510
rect 262468 327508 262474 327572
rect 52638 327372 52644 327436
rect 52708 327434 52714 327436
rect 53057 327434 53123 327437
rect 52708 327432 53123 327434
rect 52708 327376 53062 327432
rect 53118 327376 53123 327432
rect 52708 327374 53123 327376
rect 52708 327372 52714 327374
rect 53057 327371 53123 327374
rect 54069 327434 54135 327437
rect 54662 327434 54668 327436
rect 54069 327432 54668 327434
rect 54069 327376 54074 327432
rect 54130 327376 54668 327432
rect 54069 327374 54668 327376
rect 54069 327371 54135 327374
rect 54662 327372 54668 327374
rect 54732 327372 54738 327436
rect 55398 327372 55404 327436
rect 55468 327434 55474 327436
rect 56093 327434 56159 327437
rect 55468 327432 56159 327434
rect 55468 327376 56098 327432
rect 56154 327376 56159 327432
rect 55468 327374 56159 327376
rect 55468 327372 55474 327374
rect 56093 327371 56159 327374
rect 158121 327434 158187 327437
rect 168558 327434 168564 327436
rect 158121 327432 168564 327434
rect 158121 327376 158126 327432
rect 158182 327376 168564 327432
rect 158121 327374 168564 327376
rect 158121 327371 158187 327374
rect 168558 327372 168564 327374
rect 168628 327372 168634 327436
rect 339177 327434 339243 327437
rect 339494 327434 339500 327436
rect 339177 327432 339500 327434
rect 339177 327376 339182 327432
rect 339238 327376 339500 327432
rect 339177 327374 339500 327376
rect 339177 327371 339243 327374
rect 339494 327372 339500 327374
rect 339564 327372 339570 327436
rect 340005 327434 340071 327437
rect 340966 327434 340972 327436
rect 340005 327432 340972 327434
rect 340005 327376 340010 327432
rect 340066 327376 340972 327432
rect 340005 327374 340972 327376
rect 340005 327371 340071 327374
rect 340966 327372 340972 327374
rect 341036 327372 341042 327436
rect 153245 326348 153311 326349
rect 153245 326344 153292 326348
rect 153356 326346 153362 326348
rect 153245 326288 153250 326344
rect 153245 326284 153292 326288
rect 153356 326286 153402 326346
rect 153356 326284 153362 326286
rect 153245 326283 153311 326284
rect 9896 323218 10376 323248
rect 13957 323218 14023 323221
rect 9896 323216 14023 323218
rect 9896 323160 13962 323216
rect 14018 323160 14023 323216
rect 9896 323158 14023 323160
rect 9896 323128 10376 323158
rect 13957 323155 14023 323158
rect 137881 320362 137947 320365
rect 230985 320362 231051 320365
rect 324549 320362 324615 320365
rect 134740 320360 137947 320362
rect 134740 320304 137886 320360
rect 137942 320304 137947 320360
rect 134740 320302 137947 320304
rect 228764 320360 231051 320362
rect 228764 320304 230990 320360
rect 231046 320304 231051 320360
rect 228764 320302 231051 320304
rect 322788 320360 324615 320362
rect 322788 320304 324554 320360
rect 324610 320304 324615 320360
rect 322788 320302 324615 320304
rect 137881 320299 137947 320302
rect 230985 320299 231051 320302
rect 324549 320299 324615 320302
rect 54069 317914 54135 317917
rect 55214 317914 55220 317916
rect 54069 317912 55220 317914
rect 54069 317856 54074 317912
rect 54130 317856 55220 317912
rect 54069 317854 55220 317856
rect 54069 317851 54135 317854
rect 55214 317852 55220 317854
rect 55284 317852 55290 317916
rect 137697 317234 137763 317237
rect 231445 317234 231511 317237
rect 324733 317234 324799 317237
rect 134740 317232 137763 317234
rect 134740 317176 137702 317232
rect 137758 317176 137763 317232
rect 134740 317174 137763 317176
rect 228764 317232 231511 317234
rect 228764 317176 231450 317232
rect 231506 317176 231511 317232
rect 228764 317174 231511 317176
rect 322788 317232 324799 317234
rect 322788 317176 324738 317232
rect 324794 317176 324799 317232
rect 322788 317174 324799 317176
rect 137697 317171 137763 317174
rect 231445 317171 231511 317174
rect 324733 317171 324799 317174
rect 52689 315874 52755 315877
rect 55398 315874 55404 315876
rect 52689 315872 55404 315874
rect 52689 315816 52694 315872
rect 52750 315816 55404 315872
rect 52689 315814 55404 315816
rect 52689 315811 52755 315814
rect 55398 315812 55404 315814
rect 55468 315812 55474 315876
rect 153286 315812 153292 315876
rect 153356 315874 153362 315876
rect 165113 315874 165179 315877
rect 153356 315872 165179 315874
rect 153356 315816 165118 315872
rect 165174 315816 165179 315872
rect 153356 315814 165179 315816
rect 153356 315812 153362 315814
rect 165113 315811 165179 315814
rect 405969 315874 406035 315877
rect 405969 315872 409114 315874
rect 405969 315816 405974 315872
rect 406030 315816 409114 315872
rect 405969 315814 409114 315816
rect 405969 315811 406035 315814
rect 38797 315602 38863 315605
rect 35748 315600 38863 315602
rect 35748 315544 38802 315600
rect 38858 315544 38863 315600
rect 409054 315572 409114 315814
rect 35748 315542 38863 315544
rect 38797 315539 38863 315542
rect 429429 315466 429495 315469
rect 434416 315466 434896 315496
rect 429429 315464 434896 315466
rect 429429 315408 429434 315464
rect 429490 315408 434896 315464
rect 429429 315406 434896 315408
rect 429429 315403 429495 315406
rect 434416 315376 434896 315406
rect 70862 314514 70922 315028
rect 340966 314860 340972 314924
rect 341036 314922 341042 314924
rect 351822 314922 351828 314924
rect 341036 314862 351828 314922
rect 341036 314860 341042 314862
rect 351822 314860 351828 314862
rect 351892 314860 351898 314924
rect 339494 314588 339500 314652
rect 339564 314588 339570 314652
rect 74217 314514 74283 314517
rect 70862 314512 74283 314514
rect 70862 314456 74222 314512
rect 74278 314456 74283 314512
rect 70862 314454 74283 314456
rect 339502 314514 339562 314588
rect 352558 314514 352564 314516
rect 339502 314454 352564 314514
rect 74217 314451 74283 314454
rect 352558 314452 352564 314454
rect 352628 314452 352634 314516
rect 16073 313834 16139 313837
rect 19894 313834 19954 314348
rect 16073 313832 19954 313834
rect 16073 313776 16078 313832
rect 16134 313776 19954 313832
rect 16073 313774 19954 313776
rect 51217 313834 51283 313837
rect 55038 313834 55098 314280
rect 137053 314106 137119 314109
rect 231353 314106 231419 314109
rect 325837 314106 325903 314109
rect 134740 314104 137119 314106
rect 134740 314048 137058 314104
rect 137114 314048 137119 314104
rect 134740 314046 137119 314048
rect 228764 314104 231419 314106
rect 228764 314048 231358 314104
rect 231414 314048 231419 314104
rect 228764 314046 231419 314048
rect 322788 314104 325903 314106
rect 322788 314048 325842 314104
rect 325898 314048 325903 314104
rect 322788 314046 325903 314048
rect 352750 314106 352810 314280
rect 356197 314106 356263 314109
rect 352750 314104 356263 314106
rect 352750 314048 356202 314104
rect 356258 314048 356263 314104
rect 352750 314046 356263 314048
rect 137053 314043 137119 314046
rect 231353 314043 231419 314046
rect 325837 314043 325903 314046
rect 356197 314043 356263 314046
rect 51217 313832 55098 313834
rect 51217 313776 51222 313832
rect 51278 313776 55098 313832
rect 51217 313774 55098 313776
rect 424694 313834 424754 314280
rect 427313 313834 427379 313837
rect 424694 313832 427379 313834
rect 424694 313776 427318 313832
rect 427374 313776 427379 313832
rect 424694 313774 427379 313776
rect 16073 313771 16139 313774
rect 51217 313771 51283 313774
rect 427313 313771 427379 313774
rect 405969 313698 406035 313701
rect 405969 313696 409114 313698
rect 405969 313640 405974 313696
rect 406030 313640 409114 313696
rect 405969 313638 409114 313640
rect 405969 313635 406035 313638
rect 81669 313562 81735 313565
rect 175509 313562 175575 313565
rect 270269 313562 270335 313565
rect 81669 313560 85060 313562
rect 81669 313504 81674 313560
rect 81730 313504 85060 313560
rect 81669 313502 85060 313504
rect 175509 313560 178900 313562
rect 175509 313504 175514 313560
rect 175570 313504 178900 313560
rect 175509 313502 178900 313504
rect 270269 313560 272924 313562
rect 270269 313504 270274 313560
rect 270330 313504 272924 313560
rect 270269 313502 272924 313504
rect 81669 313499 81735 313502
rect 175509 313499 175575 313502
rect 270269 313499 270335 313502
rect 38429 313154 38495 313157
rect 35748 313152 38495 313154
rect 35748 313096 38434 313152
rect 38490 313096 38495 313152
rect 409054 313124 409114 313638
rect 35748 313094 38495 313096
rect 38429 313091 38495 313094
rect 70862 311114 70922 311356
rect 74125 311114 74191 311117
rect 70862 311112 74191 311114
rect 70862 311056 74130 311112
rect 74186 311056 74191 311112
rect 70862 311054 74191 311056
rect 74125 311051 74191 311054
rect 137513 310978 137579 310981
rect 230893 310978 230959 310981
rect 325193 310978 325259 310981
rect 134740 310976 137579 310978
rect 134740 310920 137518 310976
rect 137574 310920 137579 310976
rect 134740 310918 137579 310920
rect 228764 310976 230959 310978
rect 228764 310920 230898 310976
rect 230954 310920 230959 310976
rect 228764 310918 230959 310920
rect 322788 310976 325259 310978
rect 322788 310920 325198 310976
rect 325254 310920 325259 310976
rect 322788 310918 325259 310920
rect 137513 310915 137579 310918
rect 230893 310915 230959 310918
rect 325193 310915 325259 310918
rect 35718 310434 35778 310472
rect 38797 310434 38863 310437
rect 35718 310432 38863 310434
rect 35718 310376 38802 310432
rect 38858 310376 38863 310432
rect 35718 310374 38863 310376
rect 38797 310371 38863 310374
rect 54069 310434 54135 310437
rect 55030 310434 55036 310436
rect 54069 310432 55036 310434
rect 54069 310376 54074 310432
rect 54130 310376 55036 310432
rect 54069 310374 55036 310376
rect 54069 310371 54135 310374
rect 55030 310372 55036 310374
rect 55100 310372 55106 310436
rect 405969 310434 406035 310437
rect 408870 310434 408930 310540
rect 405969 310432 408930 310434
rect 405969 310376 405974 310432
rect 406030 310376 408930 310432
rect 405969 310374 408930 310376
rect 405969 310371 406035 310374
rect 148326 310170 148908 310230
rect 242350 310170 242932 310230
rect 145517 310162 145583 310165
rect 148326 310162 148386 310170
rect 145517 310160 148386 310162
rect 145517 310104 145522 310160
rect 145578 310104 148386 310160
rect 145517 310102 148386 310104
rect 240645 310162 240711 310165
rect 242350 310162 242410 310170
rect 240645 310160 242410 310162
rect 240645 310104 240650 310160
rect 240706 310104 242410 310160
rect 240645 310102 242410 310104
rect 145517 310099 145583 310102
rect 240645 310099 240711 310102
rect 9896 309890 10376 309920
rect 13957 309890 14023 309893
rect 9896 309888 14023 309890
rect 9896 309832 13962 309888
rect 14018 309832 14023 309888
rect 9896 309830 14023 309832
rect 9896 309800 10376 309830
rect 13957 309827 14023 309830
rect 334209 309754 334275 309757
rect 336926 309754 336986 310200
rect 334209 309752 336986 309754
rect 334209 309696 334214 309752
rect 334270 309696 336986 309752
rect 334209 309694 336986 309696
rect 334209 309691 334275 309694
rect 16165 308394 16231 308397
rect 19894 308394 19954 309316
rect 51217 308666 51283 308669
rect 55038 308666 55098 309248
rect 51217 308664 55098 308666
rect 51217 308608 51222 308664
rect 51278 308608 55098 308664
rect 51217 308606 55098 308608
rect 352750 308666 352810 309248
rect 356197 308666 356263 308669
rect 352750 308664 356263 308666
rect 352750 308608 356202 308664
rect 356258 308608 356263 308664
rect 352750 308606 356263 308608
rect 424694 308666 424754 309248
rect 428693 308666 428759 308669
rect 424694 308664 428759 308666
rect 424694 308608 428698 308664
rect 428754 308608 428759 308664
rect 424694 308606 428759 308608
rect 51217 308603 51283 308606
rect 356197 308603 356263 308606
rect 428693 308603 428759 308606
rect 16165 308392 19954 308394
rect 16165 308336 16170 308392
rect 16226 308336 19954 308392
rect 16165 308334 19954 308336
rect 16165 308331 16231 308334
rect 405969 308258 406035 308261
rect 405969 308256 409114 308258
rect 405969 308200 405974 308256
rect 406030 308200 409114 308256
rect 405969 308198 409114 308200
rect 405969 308195 406035 308198
rect 38797 308122 38863 308125
rect 35748 308120 38863 308122
rect 35748 308064 38802 308120
rect 38858 308064 38863 308120
rect 409054 308092 409114 308198
rect 35748 308062 38863 308064
rect 38797 308059 38863 308062
rect 136869 307850 136935 307853
rect 230801 307850 230867 307853
rect 325745 307850 325811 307853
rect 134740 307848 136935 307850
rect 134740 307792 136874 307848
rect 136930 307792 136935 307848
rect 134740 307790 136935 307792
rect 228764 307848 230867 307850
rect 228764 307792 230806 307848
rect 230862 307792 230867 307848
rect 228764 307790 230867 307792
rect 322788 307848 325811 307850
rect 322788 307792 325750 307848
rect 325806 307792 325811 307848
rect 322788 307790 325811 307792
rect 136869 307787 136935 307790
rect 230801 307787 230867 307790
rect 325745 307787 325811 307790
rect 70862 307170 70922 307684
rect 73389 307170 73455 307173
rect 70862 307168 73455 307170
rect 70862 307112 73394 307168
rect 73450 307112 73455 307168
rect 70862 307110 73455 307112
rect 73389 307107 73455 307110
rect 54437 306218 54503 306221
rect 54662 306218 54668 306220
rect 54437 306216 54668 306218
rect 54437 306160 54442 306216
rect 54498 306160 54668 306216
rect 54437 306158 54668 306160
rect 54437 306155 54503 306158
rect 54662 306156 54668 306158
rect 54732 306156 54738 306220
rect 164702 306218 164762 306800
rect 167873 306218 167939 306221
rect 164702 306216 167939 306218
rect 164702 306160 167878 306216
rect 167934 306160 167939 306216
rect 164702 306158 167939 306160
rect 258726 306218 258786 306800
rect 261713 306218 261779 306221
rect 258726 306216 261779 306218
rect 258726 306160 261718 306216
rect 261774 306160 261779 306216
rect 258726 306158 261779 306160
rect 167873 306155 167939 306158
rect 261713 306155 261779 306158
rect 406061 306218 406127 306221
rect 406061 306216 409114 306218
rect 406061 306160 406066 306216
rect 406122 306160 409114 306216
rect 406061 306158 409114 306160
rect 406061 306155 406127 306158
rect 38797 305674 38863 305677
rect 35748 305672 38863 305674
rect 35748 305616 38802 305672
rect 38858 305616 38863 305672
rect 35748 305614 38863 305616
rect 38797 305611 38863 305614
rect 73389 305674 73455 305677
rect 74534 305674 74540 305676
rect 73389 305672 74540 305674
rect 73389 305616 73394 305672
rect 73450 305616 74540 305672
rect 73389 305614 74540 305616
rect 73389 305611 73455 305614
rect 74534 305612 74540 305614
rect 74604 305674 74610 305676
rect 76885 305674 76951 305677
rect 74604 305672 76951 305674
rect 74604 305616 76890 305672
rect 76946 305616 76951 305672
rect 409054 305644 409114 306158
rect 74604 305614 76951 305616
rect 74604 305612 74610 305614
rect 76885 305611 76951 305614
rect 325101 305538 325167 305541
rect 325469 305538 325535 305541
rect 325101 305536 325535 305538
rect 325101 305480 325106 305536
rect 325162 305480 325474 305536
rect 325530 305480 325535 305536
rect 325101 305478 325535 305480
rect 325101 305475 325167 305478
rect 325469 305475 325535 305478
rect 325561 305402 325627 305405
rect 322758 305400 325627 305402
rect 322758 305344 325566 305400
rect 325622 305344 325627 305400
rect 322758 305342 325627 305344
rect 231997 304722 232063 304725
rect 228764 304720 232063 304722
rect 228764 304664 232002 304720
rect 232058 304664 232063 304720
rect 322758 304692 322818 305342
rect 325561 305339 325627 305342
rect 228764 304662 232063 304664
rect 231997 304659 232063 304662
rect 16257 304178 16323 304181
rect 19894 304178 19954 304284
rect 70678 304254 74050 304314
rect 16257 304176 19954 304178
rect 16257 304120 16262 304176
rect 16318 304120 19954 304176
rect 16257 304118 19954 304120
rect 51401 304178 51467 304181
rect 55038 304178 55098 304216
rect 51401 304176 55098 304178
rect 51401 304120 51406 304176
rect 51462 304120 55098 304176
rect 70678 304148 70738 304254
rect 51401 304118 55098 304120
rect 16257 304115 16323 304118
rect 51401 304115 51467 304118
rect 73990 304044 74050 304254
rect 134710 304178 134770 304624
rect 136961 304178 137027 304181
rect 137513 304178 137579 304181
rect 134710 304176 137579 304178
rect 134710 304120 136966 304176
rect 137022 304120 137518 304176
rect 137574 304120 137579 304176
rect 134710 304118 137579 304120
rect 352750 304178 352810 304216
rect 356197 304178 356263 304181
rect 352750 304176 356263 304178
rect 352750 304120 356202 304176
rect 356258 304120 356263 304176
rect 352750 304118 356263 304120
rect 424694 304178 424754 304216
rect 427405 304178 427471 304181
rect 424694 304176 427471 304178
rect 424694 304120 427410 304176
rect 427466 304120 427471 304176
rect 424694 304118 427471 304120
rect 136961 304115 137027 304118
rect 137513 304115 137579 304118
rect 356197 304115 356263 304118
rect 427405 304115 427471 304118
rect 73982 303980 73988 304044
rect 74052 304042 74058 304044
rect 75505 304042 75571 304045
rect 74052 304040 75571 304042
rect 74052 303984 75510 304040
rect 75566 303984 75571 304040
rect 74052 303982 75571 303984
rect 74052 303980 74058 303982
rect 75505 303979 75571 303982
rect 405969 303634 406035 303637
rect 405969 303632 409114 303634
rect 405969 303576 405974 303632
rect 406030 303576 409114 303632
rect 405969 303574 409114 303576
rect 405969 303571 406035 303574
rect 38613 303090 38679 303093
rect 35748 303088 38679 303090
rect 35748 303032 38618 303088
rect 38674 303032 38679 303088
rect 409054 303060 409114 303574
rect 35748 303030 38679 303032
rect 38613 303027 38679 303030
rect 430165 302954 430231 302957
rect 434416 302954 434896 302984
rect 430165 302952 434896 302954
rect 430165 302896 430170 302952
rect 430226 302896 434896 302952
rect 430165 302894 434896 302896
rect 430165 302891 430231 302894
rect 434416 302864 434896 302894
rect 136869 301594 136935 301597
rect 137789 301594 137855 301597
rect 231997 301594 232063 301597
rect 325653 301594 325719 301597
rect 134740 301592 137855 301594
rect 134740 301536 136874 301592
rect 136930 301536 137794 301592
rect 137850 301536 137855 301592
rect 134740 301534 137855 301536
rect 228764 301592 232063 301594
rect 228764 301536 232002 301592
rect 232058 301536 232063 301592
rect 228764 301534 232063 301536
rect 322788 301592 325719 301594
rect 322788 301536 325658 301592
rect 325714 301536 325719 301592
rect 322788 301534 325719 301536
rect 136869 301531 136935 301534
rect 137789 301531 137855 301534
rect 231997 301531 232063 301534
rect 325653 301531 325719 301534
rect 38797 300642 38863 300645
rect 35748 300640 38863 300642
rect 35748 300584 38802 300640
rect 38858 300584 38863 300640
rect 35748 300582 38863 300584
rect 38797 300579 38863 300582
rect 50297 300642 50363 300645
rect 52638 300642 52644 300644
rect 50297 300640 52644 300642
rect 50297 300584 50302 300640
rect 50358 300584 52644 300640
rect 50297 300582 52644 300584
rect 50297 300579 50363 300582
rect 52638 300580 52644 300582
rect 52708 300580 52714 300644
rect 405969 300506 406035 300509
rect 408870 300506 408930 300612
rect 405969 300504 408930 300506
rect 70862 300098 70922 300476
rect 405969 300448 405974 300504
rect 406030 300448 408930 300504
rect 405969 300446 408930 300448
rect 405969 300443 406035 300446
rect 73798 300098 73804 300100
rect 70862 300038 73804 300098
rect 73798 300036 73804 300038
rect 73868 300036 73874 300100
rect 73806 299962 73866 300036
rect 75413 299962 75479 299965
rect 73806 299960 75479 299962
rect 73806 299904 75418 299960
rect 75474 299904 75479 299960
rect 73806 299902 75479 299904
rect 75413 299899 75479 299902
rect 16441 298738 16507 298741
rect 19894 298738 19954 299388
rect 51401 298874 51467 298877
rect 55038 298874 55098 299320
rect 51401 298872 55098 298874
rect 51401 298816 51406 298872
rect 51462 298816 55098 298872
rect 51401 298814 55098 298816
rect 352750 298874 352810 299320
rect 356197 298874 356263 298877
rect 352750 298872 356263 298874
rect 352750 298816 356202 298872
rect 356258 298816 356263 298872
rect 352750 298814 356263 298816
rect 51401 298811 51467 298814
rect 356197 298811 356263 298814
rect 16441 298736 19954 298738
rect 16441 298680 16446 298736
rect 16502 298680 19954 298736
rect 16441 298678 19954 298680
rect 424694 298738 424754 299320
rect 427497 298738 427563 298741
rect 424694 298736 427563 298738
rect 424694 298680 427502 298736
rect 427558 298680 427563 298736
rect 424694 298678 427563 298680
rect 16441 298675 16507 298678
rect 427497 298675 427563 298678
rect 137605 298602 137671 298605
rect 134710 298600 137671 298602
rect 134710 298544 137610 298600
rect 137666 298544 137671 298600
rect 134710 298542 137671 298544
rect 38245 298194 38311 298197
rect 134710 298196 134770 298542
rect 137605 298539 137671 298542
rect 230709 298466 230775 298469
rect 325101 298466 325167 298469
rect 228764 298464 230775 298466
rect 228764 298408 230714 298464
rect 230770 298408 230775 298464
rect 228764 298406 230775 298408
rect 322788 298464 325167 298466
rect 322788 298408 325106 298464
rect 325162 298408 325167 298464
rect 322788 298406 325167 298408
rect 230709 298403 230775 298406
rect 325101 298403 325167 298406
rect 405969 298330 406035 298333
rect 405969 298328 409114 298330
rect 405969 298272 405974 298328
rect 406030 298272 409114 298328
rect 405969 298270 409114 298272
rect 405969 298267 406035 298270
rect 35748 298192 38311 298194
rect 35748 298136 38250 298192
rect 38306 298136 38311 298192
rect 35748 298134 38311 298136
rect 38245 298131 38311 298134
rect 134702 298132 134708 298196
rect 134772 298132 134778 298196
rect 409054 298164 409114 298270
rect 352793 297242 352859 297245
rect 353989 297242 354055 297245
rect 352793 297240 354055 297242
rect 352793 297184 352798 297240
rect 352854 297184 353994 297240
rect 354050 297184 354055 297240
rect 352793 297182 354055 297184
rect 352793 297179 352859 297182
rect 353989 297179 354055 297182
rect 74217 296970 74283 296973
rect 75965 296970 76031 296973
rect 70678 296968 76031 296970
rect 70678 296912 74222 296968
rect 74278 296912 75970 296968
rect 76026 296912 76031 296968
rect 70678 296910 76031 296912
rect 70678 296804 70738 296910
rect 74217 296907 74283 296910
rect 75965 296907 76031 296910
rect 148326 296842 148908 296902
rect 242350 296842 242932 296902
rect 81669 296834 81735 296837
rect 145425 296834 145491 296837
rect 148326 296834 148386 296842
rect 81669 296832 85060 296834
rect 81669 296776 81674 296832
rect 81730 296776 85060 296832
rect 81669 296774 85060 296776
rect 145425 296832 148386 296834
rect 145425 296776 145430 296832
rect 145486 296776 148386 296832
rect 145425 296774 148386 296776
rect 175509 296834 175575 296837
rect 240921 296834 240987 296837
rect 242350 296834 242410 296842
rect 175509 296832 178900 296834
rect 175509 296776 175514 296832
rect 175570 296776 178900 296832
rect 175509 296774 178900 296776
rect 240921 296832 242410 296834
rect 240921 296776 240926 296832
rect 240982 296776 242410 296832
rect 240921 296774 242410 296776
rect 270361 296834 270427 296837
rect 270361 296832 272924 296834
rect 270361 296776 270366 296832
rect 270422 296776 272924 296832
rect 270361 296774 272924 296776
rect 81669 296771 81735 296774
rect 145425 296771 145491 296774
rect 175509 296771 175575 296774
rect 240921 296771 240987 296774
rect 270361 296771 270427 296774
rect 9896 296426 10376 296456
rect 13681 296426 13747 296429
rect 9896 296424 13747 296426
rect 9896 296368 13686 296424
rect 13742 296368 13747 296424
rect 9896 296366 13747 296368
rect 9896 296336 10376 296366
rect 13681 296363 13747 296366
rect 334209 296290 334275 296293
rect 336926 296290 336986 296872
rect 334209 296288 336986 296290
rect 334209 296232 334214 296288
rect 334270 296232 336986 296288
rect 334209 296230 336986 296232
rect 334209 296227 334275 296230
rect 35718 295474 35778 295512
rect 38797 295474 38863 295477
rect 323486 295474 323492 295476
rect 35718 295472 38863 295474
rect 35718 295416 38802 295472
rect 38858 295416 38863 295472
rect 35718 295414 38863 295416
rect 38797 295411 38863 295414
rect 322758 295414 323492 295474
rect 322758 295308 322818 295414
rect 323486 295412 323492 295414
rect 323556 295412 323562 295476
rect 405969 295474 406035 295477
rect 408870 295474 408930 295580
rect 405969 295472 408930 295474
rect 405969 295416 405974 295472
rect 406030 295416 408930 295472
rect 405969 295414 408930 295416
rect 405969 295411 406035 295414
rect 134710 294794 134770 295240
rect 228734 294796 228794 295240
rect 136910 294794 136916 294796
rect 134710 294734 136916 294794
rect 136910 294732 136916 294734
rect 136980 294732 136986 294796
rect 228726 294732 228732 294796
rect 228796 294732 228802 294796
rect 228734 294658 228794 294732
rect 230801 294658 230867 294661
rect 231854 294658 231860 294660
rect 228734 294656 231860 294658
rect 228734 294600 230806 294656
rect 230862 294600 231860 294656
rect 228734 294598 231860 294600
rect 230801 294595 230867 294598
rect 231854 294596 231860 294598
rect 231924 294596 231930 294660
rect 17453 293842 17519 293845
rect 19894 293842 19954 294356
rect 17453 293840 19954 293842
rect 17453 293784 17458 293840
rect 17514 293784 19954 293840
rect 17453 293782 19954 293784
rect 51309 293842 51375 293845
rect 55038 293842 55098 294288
rect 51309 293840 55098 293842
rect 51309 293784 51314 293840
rect 51370 293784 55098 293840
rect 51309 293782 55098 293784
rect 352750 293842 352810 294288
rect 356197 293842 356263 293845
rect 352750 293840 356263 293842
rect 352750 293784 356202 293840
rect 356258 293784 356263 293840
rect 352750 293782 356263 293784
rect 17453 293779 17519 293782
rect 51309 293779 51375 293782
rect 356197 293779 356263 293782
rect 405969 293706 406035 293709
rect 424694 293706 424754 294288
rect 427589 293706 427655 293709
rect 405969 293704 409114 293706
rect 405969 293648 405974 293704
rect 406030 293648 409114 293704
rect 405969 293646 409114 293648
rect 424694 293704 427655 293706
rect 424694 293648 427594 293704
rect 427650 293648 427655 293704
rect 424694 293646 427655 293648
rect 405969 293643 406035 293646
rect 70678 293238 74234 293298
rect 38429 293162 38495 293165
rect 35748 293160 38495 293162
rect 35748 293104 38434 293160
rect 38490 293104 38495 293160
rect 70678 293132 70738 293238
rect 35748 293102 38495 293104
rect 38429 293099 38495 293102
rect 74174 293028 74234 293238
rect 409054 293132 409114 293646
rect 427589 293643 427655 293646
rect 74166 292964 74172 293028
rect 74236 293026 74242 293028
rect 75873 293026 75939 293029
rect 74236 293024 75939 293026
rect 74236 292968 75878 293024
rect 75934 292968 75939 293024
rect 74236 292966 75939 292968
rect 74236 292964 74242 292966
rect 75873 292963 75939 292966
rect 136910 292210 136916 292212
rect 134740 292150 136916 292210
rect 136910 292148 136916 292150
rect 136980 292148 136986 292212
rect 324549 292210 324615 292213
rect 325285 292210 325351 292213
rect 322788 292208 325351 292210
rect 322788 292180 324554 292208
rect 322758 292152 324554 292180
rect 324610 292152 325290 292208
rect 325346 292152 325351 292208
rect 322758 292150 325351 292152
rect 228764 292082 229162 292142
rect 229102 292074 229162 292082
rect 230750 292074 230756 292076
rect 229102 292014 230756 292074
rect 230750 292012 230756 292014
rect 230820 292012 230826 292076
rect 322758 291940 322818 292150
rect 324549 292147 324615 292150
rect 325285 292147 325351 292150
rect 322750 291876 322756 291940
rect 322820 291876 322826 291940
rect 73430 291740 73436 291804
rect 73500 291802 73506 291804
rect 73982 291802 73988 291804
rect 73500 291742 73988 291802
rect 73500 291740 73506 291742
rect 73982 291740 73988 291742
rect 74052 291740 74058 291804
rect 261110 290652 261116 290716
rect 261180 290714 261186 290716
rect 270494 290714 270500 290716
rect 261180 290654 270500 290714
rect 261180 290652 261186 290654
rect 270494 290652 270500 290654
rect 270564 290652 270570 290716
rect 405969 290714 406035 290717
rect 405969 290712 409114 290714
rect 405969 290656 405974 290712
rect 406030 290656 409114 290712
rect 405969 290654 409114 290656
rect 405969 290651 406035 290654
rect 38613 290578 38679 290581
rect 35748 290576 38679 290578
rect 35748 290520 38618 290576
rect 38674 290520 38679 290576
rect 409054 290548 409114 290654
rect 35748 290518 38679 290520
rect 38613 290515 38679 290518
rect 429429 290442 429495 290445
rect 434416 290442 434896 290472
rect 429429 290440 434896 290442
rect 429429 290384 429434 290440
rect 429490 290384 434896 290440
rect 429429 290382 434896 290384
rect 429429 290379 429495 290382
rect 434416 290352 434896 290382
rect 74033 290170 74099 290173
rect 70678 290168 74099 290170
rect 70678 290112 74038 290168
rect 74094 290112 74099 290168
rect 70678 290110 74099 290112
rect 70678 289596 70738 290110
rect 74033 290107 74099 290110
rect 138014 289354 138020 289356
rect 16717 289082 16783 289085
rect 19894 289082 19954 289324
rect 134710 289294 138020 289354
rect 16717 289080 19954 289082
rect 16717 289024 16722 289080
rect 16778 289024 19954 289080
rect 16717 289022 19954 289024
rect 51309 289082 51375 289085
rect 55038 289082 55098 289256
rect 51309 289080 55098 289082
rect 51309 289024 51314 289080
rect 51370 289024 55098 289080
rect 134710 289052 134770 289294
rect 138014 289292 138020 289294
rect 138084 289292 138090 289356
rect 228726 289292 228732 289356
rect 228796 289292 228802 289356
rect 228734 289082 228794 289292
rect 231077 289082 231143 289085
rect 323118 289082 323124 289084
rect 228734 289080 231143 289082
rect 228734 289052 231082 289080
rect 51309 289022 55098 289024
rect 228764 289024 231082 289052
rect 231138 289024 231143 289080
rect 228764 289022 231143 289024
rect 322788 289022 323124 289082
rect 16717 289019 16783 289022
rect 51309 289019 51375 289022
rect 231077 289019 231143 289022
rect 323118 289020 323124 289022
rect 323188 289020 323194 289084
rect 352750 289082 352810 289256
rect 356197 289082 356263 289085
rect 352750 289080 356263 289082
rect 352750 289024 356202 289080
rect 356258 289024 356263 289080
rect 352750 289022 356263 289024
rect 424694 289082 424754 289256
rect 427221 289082 427287 289085
rect 424694 289080 427287 289082
rect 424694 289024 427226 289080
rect 427282 289024 427287 289080
rect 424694 289022 427287 289024
rect 356197 289019 356263 289022
rect 427221 289019 427287 289022
rect 406061 288674 406127 288677
rect 406061 288672 409114 288674
rect 406061 288616 406066 288672
rect 406122 288616 409114 288672
rect 406061 288614 409114 288616
rect 406061 288611 406127 288614
rect 38797 288130 38863 288133
rect 35748 288128 38863 288130
rect 35748 288072 38802 288128
rect 38858 288072 38863 288128
rect 409054 288100 409114 288614
rect 35748 288070 38863 288072
rect 38797 288067 38863 288070
rect 73430 286300 73436 286364
rect 73500 286362 73506 286364
rect 74166 286362 74172 286364
rect 73500 286302 74172 286362
rect 73500 286300 73506 286302
rect 74166 286300 74172 286302
rect 74236 286300 74242 286364
rect 164702 286362 164762 286808
rect 168057 286362 168123 286365
rect 164702 286360 168123 286362
rect 164702 286304 168062 286360
rect 168118 286304 168123 286360
rect 164702 286302 168123 286304
rect 258726 286362 258786 286808
rect 261253 286362 261319 286365
rect 258726 286360 261319 286362
rect 258726 286304 261258 286360
rect 261314 286304 261319 286360
rect 258726 286302 261319 286304
rect 168057 286299 168123 286302
rect 261253 286299 261319 286302
rect 325285 285954 325351 285957
rect 322788 285952 325351 285954
rect 35718 285546 35778 285584
rect 38797 285546 38863 285549
rect 35718 285544 38863 285546
rect 35718 285488 38802 285544
rect 38858 285488 38863 285544
rect 35718 285486 38863 285488
rect 38797 285483 38863 285486
rect 70862 285410 70922 285924
rect 322788 285896 325290 285952
rect 325346 285896 325351 285952
rect 322788 285894 325351 285896
rect 325285 285891 325351 285894
rect 70862 285350 71106 285410
rect 71046 285002 71106 285350
rect 134710 285274 134770 285856
rect 137605 285274 137671 285277
rect 134710 285272 137671 285274
rect 134710 285216 137610 285272
rect 137666 285216 137671 285272
rect 134710 285214 137671 285216
rect 228734 285274 228794 285856
rect 405969 285546 406035 285549
rect 408870 285546 408930 285652
rect 405969 285544 408930 285546
rect 405969 285488 405974 285544
rect 406030 285488 408930 285544
rect 405969 285486 408930 285488
rect 405969 285483 406035 285486
rect 231353 285274 231419 285277
rect 228734 285272 231419 285274
rect 228734 285216 231358 285272
rect 231414 285216 231419 285272
rect 228734 285214 231419 285216
rect 137605 285211 137671 285214
rect 231353 285211 231419 285214
rect 353662 285212 353668 285276
rect 353732 285274 353738 285276
rect 354265 285274 354331 285277
rect 353732 285272 354331 285274
rect 353732 285216 354270 285272
rect 354326 285216 354331 285272
rect 353732 285214 354331 285216
rect 353732 285212 353738 285214
rect 354265 285211 354331 285214
rect 84654 285002 84660 285004
rect 71046 284942 84660 285002
rect 84654 284940 84660 284942
rect 84724 284940 84730 285004
rect 134886 284804 134892 284868
rect 134956 284866 134962 284868
rect 136869 284866 136935 284869
rect 134956 284864 136935 284866
rect 134956 284808 136874 284864
rect 136930 284808 136935 284864
rect 134956 284806 136935 284808
rect 134956 284804 134962 284806
rect 136869 284803 136935 284806
rect 427681 284322 427747 284325
rect 424724 284320 427747 284322
rect 16533 283506 16599 283509
rect 19894 283506 19954 284292
rect 424724 284264 427686 284320
rect 427742 284264 427747 284320
rect 424724 284262 427747 284264
rect 427681 284259 427747 284262
rect 51493 283778 51559 283781
rect 55038 283778 55098 284224
rect 51493 283776 55098 283778
rect 51493 283720 51498 283776
rect 51554 283720 55098 283776
rect 51493 283718 55098 283720
rect 352750 283778 352810 284224
rect 356197 283778 356263 283781
rect 352750 283776 356263 283778
rect 352750 283720 356202 283776
rect 356258 283720 356263 283776
rect 352750 283718 356263 283720
rect 51493 283715 51559 283718
rect 356197 283715 356263 283718
rect 334209 283642 334275 283645
rect 334209 283640 336956 283642
rect 334209 283584 334214 283640
rect 334270 283584 336956 283640
rect 334209 283582 336956 283584
rect 334209 283579 334275 283582
rect 148326 283514 148908 283574
rect 242350 283514 242932 283574
rect 16533 283504 19954 283506
rect 16533 283448 16538 283504
rect 16594 283448 19954 283504
rect 16533 283446 19954 283448
rect 145149 283506 145215 283509
rect 148326 283506 148386 283514
rect 145149 283504 148386 283506
rect 145149 283448 145154 283504
rect 145210 283448 148386 283504
rect 145149 283446 148386 283448
rect 240369 283506 240435 283509
rect 242350 283506 242410 283514
rect 240369 283504 242410 283506
rect 240369 283448 240374 283504
rect 240430 283448 242410 283504
rect 240369 283446 242410 283448
rect 16533 283443 16599 283446
rect 145149 283443 145215 283446
rect 240369 283443 240435 283446
rect 405969 283370 406035 283373
rect 405969 283368 409114 283370
rect 405969 283312 405974 283368
rect 406030 283312 409114 283368
rect 405969 283310 409114 283312
rect 405969 283307 406035 283310
rect 9896 283098 10376 283128
rect 12669 283098 12735 283101
rect 38061 283098 38127 283101
rect 9896 283096 12735 283098
rect 9896 283040 12674 283096
rect 12730 283040 12735 283096
rect 9896 283038 12735 283040
rect 35748 283096 38127 283098
rect 35748 283040 38066 283096
rect 38122 283040 38127 283096
rect 409054 283068 409114 283310
rect 35748 283038 38127 283040
rect 9896 283008 10376 283038
rect 12669 283035 12735 283038
rect 38061 283035 38127 283038
rect 73614 282826 73620 282828
rect 70678 282766 73620 282826
rect 70678 282252 70738 282766
rect 73614 282764 73620 282766
rect 73684 282826 73690 282828
rect 84470 282826 84476 282828
rect 73684 282766 84476 282826
rect 73684 282764 73690 282766
rect 84470 282764 84476 282766
rect 84540 282764 84546 282828
rect 231629 282826 231695 282829
rect 325837 282826 325903 282829
rect 228764 282824 231695 282826
rect 228764 282768 231634 282824
rect 231690 282768 231695 282824
rect 228764 282766 231695 282768
rect 322788 282824 325903 282826
rect 322788 282768 325842 282824
rect 325898 282768 325903 282824
rect 322788 282766 325903 282768
rect 231629 282763 231695 282766
rect 325837 282763 325903 282766
rect 134710 282554 134770 282728
rect 138157 282554 138223 282557
rect 134710 282552 138223 282554
rect 134710 282496 138162 282552
rect 138218 282496 138223 282552
rect 134710 282494 138223 282496
rect 138157 282491 138223 282494
rect 73430 281948 73436 282012
rect 73500 282010 73506 282012
rect 74166 282010 74172 282012
rect 73500 281950 74172 282010
rect 73500 281948 73506 281950
rect 74166 281948 74172 281950
rect 74236 281948 74242 282012
rect 35718 280378 35778 280552
rect 38061 280378 38127 280381
rect 35718 280376 38127 280378
rect 35718 280320 38066 280376
rect 38122 280320 38127 280376
rect 35718 280318 38127 280320
rect 38061 280315 38127 280318
rect 81669 280242 81735 280245
rect 175417 280242 175483 280245
rect 269257 280242 269323 280245
rect 81669 280240 85060 280242
rect 81669 280184 81674 280240
rect 81730 280184 85060 280240
rect 81669 280182 85060 280184
rect 175417 280240 178900 280242
rect 175417 280184 175422 280240
rect 175478 280184 178900 280240
rect 175417 280182 178900 280184
rect 269257 280240 272924 280242
rect 269257 280184 269262 280240
rect 269318 280184 272924 280240
rect 269257 280182 272924 280184
rect 81669 280179 81735 280182
rect 175417 280179 175483 280182
rect 269257 280179 269323 280182
rect 137697 279698 137763 279701
rect 231445 279698 231511 279701
rect 325377 279698 325443 279701
rect 134740 279696 137763 279698
rect 134740 279640 137702 279696
rect 137758 279640 137763 279696
rect 134740 279638 137763 279640
rect 228764 279696 231511 279698
rect 228764 279640 231450 279696
rect 231506 279640 231511 279696
rect 228764 279638 231511 279640
rect 322788 279696 325443 279698
rect 322788 279640 325382 279696
rect 325438 279640 325443 279696
rect 322788 279638 325443 279640
rect 137697 279635 137763 279638
rect 231445 279635 231511 279638
rect 325377 279635 325443 279638
rect 352742 279636 352748 279700
rect 352812 279698 352818 279700
rect 408870 279698 408930 280620
rect 352812 279638 408930 279698
rect 352812 279636 352818 279638
rect 16717 279426 16783 279429
rect 51493 279426 51559 279429
rect 136869 279426 136935 279429
rect 138382 279426 138388 279428
rect 16717 279424 19770 279426
rect 16717 279368 16722 279424
rect 16778 279368 19770 279424
rect 51493 279424 55068 279426
rect 16717 279366 19770 279368
rect 16717 279363 16783 279366
rect 19710 279290 19770 279366
rect 19894 279290 19954 279396
rect 51493 279368 51498 279424
rect 51554 279368 55068 279424
rect 51493 279366 55068 279368
rect 136869 279424 138388 279426
rect 136869 279368 136874 279424
rect 136930 279368 138388 279424
rect 136869 279366 138388 279368
rect 51493 279363 51559 279366
rect 136869 279363 136935 279366
rect 138382 279364 138388 279366
rect 138452 279364 138458 279428
rect 356197 279426 356263 279429
rect 427865 279426 427931 279429
rect 352780 279424 356263 279426
rect 352780 279368 356202 279424
rect 356258 279368 356263 279424
rect 352780 279366 356263 279368
rect 424724 279424 427931 279426
rect 424724 279368 427870 279424
rect 427926 279368 427931 279424
rect 424724 279366 427931 279368
rect 356197 279363 356263 279366
rect 427865 279363 427931 279366
rect 138433 279292 138499 279293
rect 138382 279290 138388 279292
rect 19710 279230 19954 279290
rect 138342 279230 138388 279290
rect 138452 279288 138499 279292
rect 138494 279232 138499 279288
rect 138382 279228 138388 279230
rect 138452 279228 138499 279232
rect 138433 279227 138499 279228
rect 405969 278746 406035 278749
rect 405969 278744 409114 278746
rect 38613 278202 38679 278205
rect 35748 278200 38679 278202
rect 35748 278144 38618 278200
rect 38674 278144 38679 278200
rect 35748 278142 38679 278144
rect 70862 278202 70922 278716
rect 405969 278688 405974 278744
rect 406030 278688 409114 278744
rect 405969 278686 409114 278688
rect 405969 278683 406035 278686
rect 74033 278202 74099 278205
rect 70862 278200 74099 278202
rect 70862 278144 74038 278200
rect 74094 278144 74099 278200
rect 409054 278172 409114 278686
rect 70862 278142 74099 278144
rect 38613 278139 38679 278142
rect 74033 278139 74099 278142
rect 430257 277930 430323 277933
rect 434416 277930 434896 277960
rect 430257 277928 434896 277930
rect 430257 277872 430262 277928
rect 430318 277872 434896 277928
rect 430257 277870 434896 277872
rect 430257 277867 430323 277870
rect 434416 277840 434896 277870
rect 73430 277324 73436 277388
rect 73500 277386 73506 277388
rect 73500 277326 74234 277386
rect 73500 277324 73506 277326
rect 73430 277188 73436 277252
rect 73500 277250 73506 277252
rect 73982 277250 73988 277252
rect 73500 277190 73988 277250
rect 73500 277188 73506 277190
rect 73982 277188 73988 277190
rect 74052 277188 74058 277252
rect 73982 277052 73988 277116
rect 74052 277114 74058 277116
rect 74174 277114 74234 277326
rect 74052 277054 74234 277114
rect 74052 277052 74058 277054
rect 137789 276570 137855 276573
rect 231537 276570 231603 276573
rect 325469 276570 325535 276573
rect 134740 276568 137855 276570
rect 134740 276512 137794 276568
rect 137850 276512 137855 276568
rect 134740 276510 137855 276512
rect 228764 276568 231603 276570
rect 228764 276512 231542 276568
rect 231598 276512 231603 276568
rect 228764 276510 231603 276512
rect 322788 276568 325535 276570
rect 322788 276512 325474 276568
rect 325530 276512 325535 276568
rect 322788 276510 325535 276512
rect 137789 276507 137855 276510
rect 231537 276507 231603 276510
rect 325469 276507 325535 276510
rect 149054 274876 149060 274940
rect 149124 274938 149130 274940
rect 159041 274938 159107 274941
rect 149124 274936 159107 274938
rect 149124 274880 159046 274936
rect 159102 274880 159107 274936
rect 149124 274878 159107 274880
rect 149124 274876 149130 274878
rect 159041 274875 159107 274878
rect 157753 274802 157819 274805
rect 168926 274802 168932 274804
rect 157753 274800 168932 274802
rect 157753 274744 157758 274800
rect 157814 274744 168932 274800
rect 157753 274742 168932 274744
rect 157753 274739 157819 274742
rect 168926 274740 168932 274742
rect 168996 274740 169002 274804
rect 253157 274802 253223 274805
rect 262030 274802 262036 274804
rect 253157 274800 262036 274802
rect 253157 274744 253162 274800
rect 253218 274744 262036 274800
rect 253157 274742 262036 274744
rect 253157 274739 253223 274742
rect 262030 274740 262036 274742
rect 262100 274740 262106 274804
rect 158397 274666 158463 274669
rect 168558 274666 168564 274668
rect 158397 274664 168564 274666
rect 158397 274608 158402 274664
rect 158458 274608 168564 274664
rect 158397 274606 168564 274608
rect 158397 274603 158463 274606
rect 168558 274604 168564 274606
rect 168628 274604 168634 274668
rect 252697 274666 252763 274669
rect 262398 274666 262404 274668
rect 252697 274664 262404 274666
rect 252697 274608 252702 274664
rect 252758 274608 262404 274664
rect 252697 274606 262404 274608
rect 252697 274603 252763 274606
rect 262398 274604 262404 274606
rect 262468 274604 262474 274668
rect 157201 274530 157267 274533
rect 167822 274530 167828 274532
rect 157201 274528 167828 274530
rect 157201 274472 157206 274528
rect 157262 274472 167828 274528
rect 157201 274470 167828 274472
rect 157201 274467 157267 274470
rect 167822 274468 167828 274470
rect 167892 274468 167898 274532
rect 252053 274530 252119 274533
rect 262582 274530 262588 274532
rect 252053 274528 262588 274530
rect 252053 274472 252058 274528
rect 252114 274472 262588 274528
rect 252053 274470 262588 274472
rect 252053 274467 252119 274470
rect 262582 274468 262588 274470
rect 262652 274468 262658 274532
rect 156557 274394 156623 274397
rect 168190 274394 168196 274396
rect 156557 274392 168196 274394
rect 156557 274336 156562 274392
rect 156618 274336 168196 274392
rect 156557 274334 168196 274336
rect 156557 274331 156623 274334
rect 168190 274332 168196 274334
rect 168260 274332 168266 274396
rect 232733 274394 232799 274397
rect 247269 274394 247335 274397
rect 232733 274392 247335 274394
rect 232733 274336 232738 274392
rect 232794 274336 247274 274392
rect 247330 274336 247335 274392
rect 232733 274334 247335 274336
rect 232733 274331 232799 274334
rect 247269 274331 247335 274334
rect 250857 274394 250923 274397
rect 261662 274394 261668 274396
rect 250857 274392 261668 274394
rect 250857 274336 250862 274392
rect 250918 274336 261668 274392
rect 250857 274334 261668 274336
rect 250857 274331 250923 274334
rect 261662 274332 261668 274334
rect 261732 274332 261738 274396
rect 247821 273988 247887 273989
rect 247821 273984 247868 273988
rect 247932 273986 247938 273988
rect 247821 273928 247826 273984
rect 247821 273924 247868 273928
rect 247932 273926 247978 273986
rect 247932 273924 247938 273926
rect 247821 273923 247887 273924
rect 136910 273788 136916 273852
rect 136980 273850 136986 273852
rect 137513 273850 137579 273853
rect 136980 273848 137579 273850
rect 136980 273792 137518 273848
rect 137574 273792 137579 273848
rect 136980 273790 137579 273792
rect 136980 273788 136986 273790
rect 137513 273787 137579 273790
rect 154574 273788 154580 273852
rect 154644 273850 154650 273852
rect 154717 273850 154783 273853
rect 154644 273848 154783 273850
rect 154644 273792 154722 273848
rect 154778 273792 154783 273848
rect 154644 273790 154783 273792
rect 154644 273788 154650 273790
rect 154717 273787 154783 273790
rect 242342 273788 242348 273852
rect 242412 273850 242418 273852
rect 250949 273850 251015 273853
rect 242412 273848 251015 273850
rect 242412 273792 250954 273848
rect 251010 273792 251015 273848
rect 242412 273790 251015 273792
rect 242412 273788 242418 273790
rect 250949 273787 251015 273790
rect 137881 273442 137947 273445
rect 231629 273442 231695 273445
rect 325561 273442 325627 273445
rect 134740 273440 137947 273442
rect 134740 273384 137886 273440
rect 137942 273384 137947 273440
rect 134740 273382 137947 273384
rect 228764 273440 231695 273442
rect 228764 273384 231634 273440
rect 231690 273384 231695 273440
rect 228764 273382 231695 273384
rect 322788 273440 325627 273442
rect 322788 273384 325566 273440
rect 325622 273384 325627 273440
rect 322788 273382 325627 273384
rect 137881 273379 137947 273382
rect 231629 273379 231695 273382
rect 325561 273379 325627 273382
rect 47077 271674 47143 271677
rect 74217 271674 74283 271677
rect 47077 271672 74283 271674
rect 47077 271616 47082 271672
rect 47138 271616 74222 271672
rect 74278 271616 74283 271672
rect 47077 271614 74283 271616
rect 47077 271611 47143 271614
rect 74217 271611 74283 271614
rect 74217 271132 74283 271133
rect 74166 271068 74172 271132
rect 74236 271130 74283 271132
rect 74236 271128 74328 271130
rect 74278 271072 74328 271128
rect 74236 271070 74328 271072
rect 74236 271068 74283 271070
rect 74217 271067 74283 271068
rect 73982 270388 73988 270452
rect 74052 270450 74058 270452
rect 74052 270390 74234 270450
rect 74052 270388 74058 270390
rect 73430 270252 73436 270316
rect 73500 270314 73506 270316
rect 73982 270314 73988 270316
rect 73500 270254 73988 270314
rect 73500 270252 73506 270254
rect 73982 270252 73988 270254
rect 74052 270252 74058 270316
rect 73430 270116 73436 270180
rect 73500 270178 73506 270180
rect 74174 270178 74234 270390
rect 73500 270118 74234 270178
rect 73500 270116 73506 270118
rect 138433 269906 138499 269909
rect 138566 269906 138572 269908
rect 138433 269904 138572 269906
rect 138433 269848 138438 269904
rect 138494 269848 138572 269904
rect 138433 269846 138572 269848
rect 138433 269843 138499 269846
rect 138566 269844 138572 269846
rect 138636 269844 138642 269908
rect 9896 269770 10376 269800
rect 12853 269770 12919 269773
rect 9896 269768 12919 269770
rect 9896 269712 12858 269768
rect 12914 269712 12919 269768
rect 9896 269710 12919 269712
rect 9896 269680 10376 269710
rect 12853 269707 12919 269710
rect 138566 269572 138572 269636
rect 138636 269634 138642 269636
rect 138750 269634 138756 269636
rect 138636 269574 138756 269634
rect 138636 269572 138642 269574
rect 138750 269572 138756 269574
rect 138820 269572 138826 269636
rect 182961 269500 183027 269501
rect 182910 269498 182916 269500
rect 182870 269438 182916 269498
rect 182980 269496 183027 269500
rect 183022 269440 183027 269496
rect 182910 269436 182916 269438
rect 182980 269436 183027 269440
rect 182961 269435 183027 269436
rect 218013 268410 218079 268413
rect 219710 268410 219716 268412
rect 218013 268408 219716 268410
rect 218013 268352 218018 268408
rect 218074 268352 219716 268408
rect 218013 268350 219716 268352
rect 218013 268347 218079 268350
rect 219710 268348 219716 268350
rect 219780 268348 219786 268412
rect 351822 266716 351828 266780
rect 351892 266778 351898 266780
rect 352057 266778 352123 266781
rect 351892 266776 352123 266778
rect 351892 266720 352062 266776
rect 352118 266720 352123 266776
rect 351892 266718 352123 266720
rect 351892 266716 351898 266718
rect 352057 266715 352123 266718
rect 55214 266580 55220 266644
rect 55284 266642 55290 266644
rect 55541 266642 55607 266645
rect 55284 266640 55607 266642
rect 55284 266584 55546 266640
rect 55602 266584 55607 266640
rect 55284 266582 55607 266584
rect 55284 266580 55290 266582
rect 55541 266579 55607 266582
rect 350953 266642 351019 266645
rect 352006 266642 352012 266644
rect 350953 266640 352012 266642
rect 350953 266584 350958 266640
rect 351014 266584 352012 266640
rect 350953 266582 352012 266584
rect 350953 266579 351019 266582
rect 352006 266580 352012 266582
rect 352076 266580 352082 266644
rect 52638 265492 52644 265556
rect 52708 265554 52714 265556
rect 53517 265554 53583 265557
rect 52708 265552 53583 265554
rect 52708 265496 53522 265552
rect 53578 265496 53583 265552
rect 52708 265494 53583 265496
rect 52708 265492 52714 265494
rect 53517 265491 53583 265494
rect 54529 265554 54595 265557
rect 54662 265554 54668 265556
rect 54529 265552 54668 265554
rect 54529 265496 54534 265552
rect 54590 265496 54668 265552
rect 54529 265494 54668 265496
rect 54529 265491 54595 265494
rect 54662 265492 54668 265494
rect 54732 265492 54738 265556
rect 55398 265492 55404 265556
rect 55468 265554 55474 265556
rect 56553 265554 56619 265557
rect 55468 265552 56619 265554
rect 55468 265496 56558 265552
rect 56614 265496 56619 265552
rect 55468 265494 56619 265496
rect 55468 265492 55474 265494
rect 56553 265491 56619 265494
rect 429429 265418 429495 265421
rect 434416 265418 434896 265448
rect 429429 265416 434896 265418
rect 429429 265360 429434 265416
rect 429490 265360 434896 265416
rect 429429 265358 434896 265360
rect 429429 265355 429495 265358
rect 434416 265328 434896 265358
rect 241422 263860 241428 263924
rect 241492 263922 241498 263924
rect 242710 263922 242716 263924
rect 241492 263862 242716 263922
rect 241492 263860 241498 263862
rect 242710 263860 242716 263862
rect 242780 263860 242786 263924
rect 73798 263588 73804 263652
rect 73868 263650 73874 263652
rect 75454 263650 75460 263652
rect 73868 263590 75460 263650
rect 73868 263588 73874 263590
rect 75454 263588 75460 263590
rect 75524 263588 75530 263652
rect 78909 263650 78975 263653
rect 76750 263648 78975 263650
rect 76750 263592 78914 263648
rect 78970 263592 78975 263648
rect 76750 263590 78975 263592
rect 73941 263514 74007 263517
rect 74534 263514 74540 263516
rect 73941 263512 74540 263514
rect 73941 263456 73946 263512
rect 74002 263456 74540 263512
rect 73941 263454 74540 263456
rect 73941 263451 74007 263454
rect 74534 263452 74540 263454
rect 74604 263452 74610 263516
rect 73430 263316 73436 263380
rect 73500 263378 73506 263380
rect 74718 263378 74724 263380
rect 73500 263318 74724 263378
rect 73500 263316 73506 263318
rect 74718 263316 74724 263318
rect 74788 263316 74794 263380
rect 76750 263144 76810 263590
rect 78909 263587 78975 263590
rect 245102 263452 245108 263516
rect 245172 263514 245178 263516
rect 251174 263514 251180 263516
rect 245172 263454 251180 263514
rect 245172 263452 245178 263454
rect 251174 263452 251180 263454
rect 251244 263452 251250 263516
rect 328413 263514 328479 263517
rect 328413 263512 331098 263514
rect 328413 263456 328418 263512
rect 328474 263456 331098 263512
rect 328413 263454 331098 263456
rect 328413 263451 328479 263454
rect 331038 263144 331098 263454
rect 139813 263106 139879 263109
rect 173485 263106 173551 263109
rect 139813 263104 143020 263106
rect 139813 263048 139818 263104
rect 139874 263048 143020 263104
rect 139813 263046 143020 263048
rect 170804 263104 173551 263106
rect 170804 263048 173490 263104
rect 173546 263048 173551 263104
rect 170804 263046 173551 263048
rect 139813 263043 139879 263046
rect 173485 263043 173551 263046
rect 233469 263106 233535 263109
rect 267417 263106 267483 263109
rect 233469 263104 237044 263106
rect 233469 263048 233474 263104
rect 233530 263048 237044 263104
rect 233469 263046 237044 263048
rect 264828 263104 267483 263106
rect 264828 263048 267422 263104
rect 267478 263048 267483 263104
rect 264828 263046 267483 263048
rect 233469 263043 233535 263046
rect 267417 263043 267483 263046
rect 49193 262698 49259 262701
rect 49150 262696 49259 262698
rect 49150 262640 49198 262696
rect 49254 262640 49259 262696
rect 49150 262635 49259 262640
rect 49150 262260 49210 262635
rect 360797 262290 360863 262293
rect 358852 262288 360863 262290
rect 358852 262232 360802 262288
rect 360858 262232 360863 262288
rect 358852 262230 360863 262232
rect 360797 262227 360863 262230
rect 183830 262092 183836 262156
rect 183900 262154 183906 262156
rect 193214 262154 193220 262156
rect 183900 262094 193220 262154
rect 183900 262092 183906 262094
rect 193214 262092 193220 262094
rect 193284 262092 193290 262156
rect 78909 261746 78975 261749
rect 76780 261744 78975 261746
rect 76780 261688 78914 261744
rect 78970 261688 78975 261744
rect 76780 261686 78975 261688
rect 78909 261683 78975 261686
rect 140365 261746 140431 261749
rect 173393 261746 173459 261749
rect 140365 261744 143020 261746
rect 140365 261688 140370 261744
rect 140426 261688 143020 261744
rect 140365 261686 143020 261688
rect 170804 261744 173459 261746
rect 170804 261688 173398 261744
rect 173454 261688 173459 261744
rect 170804 261686 173459 261688
rect 140365 261683 140431 261686
rect 173393 261683 173459 261686
rect 233469 261746 233535 261749
rect 267509 261746 267575 261749
rect 233469 261744 237044 261746
rect 233469 261688 233474 261744
rect 233530 261688 237044 261744
rect 233469 261686 237044 261688
rect 264828 261744 267575 261746
rect 264828 261688 267514 261744
rect 267570 261688 267575 261744
rect 264828 261686 267575 261688
rect 233469 261683 233535 261686
rect 267509 261683 267575 261686
rect 327677 261746 327743 261749
rect 327677 261744 331068 261746
rect 327677 261688 327682 261744
rect 327738 261688 331068 261744
rect 327677 261686 331068 261688
rect 327677 261683 327743 261686
rect 278958 261412 278964 261476
rect 279028 261474 279034 261476
rect 288526 261474 288532 261476
rect 279028 261414 288532 261474
rect 279028 261412 279034 261414
rect 288526 261412 288532 261414
rect 288596 261412 288602 261476
rect 298278 261412 298284 261476
rect 298348 261474 298354 261476
rect 307846 261474 307852 261476
rect 298348 261414 307852 261474
rect 298348 261412 298354 261414
rect 307846 261412 307852 261414
rect 307916 261412 307922 261476
rect 317598 261412 317604 261476
rect 317668 261474 317674 261476
rect 327166 261474 327172 261476
rect 317668 261414 327172 261474
rect 317668 261412 317674 261414
rect 327166 261412 327172 261414
rect 327236 261412 327242 261476
rect 203150 260732 203156 260796
rect 203220 260794 203226 260796
rect 212534 260794 212540 260796
rect 203220 260734 212540 260794
rect 203220 260732 203226 260734
rect 212534 260732 212540 260734
rect 212604 260732 212610 260796
rect 78909 260386 78975 260389
rect 76780 260384 78975 260386
rect 76780 260328 78914 260384
rect 78970 260328 78975 260384
rect 76780 260326 78975 260328
rect 78909 260323 78975 260326
rect 140365 260386 140431 260389
rect 173761 260386 173827 260389
rect 140365 260384 143020 260386
rect 140365 260328 140370 260384
rect 140426 260328 143020 260384
rect 140365 260326 143020 260328
rect 170804 260384 173827 260386
rect 170804 260328 173766 260384
rect 173822 260328 173827 260384
rect 170804 260326 173827 260328
rect 140365 260323 140431 260326
rect 173761 260323 173827 260326
rect 233469 260386 233535 260389
rect 267601 260386 267667 260389
rect 233469 260384 237044 260386
rect 233469 260328 233474 260384
rect 233530 260328 237044 260384
rect 233469 260326 237044 260328
rect 264828 260384 267667 260386
rect 264828 260328 267606 260384
rect 267662 260328 267667 260384
rect 264828 260326 267667 260328
rect 233469 260323 233535 260326
rect 267601 260323 267667 260326
rect 327953 260386 328019 260389
rect 327953 260384 331068 260386
rect 327953 260328 327958 260384
rect 328014 260328 331068 260384
rect 327953 260326 331068 260328
rect 327953 260323 328019 260326
rect 138801 259980 138867 259981
rect 138750 259916 138756 259980
rect 138820 259978 138867 259980
rect 138820 259976 138912 259978
rect 138862 259920 138912 259976
rect 138820 259918 138912 259920
rect 138820 259916 138867 259918
rect 138801 259915 138867 259916
rect 48958 259372 48964 259436
rect 49028 259372 49034 259436
rect 46617 259162 46683 259165
rect 48966 259162 49026 259372
rect 360613 259162 360679 259165
rect 46617 259160 49026 259162
rect 46617 259104 46622 259160
rect 46678 259132 49026 259160
rect 358852 259160 360679 259162
rect 46678 259104 48996 259132
rect 46617 259102 48996 259104
rect 358852 259104 360618 259160
rect 360674 259104 360679 259160
rect 358852 259102 360679 259104
rect 46617 259099 46683 259102
rect 360613 259099 360679 259102
rect 78909 258890 78975 258893
rect 76780 258888 78975 258890
rect 76780 258832 78914 258888
rect 78970 258832 78975 258888
rect 76780 258830 78975 258832
rect 78909 258827 78975 258830
rect 140549 258890 140615 258893
rect 173853 258890 173919 258893
rect 140549 258888 143020 258890
rect 140549 258832 140554 258888
rect 140610 258832 143020 258888
rect 140549 258830 143020 258832
rect 170804 258888 173919 258890
rect 170804 258832 173858 258888
rect 173914 258832 173919 258888
rect 170804 258830 173919 258832
rect 140549 258827 140615 258830
rect 173853 258827 173919 258830
rect 233469 258890 233535 258893
rect 267325 258890 267391 258893
rect 233469 258888 237044 258890
rect 233469 258832 233474 258888
rect 233530 258832 237044 258888
rect 233469 258830 237044 258832
rect 264828 258888 267391 258890
rect 264828 258832 267330 258888
rect 267386 258832 267391 258888
rect 264828 258830 267391 258832
rect 233469 258827 233535 258830
rect 267325 258827 267391 258830
rect 327217 258890 327283 258893
rect 327217 258888 331068 258890
rect 327217 258832 327222 258888
rect 327278 258832 331068 258888
rect 327217 258830 331068 258832
rect 327217 258827 327283 258830
rect 87189 258074 87255 258077
rect 87189 258072 90058 258074
rect 87189 258016 87194 258072
rect 87250 258016 90058 258072
rect 87189 258014 90058 258016
rect 87189 258011 87255 258014
rect 78909 257530 78975 257533
rect 76780 257528 78975 257530
rect 76780 257472 78914 257528
rect 78970 257472 78975 257528
rect 76780 257470 78975 257472
rect 78909 257467 78975 257470
rect 89998 257432 90058 258014
rect 140549 257530 140615 257533
rect 173669 257530 173735 257533
rect 140549 257528 143020 257530
rect 140549 257472 140554 257528
rect 140610 257472 143020 257528
rect 140549 257470 143020 257472
rect 170804 257528 173735 257530
rect 170804 257472 173674 257528
rect 173730 257472 173735 257528
rect 170804 257470 173735 257472
rect 140549 257467 140615 257470
rect 173669 257467 173735 257470
rect 233469 257530 233535 257533
rect 267785 257530 267851 257533
rect 233469 257528 237044 257530
rect 233469 257472 233474 257528
rect 233530 257472 237044 257528
rect 233469 257470 237044 257472
rect 264828 257528 267851 257530
rect 264828 257472 267790 257528
rect 267846 257472 267851 257528
rect 264828 257470 267851 257472
rect 233469 257467 233535 257470
rect 267785 257467 267851 257470
rect 327125 257530 327191 257533
rect 327125 257528 331068 257530
rect 327125 257472 327130 257528
rect 327186 257472 331068 257528
rect 327125 257470 331068 257472
rect 327125 257467 327191 257470
rect 131349 257394 131415 257397
rect 129772 257392 131415 257394
rect 129772 257336 131354 257392
rect 131410 257336 131415 257392
rect 129772 257334 131415 257336
rect 131349 257331 131415 257334
rect 181029 257394 181095 257397
rect 226477 257394 226543 257397
rect 181029 257392 184052 257394
rect 181029 257336 181034 257392
rect 181090 257336 184052 257392
rect 181029 257334 184052 257336
rect 223796 257392 226543 257394
rect 223796 257336 226482 257392
rect 226538 257336 226543 257392
rect 223796 257334 226543 257336
rect 181029 257331 181095 257334
rect 226477 257331 226543 257334
rect 276157 257394 276223 257397
rect 321053 257394 321119 257397
rect 276157 257392 278076 257394
rect 276157 257336 276162 257392
rect 276218 257336 278076 257392
rect 276157 257334 278076 257336
rect 317820 257392 321119 257394
rect 317820 257336 321058 257392
rect 321114 257336 321119 257392
rect 317820 257334 321119 257336
rect 276157 257331 276223 257334
rect 321053 257331 321119 257334
rect 87189 256850 87255 256853
rect 87189 256848 90058 256850
rect 87189 256792 87194 256848
rect 87250 256792 90058 256848
rect 87189 256790 90058 256792
rect 87189 256787 87255 256790
rect 89998 256480 90058 256790
rect 132361 256442 132427 256445
rect 129772 256440 132427 256442
rect 129772 256384 132366 256440
rect 132422 256384 132427 256440
rect 129772 256382 132427 256384
rect 132361 256379 132427 256382
rect 181029 256442 181095 256445
rect 226477 256442 226543 256445
rect 181029 256440 184052 256442
rect 181029 256384 181034 256440
rect 181090 256384 184052 256440
rect 181029 256382 184052 256384
rect 223796 256440 226543 256442
rect 223796 256384 226482 256440
rect 226538 256384 226543 256440
rect 223796 256382 226543 256384
rect 181029 256379 181095 256382
rect 226477 256379 226543 256382
rect 274961 256442 275027 256445
rect 321053 256442 321119 256445
rect 274961 256440 278076 256442
rect 274961 256384 274966 256440
rect 275022 256384 278076 256440
rect 274961 256382 278076 256384
rect 317820 256440 321119 256442
rect 317820 256384 321058 256440
rect 321114 256384 321119 256440
rect 317820 256382 321119 256384
rect 274961 256379 275027 256382
rect 321053 256379 321119 256382
rect 9896 256306 10376 256336
rect 12853 256306 12919 256309
rect 9896 256304 12919 256306
rect 9896 256248 12858 256304
rect 12914 256248 12919 256304
rect 9896 256246 12919 256248
rect 9896 256216 10376 256246
rect 12853 256243 12919 256246
rect 78909 256170 78975 256173
rect 76780 256168 78975 256170
rect 76780 256112 78914 256168
rect 78970 256112 78975 256168
rect 76780 256110 78975 256112
rect 78909 256107 78975 256110
rect 140457 256170 140523 256173
rect 173301 256170 173367 256173
rect 140457 256168 143020 256170
rect 140457 256112 140462 256168
rect 140518 256112 143020 256168
rect 140457 256110 143020 256112
rect 170804 256168 173367 256170
rect 170804 256112 173306 256168
rect 173362 256112 173367 256168
rect 170804 256110 173367 256112
rect 140457 256107 140523 256110
rect 173301 256107 173367 256110
rect 233469 256170 233535 256173
rect 266589 256170 266655 256173
rect 233469 256168 237044 256170
rect 233469 256112 233474 256168
rect 233530 256112 237044 256168
rect 233469 256110 237044 256112
rect 264828 256168 266655 256170
rect 264828 256112 266594 256168
rect 266650 256112 266655 256168
rect 264828 256110 266655 256112
rect 233469 256107 233535 256110
rect 266589 256107 266655 256110
rect 328505 256170 328571 256173
rect 328505 256168 331068 256170
rect 328505 256112 328510 256168
rect 328566 256112 331068 256168
rect 328505 256110 331068 256112
rect 328505 256107 328571 256110
rect 46525 256034 46591 256037
rect 360521 256034 360587 256037
rect 361165 256034 361231 256037
rect 46525 256032 48996 256034
rect 46525 255976 46530 256032
rect 46586 256004 48996 256032
rect 358852 256032 361231 256034
rect 46586 255976 49026 256004
rect 46525 255974 49026 255976
rect 358852 255976 360526 256032
rect 360582 255976 361170 256032
rect 361226 255976 361231 256032
rect 358852 255974 361231 255976
rect 46525 255971 46591 255974
rect 48966 255900 49026 255974
rect 360521 255971 360587 255974
rect 361165 255971 361231 255974
rect 48958 255836 48964 255900
rect 49028 255836 49034 255900
rect 87281 255626 87347 255629
rect 131993 255626 132059 255629
rect 87281 255624 90028 255626
rect 87281 255568 87286 255624
rect 87342 255568 90028 255624
rect 87281 255566 90028 255568
rect 129772 255624 132059 255626
rect 129772 255568 131998 255624
rect 132054 255568 132059 255624
rect 129772 255566 132059 255568
rect 87281 255563 87347 255566
rect 131993 255563 132059 255566
rect 181581 255626 181647 255629
rect 225925 255626 225991 255629
rect 181581 255624 184052 255626
rect 181581 255568 181586 255624
rect 181642 255568 184052 255624
rect 181581 255566 184052 255568
rect 223796 255624 225991 255626
rect 223796 255568 225930 255624
rect 225986 255568 225991 255624
rect 223796 255566 225991 255568
rect 181581 255563 181647 255566
rect 225925 255563 225991 255566
rect 274869 255626 274935 255629
rect 321605 255626 321671 255629
rect 274869 255624 278076 255626
rect 274869 255568 274874 255624
rect 274930 255568 278076 255624
rect 274869 255566 278076 255568
rect 317820 255624 321671 255626
rect 317820 255568 321610 255624
rect 321666 255568 321671 255624
rect 317820 255566 321671 255568
rect 274869 255563 274935 255566
rect 321605 255563 321671 255566
rect 87189 255354 87255 255357
rect 87189 255352 90058 255354
rect 87189 255296 87194 255352
rect 87250 255296 90058 255352
rect 87189 255294 90058 255296
rect 87189 255291 87255 255294
rect 89998 254712 90058 255294
rect 78909 254674 78975 254677
rect 131349 254674 131415 254677
rect 76780 254672 78975 254674
rect 76780 254616 78914 254672
rect 78970 254616 78975 254672
rect 76780 254614 78975 254616
rect 129772 254672 131415 254674
rect 129772 254616 131354 254672
rect 131410 254616 131415 254672
rect 129772 254614 131415 254616
rect 78909 254611 78975 254614
rect 131349 254611 131415 254614
rect 140549 254674 140615 254677
rect 173301 254674 173367 254677
rect 140549 254672 143020 254674
rect 140549 254616 140554 254672
rect 140610 254616 143020 254672
rect 140549 254614 143020 254616
rect 170804 254672 173367 254674
rect 170804 254616 173306 254672
rect 173362 254616 173367 254672
rect 170804 254614 173367 254616
rect 140549 254611 140615 254614
rect 173301 254611 173367 254614
rect 181029 254674 181095 254677
rect 226385 254674 226451 254677
rect 181029 254672 184052 254674
rect 181029 254616 181034 254672
rect 181090 254616 184052 254672
rect 181029 254614 184052 254616
rect 223796 254672 226451 254674
rect 223796 254616 226390 254672
rect 226446 254616 226451 254672
rect 223796 254614 226451 254616
rect 181029 254611 181095 254614
rect 226385 254611 226451 254614
rect 232733 254674 232799 254677
rect 266589 254674 266655 254677
rect 232733 254672 237044 254674
rect 232733 254616 232738 254672
rect 232794 254616 237044 254672
rect 232733 254614 237044 254616
rect 264828 254672 266655 254674
rect 264828 254616 266594 254672
rect 266650 254616 266655 254672
rect 264828 254614 266655 254616
rect 232733 254611 232799 254614
rect 266589 254611 266655 254614
rect 275789 254674 275855 254677
rect 320593 254674 320659 254677
rect 275789 254672 278076 254674
rect 275789 254616 275794 254672
rect 275850 254616 278076 254672
rect 275789 254614 278076 254616
rect 317820 254672 320659 254674
rect 317820 254616 320598 254672
rect 320654 254616 320659 254672
rect 317820 254614 320659 254616
rect 275789 254611 275855 254614
rect 320593 254611 320659 254614
rect 328413 254674 328479 254677
rect 328413 254672 331068 254674
rect 328413 254616 328418 254672
rect 328474 254616 331068 254672
rect 328413 254614 331068 254616
rect 328413 254611 328479 254614
rect 87189 254402 87255 254405
rect 87189 254400 90058 254402
rect 87189 254344 87194 254400
rect 87250 254344 90058 254400
rect 87189 254342 90058 254344
rect 87189 254339 87255 254342
rect 89998 253896 90058 254342
rect 131349 253858 131415 253861
rect 129772 253856 131415 253858
rect 129772 253800 131354 253856
rect 131410 253800 131415 253856
rect 129772 253798 131415 253800
rect 131349 253795 131415 253798
rect 181029 253858 181095 253861
rect 225741 253858 225807 253861
rect 181029 253856 184052 253858
rect 181029 253800 181034 253856
rect 181090 253800 184052 253856
rect 181029 253798 184052 253800
rect 223796 253856 225807 253858
rect 223796 253800 225746 253856
rect 225802 253800 225807 253856
rect 223796 253798 225807 253800
rect 181029 253795 181095 253798
rect 225741 253795 225807 253798
rect 275881 253858 275947 253861
rect 321605 253858 321671 253861
rect 275881 253856 278076 253858
rect 275881 253800 275886 253856
rect 275942 253800 278076 253856
rect 275881 253798 278076 253800
rect 317820 253856 321671 253858
rect 317820 253800 321610 253856
rect 321666 253800 321671 253856
rect 317820 253798 321671 253800
rect 275881 253795 275947 253798
rect 321605 253795 321671 253798
rect 78909 253314 78975 253317
rect 76780 253312 78975 253314
rect 76780 253256 78914 253312
rect 78970 253256 78975 253312
rect 76780 253254 78975 253256
rect 78909 253251 78975 253254
rect 139813 253314 139879 253317
rect 173945 253314 174011 253317
rect 139813 253312 143020 253314
rect 139813 253256 139818 253312
rect 139874 253256 143020 253312
rect 139813 253254 143020 253256
rect 170804 253312 174011 253314
rect 170804 253256 173950 253312
rect 174006 253256 174011 253312
rect 170804 253254 174011 253256
rect 139813 253251 139879 253254
rect 173945 253251 174011 253254
rect 233469 253314 233535 253317
rect 266589 253314 266655 253317
rect 233469 253312 237044 253314
rect 233469 253256 233474 253312
rect 233530 253256 237044 253312
rect 233469 253254 237044 253256
rect 264828 253312 266655 253314
rect 264828 253256 266594 253312
rect 266650 253256 266655 253312
rect 264828 253254 266655 253256
rect 233469 253251 233535 253254
rect 266589 253251 266655 253254
rect 327125 253314 327191 253317
rect 327125 253312 331068 253314
rect 327125 253256 327130 253312
rect 327186 253256 331068 253312
rect 327125 253254 331068 253256
rect 327125 253251 327191 253254
rect 47077 252906 47143 252909
rect 87189 252906 87255 252909
rect 131349 252906 131415 252909
rect 47077 252904 48996 252906
rect 47077 252848 47082 252904
rect 47138 252848 48996 252904
rect 47077 252846 48996 252848
rect 87189 252904 90028 252906
rect 87189 252848 87194 252904
rect 87250 252848 90028 252904
rect 87189 252846 90028 252848
rect 129772 252904 131415 252906
rect 129772 252848 131354 252904
rect 131410 252848 131415 252904
rect 129772 252846 131415 252848
rect 47077 252843 47143 252846
rect 87189 252843 87255 252846
rect 131349 252843 131415 252846
rect 181581 252906 181647 252909
rect 226477 252906 226543 252909
rect 181581 252904 184052 252906
rect 181581 252848 181586 252904
rect 181642 252848 184052 252904
rect 181581 252846 184052 252848
rect 223796 252904 226543 252906
rect 223796 252848 226482 252904
rect 226538 252848 226543 252904
rect 223796 252846 226543 252848
rect 181581 252843 181647 252846
rect 226477 252843 226543 252846
rect 274869 252906 274935 252909
rect 320501 252906 320567 252909
rect 360705 252906 360771 252909
rect 361165 252906 361231 252909
rect 274869 252904 278076 252906
rect 274869 252848 274874 252904
rect 274930 252848 278076 252904
rect 274869 252846 278076 252848
rect 317820 252904 320567 252906
rect 317820 252848 320506 252904
rect 320562 252848 320567 252904
rect 317820 252846 320567 252848
rect 358852 252904 361231 252906
rect 358852 252848 360710 252904
rect 360766 252848 361170 252904
rect 361226 252848 361231 252904
rect 358852 252846 361231 252848
rect 274869 252843 274935 252846
rect 320501 252843 320567 252846
rect 360705 252843 360771 252846
rect 361165 252843 361231 252846
rect 429429 252906 429495 252909
rect 434416 252906 434896 252936
rect 429429 252904 434896 252906
rect 429429 252848 429434 252904
rect 429490 252848 434896 252904
rect 429429 252846 434896 252848
rect 429429 252843 429495 252846
rect 434416 252816 434896 252846
rect 87281 252770 87347 252773
rect 87281 252768 90058 252770
rect 87281 252712 87286 252768
rect 87342 252712 90058 252768
rect 87281 252710 90058 252712
rect 87281 252707 87347 252710
rect 89998 252128 90058 252710
rect 133373 252090 133439 252093
rect 129772 252088 133439 252090
rect 129772 252032 133378 252088
rect 133434 252032 133439 252088
rect 129772 252030 133439 252032
rect 133373 252027 133439 252030
rect 181673 252090 181739 252093
rect 227213 252090 227279 252093
rect 181673 252088 184052 252090
rect 181673 252032 181678 252088
rect 181734 252032 184052 252088
rect 181673 252030 184052 252032
rect 223796 252088 227279 252090
rect 223796 252032 227218 252088
rect 227274 252032 227279 252088
rect 223796 252030 227279 252032
rect 181673 252027 181739 252030
rect 227213 252027 227279 252030
rect 275605 252090 275671 252093
rect 321605 252090 321671 252093
rect 275605 252088 278076 252090
rect 275605 252032 275610 252088
rect 275666 252032 278076 252088
rect 275605 252030 278076 252032
rect 317820 252088 321671 252090
rect 317820 252032 321610 252088
rect 321666 252032 321671 252088
rect 317820 252030 321671 252032
rect 275605 252027 275671 252030
rect 321605 252027 321671 252030
rect 78909 251954 78975 251957
rect 76780 251952 78975 251954
rect 76780 251896 78914 251952
rect 78970 251896 78975 251952
rect 76780 251894 78975 251896
rect 78909 251891 78975 251894
rect 140549 251954 140615 251957
rect 174037 251954 174103 251957
rect 140549 251952 143020 251954
rect 140549 251896 140554 251952
rect 140610 251896 143020 251952
rect 140549 251894 143020 251896
rect 170804 251952 174103 251954
rect 170804 251896 174042 251952
rect 174098 251896 174103 251952
rect 170804 251894 174103 251896
rect 140549 251891 140615 251894
rect 174037 251891 174103 251894
rect 233561 251954 233627 251957
rect 266589 251954 266655 251957
rect 233561 251952 237044 251954
rect 233561 251896 233566 251952
rect 233622 251896 237044 251952
rect 233561 251894 237044 251896
rect 264828 251952 266655 251954
rect 264828 251896 266594 251952
rect 266650 251896 266655 251952
rect 264828 251894 266655 251896
rect 233561 251891 233627 251894
rect 266589 251891 266655 251894
rect 327217 251954 327283 251957
rect 327217 251952 331068 251954
rect 327217 251896 327222 251952
rect 327278 251896 331068 251952
rect 327217 251894 331068 251896
rect 327217 251891 327283 251894
rect 87189 251546 87255 251549
rect 87189 251544 90058 251546
rect 87189 251488 87194 251544
rect 87250 251488 90058 251544
rect 87189 251486 90058 251488
rect 87189 251483 87255 251486
rect 89998 251176 90058 251486
rect 132177 251138 132243 251141
rect 129772 251136 132243 251138
rect 129772 251080 132182 251136
rect 132238 251080 132243 251136
rect 129772 251078 132243 251080
rect 132177 251075 132243 251078
rect 182317 251138 182383 251141
rect 226017 251138 226083 251141
rect 182317 251136 184052 251138
rect 182317 251080 182322 251136
rect 182378 251080 184052 251136
rect 182317 251078 184052 251080
rect 223796 251136 226083 251138
rect 223796 251080 226022 251136
rect 226078 251080 226083 251136
rect 223796 251078 226083 251080
rect 182317 251075 182383 251078
rect 226017 251075 226083 251078
rect 275513 251138 275579 251141
rect 321605 251138 321671 251141
rect 275513 251136 278076 251138
rect 275513 251080 275518 251136
rect 275574 251080 278076 251136
rect 275513 251078 278076 251080
rect 317820 251136 321671 251138
rect 317820 251080 321610 251136
rect 321666 251080 321671 251136
rect 317820 251078 321671 251080
rect 275513 251075 275579 251078
rect 321605 251075 321671 251078
rect 233469 251002 233535 251005
rect 233469 251000 237074 251002
rect 233469 250944 233474 251000
rect 233530 250944 237074 251000
rect 233469 250942 237074 250944
rect 233469 250939 233535 250942
rect 237014 250632 237074 250942
rect 79737 250594 79803 250597
rect 138801 250594 138867 250597
rect 76780 250592 79803 250594
rect 76780 250536 79742 250592
rect 79798 250536 79803 250592
rect 76780 250534 79803 250536
rect 79737 250531 79803 250534
rect 138758 250592 138867 250594
rect 138758 250536 138806 250592
rect 138862 250536 138867 250592
rect 138758 250531 138867 250536
rect 140733 250594 140799 250597
rect 173577 250594 173643 250597
rect 267325 250594 267391 250597
rect 140733 250592 143020 250594
rect 140733 250536 140738 250592
rect 140794 250536 143020 250592
rect 140733 250534 143020 250536
rect 170804 250592 173643 250594
rect 170804 250536 173582 250592
rect 173638 250536 173643 250592
rect 170804 250534 173643 250536
rect 264828 250592 267391 250594
rect 264828 250536 267330 250592
rect 267386 250536 267391 250592
rect 264828 250534 267391 250536
rect 140733 250531 140799 250534
rect 173577 250531 173643 250534
rect 267325 250531 267391 250534
rect 327217 250594 327283 250597
rect 327217 250592 331068 250594
rect 327217 250536 327222 250592
rect 327278 250536 331068 250592
rect 327217 250534 331068 250536
rect 327217 250531 327283 250534
rect 138758 250460 138818 250531
rect 138750 250396 138756 250460
rect 138820 250396 138826 250460
rect 87189 250322 87255 250325
rect 131993 250322 132059 250325
rect 87189 250320 90028 250322
rect 87189 250264 87194 250320
rect 87250 250264 90028 250320
rect 87189 250262 90028 250264
rect 129772 250320 132059 250322
rect 129772 250264 131998 250320
rect 132054 250264 132059 250320
rect 129772 250262 132059 250264
rect 87189 250259 87255 250262
rect 131993 250259 132059 250262
rect 181765 250322 181831 250325
rect 225833 250322 225899 250325
rect 181765 250320 184052 250322
rect 181765 250264 181770 250320
rect 181826 250264 184052 250320
rect 181765 250262 184052 250264
rect 223796 250320 225899 250322
rect 223796 250264 225838 250320
rect 225894 250264 225899 250320
rect 223796 250262 225899 250264
rect 181765 250259 181831 250262
rect 225833 250259 225899 250262
rect 275697 250322 275763 250325
rect 321053 250322 321119 250325
rect 275697 250320 278076 250322
rect 275697 250264 275702 250320
rect 275758 250264 278076 250320
rect 275697 250262 278076 250264
rect 317820 250320 321119 250322
rect 317820 250264 321058 250320
rect 321114 250264 321119 250320
rect 317820 250262 321119 250264
rect 275697 250259 275763 250262
rect 321053 250259 321119 250262
rect 131809 250050 131875 250053
rect 129742 250048 131875 250050
rect 129742 249992 131814 250048
rect 131870 249992 131875 250048
rect 129742 249990 131875 249992
rect 46433 249778 46499 249781
rect 46433 249776 48996 249778
rect 46433 249720 46438 249776
rect 46494 249748 48996 249776
rect 46494 249720 49026 249748
rect 46433 249718 49026 249720
rect 46433 249715 46499 249718
rect 48966 249236 49026 249718
rect 129742 249408 129802 249990
rect 131809 249987 131875 249990
rect 274869 250050 274935 250053
rect 274869 250048 278106 250050
rect 274869 249992 274874 250048
rect 274930 249992 278106 250048
rect 274869 249990 278106 249992
rect 274869 249987 274935 249990
rect 140641 249778 140707 249781
rect 181489 249778 181555 249781
rect 232825 249778 232891 249781
rect 140641 249776 143050 249778
rect 140641 249720 140646 249776
rect 140702 249720 143050 249776
rect 140641 249718 143050 249720
rect 140641 249715 140707 249718
rect 78909 249370 78975 249373
rect 76750 249368 78975 249370
rect 76750 249312 78914 249368
rect 78970 249312 78975 249368
rect 76750 249310 78975 249312
rect 48958 249172 48964 249236
rect 49028 249172 49034 249236
rect 76750 249136 76810 249310
rect 78909 249307 78975 249310
rect 87189 249370 87255 249373
rect 87189 249368 90028 249370
rect 87189 249312 87194 249368
rect 87250 249312 90028 249368
rect 87189 249310 90028 249312
rect 87189 249307 87255 249310
rect 142990 249136 143050 249718
rect 181489 249776 184082 249778
rect 181489 249720 181494 249776
rect 181550 249720 184082 249776
rect 181489 249718 184082 249720
rect 181489 249715 181555 249718
rect 184022 249408 184082 249718
rect 232825 249776 237074 249778
rect 232825 249720 232830 249776
rect 232886 249720 237074 249776
rect 232825 249718 237074 249720
rect 232825 249715 232891 249718
rect 225741 249370 225807 249373
rect 223796 249368 225807 249370
rect 223796 249312 225746 249368
rect 225802 249312 225807 249368
rect 223796 249310 225807 249312
rect 225741 249307 225807 249310
rect 237014 249136 237074 249718
rect 278046 249408 278106 249990
rect 360705 249778 360771 249781
rect 358852 249776 360771 249778
rect 358852 249720 360710 249776
rect 360766 249720 360771 249776
rect 358852 249718 360771 249720
rect 360705 249715 360771 249718
rect 321605 249370 321671 249373
rect 317820 249368 321671 249370
rect 317820 249312 321610 249368
rect 321666 249312 321671 249368
rect 317820 249310 321671 249312
rect 321605 249307 321671 249310
rect 173301 249098 173367 249101
rect 266589 249098 266655 249101
rect 170804 249096 173367 249098
rect 170804 249040 173306 249096
rect 173362 249040 173367 249096
rect 170804 249038 173367 249040
rect 264828 249096 266655 249098
rect 264828 249040 266594 249096
rect 266650 249040 266655 249096
rect 264828 249038 266655 249040
rect 173301 249035 173367 249038
rect 266589 249035 266655 249038
rect 328413 249098 328479 249101
rect 328413 249096 331068 249098
rect 328413 249040 328418 249096
rect 328474 249040 331068 249096
rect 328413 249038 331068 249040
rect 328413 249035 328479 249038
rect 132085 248962 132151 248965
rect 129742 248960 132151 248962
rect 129742 248904 132090 248960
rect 132146 248904 132151 248960
rect 129742 248902 132151 248904
rect 129742 248456 129802 248902
rect 132085 248899 132151 248902
rect 274869 248826 274935 248829
rect 274869 248824 278106 248826
rect 274869 248768 274874 248824
rect 274930 248768 278106 248824
rect 274869 248766 278106 248768
rect 274869 248763 274935 248766
rect 181949 248690 182015 248693
rect 181949 248688 184082 248690
rect 181949 248632 181954 248688
rect 182010 248632 184082 248688
rect 181949 248630 184082 248632
rect 181949 248627 182015 248630
rect 184022 248456 184082 248630
rect 278046 248456 278106 248766
rect 87189 248418 87255 248421
rect 139721 248418 139787 248421
rect 225925 248418 225991 248421
rect 87189 248416 90028 248418
rect 87189 248360 87194 248416
rect 87250 248360 90028 248416
rect 87189 248358 90028 248360
rect 139721 248416 143050 248418
rect 139721 248360 139726 248416
rect 139782 248360 143050 248416
rect 139721 248358 143050 248360
rect 223796 248416 225991 248418
rect 223796 248360 225930 248416
rect 225986 248360 225991 248416
rect 223796 248358 225991 248360
rect 87189 248355 87255 248358
rect 139721 248355 139787 248358
rect 132453 248282 132519 248285
rect 129742 248280 132519 248282
rect 129742 248224 132458 248280
rect 132514 248224 132519 248280
rect 129742 248222 132519 248224
rect 78909 248010 78975 248013
rect 76750 248008 78975 248010
rect 76750 247952 78914 248008
rect 78970 247952 78975 248008
rect 76750 247950 78975 247952
rect 76750 247776 76810 247950
rect 78909 247947 78975 247950
rect 129742 247640 129802 248222
rect 132453 248219 132519 248222
rect 142990 247776 143050 248358
rect 225925 248355 225991 248358
rect 233469 248418 233535 248421
rect 321605 248418 321671 248421
rect 233469 248416 237074 248418
rect 233469 248360 233474 248416
rect 233530 248360 237074 248416
rect 233469 248358 237074 248360
rect 317820 248416 321671 248418
rect 317820 248360 321610 248416
rect 321666 248360 321671 248416
rect 317820 248358 321671 248360
rect 233469 248355 233535 248358
rect 181857 248282 181923 248285
rect 181857 248280 184082 248282
rect 181857 248224 181862 248280
rect 181918 248224 184082 248280
rect 181857 248222 184082 248224
rect 181857 248219 181923 248222
rect 173485 247738 173551 247741
rect 170804 247736 173551 247738
rect 170804 247680 173490 247736
rect 173546 247680 173551 247736
rect 170804 247678 173551 247680
rect 173485 247675 173551 247678
rect 184022 247640 184082 248222
rect 237014 247776 237074 248358
rect 321605 248355 321671 248358
rect 274961 248282 275027 248285
rect 274961 248280 278106 248282
rect 274961 248224 274966 248280
rect 275022 248224 278106 248280
rect 274961 248222 278106 248224
rect 274961 248219 275027 248222
rect 266589 247738 266655 247741
rect 264828 247736 266655 247738
rect 264828 247680 266594 247736
rect 266650 247680 266655 247736
rect 264828 247678 266655 247680
rect 266589 247675 266655 247678
rect 278046 247640 278106 248222
rect 328413 247738 328479 247741
rect 328413 247736 331068 247738
rect 328413 247680 328418 247736
rect 328474 247680 331068 247736
rect 328413 247678 331068 247680
rect 328413 247675 328479 247678
rect 88477 247602 88543 247605
rect 226201 247602 226267 247605
rect 321789 247602 321855 247605
rect 88477 247600 90028 247602
rect 88477 247544 88482 247600
rect 88538 247544 90028 247600
rect 88477 247542 90028 247544
rect 223796 247600 226267 247602
rect 223796 247544 226206 247600
rect 226262 247544 226267 247600
rect 223796 247542 226267 247544
rect 317820 247600 321855 247602
rect 317820 247544 321794 247600
rect 321850 247544 321855 247600
rect 317820 247542 321855 247544
rect 88477 247539 88543 247542
rect 226201 247539 226267 247542
rect 321789 247539 321855 247542
rect 274869 247330 274935 247333
rect 274869 247328 278106 247330
rect 274869 247272 274874 247328
rect 274930 247272 278106 247328
rect 274869 247270 278106 247272
rect 274869 247267 274935 247270
rect 182317 247194 182383 247197
rect 182317 247192 184082 247194
rect 182317 247136 182322 247192
rect 182378 247136 184082 247192
rect 182317 247134 184082 247136
rect 182317 247131 182383 247134
rect 132361 247058 132427 247061
rect 129742 247056 132427 247058
rect 129742 247000 132366 247056
rect 132422 247000 132427 247056
rect 129742 246998 132427 247000
rect 78909 246922 78975 246925
rect 76750 246920 78975 246922
rect 76750 246864 78914 246920
rect 78970 246864 78975 246920
rect 76750 246862 78975 246864
rect 49150 246108 49210 246620
rect 76750 246416 76810 246862
rect 78909 246859 78975 246862
rect 129742 246688 129802 246998
rect 132361 246995 132427 246998
rect 140641 246786 140707 246789
rect 140641 246784 143050 246786
rect 140641 246728 140646 246784
rect 140702 246728 143050 246784
rect 140641 246726 143050 246728
rect 140641 246723 140707 246726
rect 87189 246650 87255 246653
rect 87189 246648 90028 246650
rect 87189 246592 87194 246648
rect 87250 246592 90028 246648
rect 87189 246590 90028 246592
rect 87189 246587 87255 246590
rect 142990 246416 143050 246726
rect 184022 246688 184082 247134
rect 234573 246922 234639 246925
rect 234573 246920 237074 246922
rect 234573 246864 234578 246920
rect 234634 246864 237074 246920
rect 234573 246862 237074 246864
rect 234573 246859 234639 246862
rect 226293 246650 226359 246653
rect 223796 246648 226359 246650
rect 223796 246592 226298 246648
rect 226354 246592 226359 246648
rect 223796 246590 226359 246592
rect 226293 246587 226359 246590
rect 237014 246416 237074 246862
rect 278046 246688 278106 247270
rect 328413 246922 328479 246925
rect 328413 246920 331098 246922
rect 328413 246864 328418 246920
rect 328474 246864 331098 246920
rect 328413 246862 331098 246864
rect 328413 246859 328479 246862
rect 321421 246650 321487 246653
rect 317820 246648 321487 246650
rect 317820 246592 321426 246648
rect 321482 246592 321487 246648
rect 317820 246590 321487 246592
rect 321421 246587 321487 246590
rect 331038 246416 331098 246862
rect 360797 246650 360863 246653
rect 358852 246648 360863 246650
rect 358852 246592 360802 246648
rect 360858 246592 360863 246648
rect 358852 246590 360863 246592
rect 360797 246587 360863 246590
rect 173301 246378 173367 246381
rect 267877 246378 267943 246381
rect 170804 246376 173367 246378
rect 170804 246320 173306 246376
rect 173362 246320 173367 246376
rect 170804 246318 173367 246320
rect 264828 246376 267943 246378
rect 264828 246320 267882 246376
rect 267938 246320 267943 246376
rect 264828 246318 267943 246320
rect 173301 246315 173367 246318
rect 267877 246315 267943 246318
rect 49142 246044 49148 246108
rect 49212 246044 49218 246108
rect 132269 246106 132335 246109
rect 129742 246104 132335 246106
rect 129742 246048 132274 246104
rect 132330 246048 132335 246104
rect 129742 246046 132335 246048
rect 129742 245872 129802 246046
rect 132269 246043 132335 246046
rect 274869 246106 274935 246109
rect 274869 246104 278106 246106
rect 274869 246048 274874 246104
rect 274930 246048 278106 246104
rect 274869 246046 278106 246048
rect 274869 246043 274935 246046
rect 278046 245872 278106 246046
rect 87189 245834 87255 245837
rect 182317 245834 182383 245837
rect 226109 245834 226175 245837
rect 321605 245834 321671 245837
rect 87189 245832 90028 245834
rect 87189 245776 87194 245832
rect 87250 245776 90028 245832
rect 87189 245774 90028 245776
rect 182317 245832 184052 245834
rect 182317 245776 182322 245832
rect 182378 245776 184052 245832
rect 182317 245774 184052 245776
rect 223796 245832 226175 245834
rect 223796 245776 226114 245832
rect 226170 245776 226175 245832
rect 223796 245774 226175 245776
rect 317820 245832 321671 245834
rect 317820 245776 321610 245832
rect 321666 245776 321671 245832
rect 317820 245774 321671 245776
rect 87189 245771 87255 245774
rect 182317 245771 182383 245774
rect 226109 245771 226175 245774
rect 321605 245771 321671 245774
rect 78909 245562 78975 245565
rect 131349 245562 131415 245565
rect 76750 245560 78975 245562
rect 76750 245504 78914 245560
rect 78970 245504 78975 245560
rect 76750 245502 78975 245504
rect 76750 244920 76810 245502
rect 78909 245499 78975 245502
rect 129742 245560 131415 245562
rect 129742 245504 131354 245560
rect 131410 245504 131415 245560
rect 129742 245502 131415 245504
rect 129742 244920 129802 245502
rect 131349 245499 131415 245502
rect 138433 245562 138499 245565
rect 138750 245562 138756 245564
rect 138433 245560 138756 245562
rect 138433 245504 138438 245560
rect 138494 245504 138756 245560
rect 138433 245502 138756 245504
rect 138433 245499 138499 245502
rect 138750 245500 138756 245502
rect 138820 245500 138826 245564
rect 140365 245562 140431 245565
rect 233469 245562 233535 245565
rect 274961 245562 275027 245565
rect 327861 245562 327927 245565
rect 140365 245560 143050 245562
rect 140365 245504 140370 245560
rect 140426 245504 143050 245560
rect 140365 245502 143050 245504
rect 140365 245499 140431 245502
rect 142990 244920 143050 245502
rect 233469 245560 237074 245562
rect 233469 245504 233474 245560
rect 233530 245504 237074 245560
rect 233469 245502 237074 245504
rect 233469 245499 233535 245502
rect 181581 245426 181647 245429
rect 181581 245424 184082 245426
rect 181581 245368 181586 245424
rect 181642 245368 184082 245424
rect 181581 245366 184082 245368
rect 181581 245363 181647 245366
rect 184022 244920 184082 245366
rect 237014 244920 237074 245502
rect 274961 245560 278106 245562
rect 274961 245504 274966 245560
rect 275022 245504 278106 245560
rect 274961 245502 278106 245504
rect 274961 245499 275027 245502
rect 278046 244920 278106 245502
rect 327861 245560 331098 245562
rect 327861 245504 327866 245560
rect 327922 245504 331098 245560
rect 327861 245502 331098 245504
rect 327861 245499 327927 245502
rect 331038 244920 331098 245502
rect 87097 244882 87163 244885
rect 172749 244882 172815 244885
rect 225557 244882 225623 244885
rect 266589 244882 266655 244885
rect 321697 244882 321763 244885
rect 87097 244880 90028 244882
rect 87097 244824 87102 244880
rect 87158 244824 90028 244880
rect 87097 244822 90028 244824
rect 170804 244880 172815 244882
rect 170804 244824 172754 244880
rect 172810 244824 172815 244880
rect 170804 244822 172815 244824
rect 223796 244880 225623 244882
rect 223796 244824 225562 244880
rect 225618 244824 225623 244880
rect 223796 244822 225623 244824
rect 264828 244880 266655 244882
rect 264828 244824 266594 244880
rect 266650 244824 266655 244880
rect 264828 244822 266655 244824
rect 317820 244880 321763 244882
rect 317820 244824 321702 244880
rect 321758 244824 321763 244880
rect 317820 244822 321763 244824
rect 87097 244819 87163 244822
rect 172749 244819 172815 244822
rect 225557 244819 225623 244822
rect 266589 244819 266655 244822
rect 321697 244819 321763 244822
rect 132545 244746 132611 244749
rect 129742 244744 132611 244746
rect 129742 244688 132550 244744
rect 132606 244688 132611 244744
rect 129742 244686 132611 244688
rect 78909 244202 78975 244205
rect 76750 244200 78975 244202
rect 76750 244144 78914 244200
rect 78970 244144 78975 244200
rect 76750 244142 78975 244144
rect 76750 243560 76810 244142
rect 78909 244139 78975 244142
rect 129742 244104 129802 244686
rect 132545 244683 132611 244686
rect 182317 244610 182383 244613
rect 274869 244610 274935 244613
rect 182317 244608 184082 244610
rect 182317 244552 182322 244608
rect 182378 244552 184082 244608
rect 182317 244550 184082 244552
rect 182317 244547 182383 244550
rect 184022 244104 184082 244550
rect 274869 244608 278106 244610
rect 274869 244552 274874 244608
rect 274930 244552 278106 244608
rect 274869 244550 278106 244552
rect 274869 244547 274935 244550
rect 234205 244202 234271 244205
rect 234205 244200 237074 244202
rect 234205 244144 234210 244200
rect 234266 244144 237074 244200
rect 234205 244142 237074 244144
rect 234205 244139 234271 244142
rect 87005 244066 87071 244069
rect 140089 244066 140155 244069
rect 225557 244066 225623 244069
rect 87005 244064 90028 244066
rect 87005 244008 87010 244064
rect 87066 244008 90028 244064
rect 87005 244006 90028 244008
rect 140089 244064 143050 244066
rect 140089 244008 140094 244064
rect 140150 244008 143050 244064
rect 140089 244006 143050 244008
rect 223796 244064 225623 244066
rect 223796 244008 225562 244064
rect 225618 244008 225623 244064
rect 223796 244006 225623 244008
rect 87005 244003 87071 244006
rect 140089 244003 140155 244006
rect 142990 243560 143050 244006
rect 225557 244003 225623 244006
rect 237014 243560 237074 244142
rect 278046 244104 278106 244550
rect 321605 244066 321671 244069
rect 317820 244064 321671 244066
rect 317820 244008 321610 244064
rect 321666 244008 321671 244064
rect 317820 244006 321671 244008
rect 321605 244003 321671 244006
rect 327861 244066 327927 244069
rect 327861 244064 331098 244066
rect 327861 244008 327866 244064
rect 327922 244008 331098 244064
rect 327861 244006 331098 244008
rect 327861 244003 327927 244006
rect 331038 243560 331098 244006
rect 46934 243460 46940 243524
rect 47004 243522 47010 243524
rect 173117 243522 173183 243525
rect 266589 243522 266655 243525
rect 360889 243522 360955 243525
rect 47004 243462 48996 243522
rect 170804 243520 173183 243522
rect 170804 243464 173122 243520
rect 173178 243464 173183 243520
rect 170804 243462 173183 243464
rect 264828 243520 266655 243522
rect 264828 243464 266594 243520
rect 266650 243464 266655 243520
rect 264828 243462 266655 243464
rect 358852 243520 360955 243522
rect 358852 243464 360894 243520
rect 360950 243464 360955 243520
rect 358852 243462 360955 243464
rect 47004 243460 47010 243462
rect 173117 243459 173183 243462
rect 266589 243459 266655 243462
rect 360889 243459 360955 243462
rect 181029 243386 181095 243389
rect 275421 243386 275487 243389
rect 181029 243384 184082 243386
rect 181029 243328 181034 243384
rect 181090 243328 184082 243384
rect 181029 243326 184082 243328
rect 181029 243323 181095 243326
rect 184022 243152 184082 243326
rect 275421 243384 278106 243386
rect 275421 243328 275426 243384
rect 275482 243328 278106 243384
rect 275421 243326 278106 243328
rect 275421 243323 275487 243326
rect 278046 243152 278106 243326
rect 87281 243114 87347 243117
rect 132545 243114 132611 243117
rect 226477 243114 226543 243117
rect 321605 243114 321671 243117
rect 87281 243112 90028 243114
rect 87281 243056 87286 243112
rect 87342 243056 90028 243112
rect 87281 243054 90028 243056
rect 129772 243112 132611 243114
rect 129772 243056 132550 243112
rect 132606 243056 132611 243112
rect 129772 243054 132611 243056
rect 223796 243112 226543 243114
rect 223796 243056 226482 243112
rect 226538 243056 226543 243112
rect 223796 243054 226543 243056
rect 317820 243112 321671 243114
rect 317820 243056 321610 243112
rect 321666 243056 321671 243112
rect 317820 243054 321671 243056
rect 87281 243051 87347 243054
rect 132545 243051 132611 243054
rect 226477 243051 226543 243054
rect 321605 243051 321671 243054
rect 9896 242978 10376 243008
rect 13129 242978 13195 242981
rect 9896 242976 13195 242978
rect 9896 242920 13134 242976
rect 13190 242920 13195 242976
rect 9896 242918 13195 242920
rect 9896 242888 10376 242918
rect 13129 242915 13195 242918
rect 132637 242842 132703 242845
rect 129742 242840 132703 242842
rect 129742 242784 132642 242840
rect 132698 242784 132703 242840
rect 129742 242782 132703 242784
rect 78909 242570 78975 242573
rect 76750 242568 78975 242570
rect 76750 242512 78914 242568
rect 78970 242512 78975 242568
rect 76750 242510 78975 242512
rect 76750 242200 76810 242510
rect 78909 242507 78975 242510
rect 129742 242336 129802 242782
rect 132637 242779 132703 242782
rect 138985 242842 139051 242845
rect 181213 242842 181279 242845
rect 233469 242842 233535 242845
rect 275973 242842 276039 242845
rect 138985 242840 143050 242842
rect 138985 242784 138990 242840
rect 139046 242784 143050 242840
rect 138985 242782 143050 242784
rect 138985 242779 139051 242782
rect 87189 242298 87255 242301
rect 87189 242296 90028 242298
rect 87189 242240 87194 242296
rect 87250 242240 90028 242296
rect 87189 242238 90028 242240
rect 87189 242235 87255 242238
rect 142990 242200 143050 242782
rect 181213 242840 184082 242842
rect 181213 242784 181218 242840
rect 181274 242784 184082 242840
rect 181213 242782 184082 242784
rect 181213 242779 181279 242782
rect 184022 242336 184082 242782
rect 233469 242840 237074 242842
rect 233469 242784 233474 242840
rect 233530 242784 237074 242840
rect 233469 242782 237074 242784
rect 233469 242779 233535 242782
rect 225741 242298 225807 242301
rect 223796 242296 225807 242298
rect 223796 242240 225746 242296
rect 225802 242240 225807 242296
rect 223796 242238 225807 242240
rect 225741 242235 225807 242238
rect 237014 242200 237074 242782
rect 275973 242840 278106 242842
rect 275973 242784 275978 242840
rect 276034 242784 278106 242840
rect 275973 242782 278106 242784
rect 275973 242779 276039 242782
rect 278046 242336 278106 242782
rect 327861 242706 327927 242709
rect 327861 242704 331098 242706
rect 327861 242648 327866 242704
rect 327922 242648 331098 242704
rect 327861 242646 331098 242648
rect 327861 242643 327927 242646
rect 320501 242298 320567 242301
rect 317820 242296 320567 242298
rect 317820 242240 320506 242296
rect 320562 242240 320567 242296
rect 317820 242238 320567 242240
rect 320501 242235 320567 242238
rect 331038 242200 331098 242646
rect 174037 242162 174103 242165
rect 267877 242162 267943 242165
rect 170804 242160 174103 242162
rect 170804 242104 174042 242160
rect 174098 242104 174103 242160
rect 170804 242102 174103 242104
rect 264828 242160 267943 242162
rect 264828 242104 267882 242160
rect 267938 242104 267943 242160
rect 264828 242102 267943 242104
rect 174037 242099 174103 242102
rect 267877 242099 267943 242102
rect 96062 241692 96068 241756
rect 96132 241754 96138 241756
rect 98919 241754 98985 241757
rect 104894 241754 104900 241756
rect 96132 241752 104900 241754
rect 96132 241696 98924 241752
rect 98980 241696 104900 241752
rect 96132 241694 104900 241696
rect 96132 241692 96138 241694
rect 98919 241691 98985 241694
rect 104894 241692 104900 241694
rect 104964 241692 104970 241756
rect 84470 241012 84476 241076
rect 84540 241074 84546 241076
rect 93854 241074 93860 241076
rect 84540 241014 93860 241074
rect 84540 241012 84546 241014
rect 93854 241012 93860 241014
rect 93924 241012 93930 241076
rect 138433 240938 138499 240941
rect 138390 240936 138499 240938
rect 138390 240880 138438 240936
rect 138494 240880 138499 240936
rect 138390 240875 138499 240880
rect 138390 240804 138450 240875
rect 138382 240740 138388 240804
rect 138452 240740 138458 240804
rect 78909 240666 78975 240669
rect 76780 240664 78975 240666
rect 76780 240608 78914 240664
rect 78970 240608 78975 240664
rect 76780 240606 78975 240608
rect 78909 240603 78975 240606
rect 140549 240666 140615 240669
rect 173577 240666 173643 240669
rect 140549 240664 143020 240666
rect 140549 240608 140554 240664
rect 140610 240608 143020 240664
rect 140549 240606 143020 240608
rect 170804 240664 173643 240666
rect 170804 240608 173582 240664
rect 173638 240608 173643 240664
rect 170804 240606 173643 240608
rect 140549 240603 140615 240606
rect 173577 240603 173643 240606
rect 222429 240666 222495 240669
rect 222797 240666 222863 240669
rect 222429 240664 222863 240666
rect 222429 240608 222434 240664
rect 222490 240608 222802 240664
rect 222858 240608 222863 240664
rect 222429 240606 222863 240608
rect 222429 240603 222495 240606
rect 222797 240603 222863 240606
rect 233469 240666 233535 240669
rect 267877 240666 267943 240669
rect 233469 240664 237044 240666
rect 233469 240608 233474 240664
rect 233530 240608 237044 240664
rect 233469 240606 237044 240608
rect 264828 240664 267943 240666
rect 264828 240608 267882 240664
rect 267938 240608 267943 240664
rect 264828 240606 267943 240608
rect 233469 240603 233535 240606
rect 267877 240603 267943 240606
rect 327217 240666 327283 240669
rect 327217 240664 331068 240666
rect 327217 240608 327222 240664
rect 327278 240608 331068 240664
rect 327217 240606 331068 240608
rect 327217 240603 327283 240606
rect 49150 239852 49210 240364
rect 196158 240332 196164 240396
rect 196228 240394 196234 240396
rect 196485 240394 196551 240397
rect 305137 240396 305203 240397
rect 196228 240392 196551 240394
rect 196228 240336 196490 240392
rect 196546 240336 196551 240392
rect 196228 240334 196551 240336
rect 196228 240332 196234 240334
rect 196485 240331 196551 240334
rect 305086 240332 305092 240396
rect 305156 240394 305203 240396
rect 360981 240394 361047 240397
rect 305156 240392 305248 240394
rect 305198 240336 305248 240392
rect 305156 240334 305248 240336
rect 358852 240392 361047 240394
rect 358852 240336 360986 240392
rect 361042 240336 361047 240392
rect 358852 240334 361047 240336
rect 305156 240332 305203 240334
rect 305137 240331 305203 240332
rect 360981 240331 361047 240334
rect 429521 240394 429587 240397
rect 434416 240394 434896 240424
rect 429521 240392 434896 240394
rect 429521 240336 429526 240392
rect 429582 240336 434896 240392
rect 429521 240334 434896 240336
rect 429521 240331 429587 240334
rect 434416 240304 434896 240334
rect 49142 239788 49148 239852
rect 49212 239788 49218 239852
rect 294189 239850 294255 239853
rect 295518 239850 295524 239852
rect 294189 239848 295524 239850
rect 294189 239792 294194 239848
rect 294250 239792 295524 239848
rect 294189 239790 295524 239792
rect 294189 239787 294255 239790
rect 295518 239788 295524 239790
rect 295588 239788 295594 239852
rect 95193 239716 95259 239717
rect 95142 239652 95148 239716
rect 95212 239714 95259 239716
rect 95212 239712 95304 239714
rect 95254 239656 95304 239712
rect 95212 239654 95304 239656
rect 95212 239652 95259 239654
rect 187878 239652 187884 239716
rect 187948 239714 187954 239716
rect 189217 239714 189283 239717
rect 187948 239712 189283 239714
rect 187948 239656 189222 239712
rect 189278 239656 189283 239712
rect 187948 239654 189283 239656
rect 187948 239652 187954 239654
rect 95193 239651 95259 239652
rect 189217 239651 189283 239654
rect 324590 239652 324596 239716
rect 324660 239714 324666 239716
rect 325837 239714 325903 239717
rect 324660 239712 325903 239714
rect 324660 239656 325842 239712
rect 325898 239656 325903 239712
rect 324660 239654 325903 239656
rect 324660 239652 324666 239654
rect 325837 239651 325903 239654
rect 91697 239442 91763 239445
rect 92566 239442 92572 239444
rect 91697 239440 92572 239442
rect 91697 239384 91702 239440
rect 91758 239384 92572 239440
rect 91697 239382 92572 239384
rect 91697 239379 91763 239382
rect 92566 239380 92572 239382
rect 92636 239380 92642 239444
rect 192110 239380 192116 239444
rect 192180 239442 192186 239444
rect 192897 239442 192963 239445
rect 283241 239444 283307 239445
rect 283190 239442 283196 239444
rect 192180 239440 192963 239442
rect 192180 239384 192902 239440
rect 192958 239384 192963 239440
rect 192180 239382 192963 239384
rect 283150 239382 283196 239442
rect 283260 239440 283307 239444
rect 283302 239384 283307 239440
rect 192180 239380 192186 239382
rect 192897 239379 192963 239382
rect 283190 239380 283196 239382
rect 283260 239380 283307 239384
rect 283241 239379 283307 239380
rect 79001 239306 79067 239309
rect 76780 239304 79067 239306
rect 76780 239248 79006 239304
rect 79062 239248 79067 239304
rect 76780 239246 79067 239248
rect 79001 239243 79067 239246
rect 140549 239306 140615 239309
rect 173301 239306 173367 239309
rect 140549 239304 143020 239306
rect 140549 239248 140554 239304
rect 140610 239248 143020 239304
rect 140549 239246 143020 239248
rect 170804 239304 173367 239306
rect 170804 239248 173306 239304
rect 173362 239248 173367 239304
rect 170804 239246 173367 239248
rect 140549 239243 140615 239246
rect 173301 239243 173367 239246
rect 233469 239306 233535 239309
rect 266773 239306 266839 239309
rect 233469 239304 237044 239306
rect 233469 239248 233474 239304
rect 233530 239248 237044 239304
rect 233469 239246 237044 239248
rect 264828 239304 266839 239306
rect 264828 239248 266778 239304
rect 266834 239248 266839 239304
rect 264828 239246 266839 239248
rect 233469 239243 233535 239246
rect 266773 239243 266839 239246
rect 328045 239306 328111 239309
rect 328045 239304 331068 239306
rect 328045 239248 328050 239304
rect 328106 239248 331068 239304
rect 328045 239246 331068 239248
rect 328045 239243 328111 239246
rect 79093 238626 79159 238629
rect 76750 238624 79159 238626
rect 76750 238568 79098 238624
rect 79154 238568 79159 238624
rect 76750 238566 79159 238568
rect 76750 237984 76810 238566
rect 79093 238563 79159 238566
rect 138893 238626 138959 238629
rect 234113 238626 234179 238629
rect 327861 238626 327927 238629
rect 138893 238624 143050 238626
rect 138893 238568 138898 238624
rect 138954 238568 143050 238624
rect 138893 238566 143050 238568
rect 138893 238563 138959 238566
rect 142990 237984 143050 238566
rect 234113 238624 237074 238626
rect 234113 238568 234118 238624
rect 234174 238568 237074 238624
rect 234113 238566 237074 238568
rect 234113 238563 234179 238566
rect 198918 238428 198924 238492
rect 198988 238490 198994 238492
rect 200165 238490 200231 238493
rect 198988 238488 200231 238490
rect 198988 238432 200170 238488
rect 200226 238432 200231 238488
rect 198988 238430 200231 238432
rect 198988 238428 198994 238430
rect 200165 238427 200231 238430
rect 237014 237984 237074 238566
rect 327861 238624 331098 238626
rect 327861 238568 327866 238624
rect 327922 238568 331098 238624
rect 327861 238566 331098 238568
rect 327861 238563 327927 238566
rect 290049 238492 290115 238493
rect 289998 238428 290004 238492
rect 290068 238490 290115 238492
rect 290068 238488 290160 238490
rect 290110 238432 290160 238488
rect 290068 238430 290160 238432
rect 290068 238428 290115 238430
rect 290049 238427 290115 238428
rect 331038 237984 331098 238566
rect 100110 237884 100116 237948
rect 100180 237946 100186 237948
rect 102461 237946 102527 237949
rect 173393 237946 173459 237949
rect 100180 237944 102527 237946
rect 100180 237888 102466 237944
rect 102522 237888 102527 237944
rect 100180 237886 102527 237888
rect 170804 237944 173459 237946
rect 170804 237888 173398 237944
rect 173454 237888 173459 237944
rect 170804 237886 173459 237888
rect 100180 237884 100186 237886
rect 102461 237883 102527 237886
rect 173393 237883 173459 237886
rect 230893 237946 230959 237949
rect 231854 237946 231860 237948
rect 230893 237944 231860 237946
rect 230893 237888 230898 237944
rect 230954 237888 231860 237944
rect 230893 237886 231860 237888
rect 230893 237883 230959 237886
rect 231854 237884 231860 237886
rect 231924 237884 231930 237948
rect 267601 237946 267667 237949
rect 264828 237944 267667 237946
rect 264828 237888 267606 237944
rect 267662 237888 267667 237944
rect 264828 237886 267667 237888
rect 267601 237883 267667 237886
rect 219761 237812 219827 237813
rect 219710 237810 219716 237812
rect 219670 237750 219716 237810
rect 219780 237808 219827 237812
rect 219822 237752 219827 237808
rect 219710 237748 219716 237750
rect 219780 237748 219827 237752
rect 219761 237747 219827 237748
rect 141142 237612 141148 237676
rect 141212 237674 141218 237676
rect 143166 237674 143172 237676
rect 141212 237614 143172 237674
rect 141212 237612 141218 237614
rect 143166 237612 143172 237614
rect 143236 237612 143242 237676
rect 47077 237402 47143 237405
rect 361257 237402 361323 237405
rect 47077 237400 48996 237402
rect 47077 237344 47082 237400
rect 47138 237344 48996 237400
rect 47077 237342 48996 237344
rect 358852 237400 361323 237402
rect 358852 237344 361262 237400
rect 361318 237344 361323 237400
rect 358852 237342 361323 237344
rect 47077 237339 47143 237342
rect 361257 237339 361323 237342
rect 140273 237266 140339 237269
rect 140273 237264 143050 237266
rect 140273 237208 140278 237264
rect 140334 237208 143050 237264
rect 140273 237206 143050 237208
rect 140273 237203 140339 237206
rect 89990 236932 89996 236996
rect 90060 236994 90066 236996
rect 100110 236994 100116 236996
rect 90060 236934 100116 236994
rect 90060 236932 90066 236934
rect 100110 236932 100116 236934
rect 100180 236932 100186 236996
rect 142990 236624 143050 237206
rect 233469 237130 233535 237133
rect 233469 237128 237074 237130
rect 233469 237072 233474 237128
rect 233530 237072 237074 237128
rect 233469 237070 237074 237072
rect 233469 237067 233535 237070
rect 186590 236932 186596 236996
rect 186660 236994 186666 236996
rect 198918 236994 198924 236996
rect 186660 236934 198924 236994
rect 186660 236932 186666 236934
rect 198918 236932 198924 236934
rect 198988 236932 198994 236996
rect 237014 236624 237074 237070
rect 264790 236932 264796 236996
rect 264860 236994 264866 236996
rect 273806 236994 273812 236996
rect 264860 236934 273812 236994
rect 264860 236932 264866 236934
rect 273806 236932 273812 236934
rect 273876 236932 273882 236996
rect 78909 236586 78975 236589
rect 172933 236586 172999 236589
rect 267233 236586 267299 236589
rect 76780 236584 78975 236586
rect 76780 236528 78914 236584
rect 78970 236528 78975 236584
rect 76780 236526 78975 236528
rect 170804 236584 172999 236586
rect 170804 236528 172938 236584
rect 172994 236528 172999 236584
rect 170804 236526 172999 236528
rect 264828 236584 267299 236586
rect 264828 236528 267238 236584
rect 267294 236528 267299 236584
rect 264828 236526 267299 236528
rect 78909 236523 78975 236526
rect 172933 236523 172999 236526
rect 267233 236523 267299 236526
rect 328413 236586 328479 236589
rect 369169 236586 369235 236589
rect 328413 236584 331068 236586
rect 328413 236528 328418 236584
rect 328474 236528 331068 236584
rect 328413 236526 331068 236528
rect 369169 236584 371916 236586
rect 369169 236528 369174 236584
rect 369230 236528 371916 236584
rect 369169 236526 371916 236528
rect 328413 236523 328479 236526
rect 369169 236523 369235 236526
rect 74534 236388 74540 236452
rect 74604 236450 74610 236452
rect 75454 236450 75460 236452
rect 74604 236390 75460 236450
rect 74604 236388 74610 236390
rect 75454 236388 75460 236390
rect 75524 236450 75530 236452
rect 81342 236450 81348 236452
rect 75524 236390 81348 236450
rect 75524 236388 75530 236390
rect 81342 236388 81348 236390
rect 81412 236388 81418 236452
rect 203109 236316 203175 236317
rect 286921 236316 286987 236317
rect 73430 236252 73436 236316
rect 73500 236314 73506 236316
rect 74718 236314 74724 236316
rect 73500 236254 74724 236314
rect 73500 236252 73506 236254
rect 74718 236252 74724 236254
rect 74788 236314 74794 236316
rect 76374 236314 76380 236316
rect 74788 236254 76380 236314
rect 74788 236252 74794 236254
rect 76374 236252 76380 236254
rect 76444 236252 76450 236316
rect 203109 236312 203156 236316
rect 203220 236314 203226 236316
rect 203109 236256 203114 236312
rect 203109 236252 203156 236256
rect 203220 236254 203266 236314
rect 203220 236252 203226 236254
rect 286870 236252 286876 236316
rect 286940 236314 286987 236316
rect 286940 236312 287032 236314
rect 286982 236256 287032 236312
rect 286940 236254 287032 236256
rect 286940 236252 286987 236254
rect 203109 236251 203175 236252
rect 286921 236251 286987 236252
rect 244233 236180 244299 236181
rect 73982 236116 73988 236180
rect 74052 236178 74058 236180
rect 76558 236178 76564 236180
rect 74052 236118 76564 236178
rect 74052 236116 74058 236118
rect 76558 236116 76564 236118
rect 76628 236116 76634 236180
rect 167822 236116 167828 236180
rect 167892 236178 167898 236180
rect 177022 236178 177028 236180
rect 167892 236118 177028 236178
rect 167892 236116 167898 236118
rect 177022 236116 177028 236118
rect 177092 236116 177098 236180
rect 244182 236116 244188 236180
rect 244252 236178 244299 236180
rect 369445 236178 369511 236181
rect 244252 236176 244344 236178
rect 244294 236120 244344 236176
rect 244252 236118 244344 236120
rect 369445 236176 371916 236178
rect 369445 236120 369450 236176
rect 369506 236120 371916 236176
rect 369445 236118 371916 236120
rect 244252 236116 244299 236118
rect 244233 236115 244299 236116
rect 369445 236115 369511 236118
rect 73614 235980 73620 236044
rect 73684 236042 73690 236044
rect 76006 236042 76012 236044
rect 73684 235982 76012 236042
rect 73684 235980 73690 235982
rect 76006 235980 76012 235982
rect 76076 235980 76082 236044
rect 147766 235980 147772 236044
rect 147836 236042 147842 236044
rect 148737 236042 148803 236045
rect 147836 236040 148803 236042
rect 147836 235984 148742 236040
rect 148798 235984 148803 236040
rect 147836 235982 148803 235984
rect 147836 235980 147842 235982
rect 148737 235979 148803 235982
rect 167965 236042 168031 236045
rect 168190 236042 168196 236044
rect 167965 236040 168196 236042
rect 167965 235984 167970 236040
rect 168026 235984 168196 236040
rect 167965 235982 168196 235984
rect 167965 235979 168031 235982
rect 168190 235980 168196 235982
rect 168260 235980 168266 236044
rect 75638 235844 75644 235908
rect 75708 235906 75714 235908
rect 76926 235906 76932 235908
rect 75708 235846 76932 235906
rect 75708 235844 75714 235846
rect 76926 235844 76932 235846
rect 76996 235844 77002 235908
rect 116118 235844 116124 235908
rect 116188 235906 116194 235908
rect 117089 235906 117155 235909
rect 136869 235906 136935 235909
rect 116188 235904 136935 235906
rect 116188 235848 117094 235904
rect 117150 235848 136874 235904
rect 136930 235848 136935 235904
rect 116188 235846 136935 235848
rect 116188 235844 116194 235846
rect 117089 235843 117155 235846
rect 136869 235843 136935 235846
rect 147265 235906 147331 235909
rect 148686 235906 148692 235908
rect 147265 235904 148692 235906
rect 147265 235848 147270 235904
rect 147326 235848 148692 235904
rect 147265 235846 148692 235848
rect 147265 235843 147331 235846
rect 148686 235844 148692 235846
rect 148756 235844 148762 235908
rect 242485 235906 242551 235909
rect 247126 235906 247132 235908
rect 242485 235904 247132 235906
rect 242485 235848 242490 235904
rect 242546 235848 247132 235904
rect 242485 235846 247132 235848
rect 242485 235843 242551 235846
rect 247126 235844 247132 235846
rect 247196 235844 247202 235908
rect 105078 235708 105084 235772
rect 105148 235770 105154 235772
rect 106141 235770 106207 235773
rect 137053 235770 137119 235773
rect 105148 235768 137119 235770
rect 105148 235712 106146 235768
rect 106202 235712 137058 235768
rect 137114 235712 137119 235768
rect 105148 235710 137119 235712
rect 105148 235708 105154 235710
rect 106141 235707 106207 235710
rect 137053 235707 137119 235710
rect 167689 235770 167755 235773
rect 262541 235772 262607 235773
rect 167822 235770 167828 235772
rect 167689 235768 167828 235770
rect 167689 235712 167694 235768
rect 167750 235712 167828 235768
rect 167689 235710 167828 235712
rect 167689 235707 167755 235710
rect 167822 235708 167828 235710
rect 167892 235708 167898 235772
rect 262541 235768 262588 235772
rect 262652 235770 262658 235772
rect 369629 235770 369695 235773
rect 262541 235712 262546 235768
rect 262541 235708 262588 235712
rect 262652 235710 262698 235770
rect 369629 235768 371916 235770
rect 369629 235712 369634 235768
rect 369690 235712 371916 235768
rect 369629 235710 371916 235712
rect 262652 235708 262658 235710
rect 262541 235707 262607 235708
rect 369629 235707 369695 235710
rect 152003 235636 152069 235637
rect 74350 235572 74356 235636
rect 74420 235634 74426 235636
rect 74902 235634 74908 235636
rect 74420 235574 74908 235634
rect 74420 235572 74426 235574
rect 74902 235572 74908 235574
rect 74972 235572 74978 235636
rect 124398 235572 124404 235636
rect 124468 235634 124474 235636
rect 133966 235634 133972 235636
rect 124468 235574 133972 235634
rect 124468 235572 124474 235574
rect 133966 235572 133972 235574
rect 134036 235572 134042 235636
rect 151998 235572 152004 235636
rect 152068 235634 152074 235636
rect 158806 235634 158812 235636
rect 152068 235574 158812 235634
rect 152068 235572 152074 235574
rect 158806 235572 158812 235574
rect 158876 235572 158882 235636
rect 246027 235634 246093 235637
rect 246206 235634 246212 235636
rect 246027 235632 246212 235634
rect 246027 235576 246032 235632
rect 246088 235576 246212 235632
rect 246027 235574 246212 235576
rect 152003 235571 152069 235572
rect 246027 235571 246093 235574
rect 246206 235572 246212 235574
rect 246276 235572 246282 235636
rect 74534 235436 74540 235500
rect 74604 235498 74610 235500
rect 75454 235498 75460 235500
rect 74604 235438 75460 235498
rect 74604 235436 74610 235438
rect 75454 235436 75460 235438
rect 75524 235436 75530 235500
rect 145149 235364 145215 235365
rect 145149 235360 145196 235364
rect 145260 235362 145266 235364
rect 369813 235362 369879 235365
rect 145149 235304 145154 235360
rect 145149 235300 145196 235304
rect 145260 235302 145306 235362
rect 369813 235360 371916 235362
rect 369813 235304 369818 235360
rect 369874 235304 371916 235360
rect 369813 235302 371916 235304
rect 145260 235300 145266 235302
rect 145149 235299 145215 235300
rect 369813 235299 369879 235302
rect 74677 235090 74743 235093
rect 75270 235090 75276 235092
rect 74677 235088 75276 235090
rect 74677 235032 74682 235088
rect 74738 235032 75276 235088
rect 74677 235030 75276 235032
rect 74677 235027 74743 235030
rect 75270 235028 75276 235030
rect 75340 235090 75346 235092
rect 76057 235090 76123 235093
rect 75340 235088 76123 235090
rect 75340 235032 76062 235088
rect 76118 235032 76123 235088
rect 75340 235030 76123 235032
rect 75340 235028 75346 235030
rect 76057 235027 76123 235030
rect 136358 235028 136364 235092
rect 136428 235090 136434 235092
rect 136869 235090 136935 235093
rect 136428 235088 136935 235090
rect 136428 235032 136874 235088
rect 136930 235032 136935 235088
rect 136428 235030 136935 235032
rect 136428 235028 136434 235030
rect 136869 235027 136935 235030
rect 136961 234954 137027 234957
rect 148185 234956 148251 234957
rect 137278 234954 137284 234956
rect 136961 234952 137284 234954
rect 136961 234896 136966 234952
rect 137022 234896 137284 234952
rect 136961 234894 137284 234896
rect 136961 234891 137027 234894
rect 137278 234892 137284 234894
rect 137348 234892 137354 234956
rect 148134 234892 148140 234956
rect 148204 234954 148251 234956
rect 231169 234954 231235 234957
rect 231302 234954 231308 234956
rect 148204 234952 148296 234954
rect 148246 234896 148296 234952
rect 148204 234894 148296 234896
rect 231169 234952 231308 234954
rect 231169 234896 231174 234952
rect 231230 234896 231308 234952
rect 231169 234894 231308 234896
rect 148204 234892 148251 234894
rect 148185 234891 148251 234892
rect 231169 234891 231235 234894
rect 231302 234892 231308 234894
rect 231372 234892 231378 234956
rect 245470 234892 245476 234956
rect 245540 234954 245546 234956
rect 246625 234954 246691 234957
rect 301089 234956 301155 234957
rect 245540 234952 246691 234954
rect 245540 234896 246630 234952
rect 246686 234896 246691 234952
rect 245540 234894 246691 234896
rect 245540 234892 245546 234894
rect 246625 234891 246691 234894
rect 301038 234892 301044 234956
rect 301108 234954 301155 234956
rect 369997 234954 370063 234957
rect 301108 234952 301200 234954
rect 301150 234896 301200 234952
rect 301108 234894 301200 234896
rect 369997 234952 371916 234954
rect 369997 234896 370002 234952
rect 370058 234896 371916 234952
rect 369997 234894 371916 234896
rect 301108 234892 301155 234894
rect 301089 234891 301155 234892
rect 369997 234891 370063 234894
rect 210009 234546 210075 234549
rect 231169 234546 231235 234549
rect 210009 234544 231235 234546
rect 210009 234488 210014 234544
rect 210070 234488 231174 234544
rect 231230 234488 231235 234544
rect 210009 234486 231235 234488
rect 210009 234483 210075 234486
rect 231169 234483 231235 234486
rect 369905 234546 369971 234549
rect 369905 234544 371916 234546
rect 369905 234488 369910 234544
rect 369966 234488 371916 234544
rect 369905 234486 371916 234488
rect 369905 234483 369971 234486
rect 207249 234412 207315 234413
rect 207198 234410 207204 234412
rect 207122 234350 207204 234410
rect 207268 234410 207315 234412
rect 230709 234410 230775 234413
rect 207268 234408 230775 234410
rect 207310 234352 230714 234408
rect 230770 234352 230775 234408
rect 207198 234348 207204 234350
rect 207268 234350 230775 234352
rect 207268 234348 207315 234350
rect 207249 234347 207315 234348
rect 230709 234347 230775 234350
rect 283190 234348 283196 234412
rect 283260 234410 283266 234412
rect 324641 234410 324707 234413
rect 283260 234408 324707 234410
rect 283260 234352 324646 234408
rect 324702 234352 324707 234408
rect 283260 234350 324707 234352
rect 283260 234348 283266 234350
rect 324641 234347 324707 234350
rect 137329 234274 137395 234277
rect 137646 234274 137652 234276
rect 137329 234272 137652 234274
rect 137329 234216 137334 234272
rect 137390 234216 137652 234272
rect 137329 234214 137652 234216
rect 137329 234211 137395 234214
rect 137646 234212 137652 234214
rect 137716 234212 137722 234276
rect 230709 234140 230775 234141
rect 73798 234076 73804 234140
rect 73868 234138 73874 234140
rect 75638 234138 75644 234140
rect 73868 234078 75644 234138
rect 73868 234076 73874 234078
rect 75638 234076 75644 234078
rect 75708 234076 75714 234140
rect 230709 234138 230756 234140
rect 230664 234136 230756 234138
rect 230664 234080 230714 234136
rect 230664 234078 230756 234080
rect 230709 234076 230756 234078
rect 230820 234076 230826 234140
rect 368709 234138 368775 234141
rect 368709 234136 371916 234138
rect 368709 234080 368714 234136
rect 368770 234080 371916 234136
rect 368709 234078 371916 234080
rect 230709 234075 230775 234076
rect 368709 234075 368775 234078
rect 74166 233804 74172 233868
rect 74236 233866 74242 233868
rect 74902 233866 74908 233868
rect 74236 233806 74908 233866
rect 74236 233804 74242 233806
rect 74902 233804 74908 233806
rect 74972 233804 74978 233868
rect 74125 233730 74191 233733
rect 74902 233730 74908 233732
rect 74125 233728 74908 233730
rect 74125 233672 74130 233728
rect 74186 233672 74908 233728
rect 74125 233670 74908 233672
rect 74125 233667 74191 233670
rect 74902 233668 74908 233670
rect 74972 233668 74978 233732
rect 150669 233730 150735 233733
rect 156782 233730 156788 233732
rect 150669 233728 156788 233730
rect 150669 233672 150674 233728
rect 150730 233672 156788 233728
rect 150669 233670 156788 233672
rect 150669 233667 150735 233670
rect 156782 233668 156788 233670
rect 156852 233668 156858 233732
rect 243037 233730 243103 233733
rect 261662 233730 261668 233732
rect 243037 233728 261668 233730
rect 243037 233672 243042 233728
rect 243098 233672 261668 233728
rect 243037 233670 261668 233672
rect 243037 233667 243103 233670
rect 261662 233668 261668 233670
rect 261732 233668 261738 233732
rect 368709 233730 368775 233733
rect 368709 233728 371916 233730
rect 368709 233672 368714 233728
rect 368770 233672 371916 233728
rect 368709 233670 371916 233672
rect 368709 233667 368775 233670
rect 241473 233458 241539 233461
rect 249886 233458 249892 233460
rect 241473 233456 249892 233458
rect 241473 233400 241478 233456
rect 241534 233400 249892 233456
rect 241473 233398 249892 233400
rect 241473 233395 241539 233398
rect 249886 233396 249892 233398
rect 249956 233396 249962 233460
rect 368801 233458 368867 233461
rect 368801 233456 371916 233458
rect 368801 233400 368806 233456
rect 368862 233400 371916 233456
rect 368801 233398 371916 233400
rect 368801 233395 368867 233398
rect 246625 233322 246691 233325
rect 262030 233322 262036 233324
rect 246625 233320 262036 233322
rect 246625 233264 246630 233320
rect 246686 233264 262036 233320
rect 246625 233262 262036 233264
rect 246625 233259 246691 233262
rect 262030 233260 262036 233262
rect 262100 233260 262106 233324
rect 368709 233050 368775 233053
rect 368709 233048 371916 233050
rect 368709 232992 368714 233048
rect 368770 232992 371916 233048
rect 368709 232990 371916 232992
rect 368709 232987 368775 232990
rect 369721 232642 369787 232645
rect 369721 232640 371916 232642
rect 369721 232584 369726 232640
rect 369782 232584 371916 232640
rect 369721 232582 371916 232584
rect 369721 232579 369787 232582
rect 52638 232444 52644 232508
rect 52708 232506 52714 232508
rect 53517 232506 53583 232509
rect 52708 232504 53583 232506
rect 52708 232448 53522 232504
rect 53578 232448 53583 232504
rect 52708 232446 53583 232448
rect 52708 232444 52714 232446
rect 53517 232443 53583 232446
rect 54529 232506 54595 232509
rect 55541 232508 55607 232509
rect 54662 232506 54668 232508
rect 54529 232504 54668 232506
rect 54529 232448 54534 232504
rect 54590 232448 54668 232504
rect 54529 232446 54668 232448
rect 54529 232443 54595 232446
rect 54662 232444 54668 232446
rect 54732 232444 54738 232508
rect 55541 232504 55588 232508
rect 55652 232506 55658 232508
rect 55541 232448 55546 232504
rect 55541 232444 55588 232448
rect 55652 232446 55698 232506
rect 55652 232444 55658 232446
rect 239582 232444 239588 232508
rect 239652 232506 239658 232508
rect 239909 232506 239975 232509
rect 239652 232504 239975 232506
rect 239652 232448 239914 232504
rect 239970 232448 239975 232504
rect 239652 232446 239975 232448
rect 239652 232444 239658 232446
rect 55541 232443 55607 232444
rect 239909 232443 239975 232446
rect 350953 232506 351019 232509
rect 351638 232506 351644 232508
rect 350953 232504 351644 232506
rect 350953 232448 350958 232504
rect 351014 232448 351644 232504
rect 350953 232446 351644 232448
rect 350953 232443 351019 232446
rect 351638 232444 351644 232446
rect 351708 232444 351714 232508
rect 351822 232444 351828 232508
rect 351892 232506 351898 232508
rect 352057 232506 352123 232509
rect 351892 232504 352123 232506
rect 351892 232448 352062 232504
rect 352118 232448 352123 232504
rect 351892 232446 352123 232448
rect 351892 232444 351898 232446
rect 352057 232443 352123 232446
rect 368709 232234 368775 232237
rect 368709 232232 371916 232234
rect 368709 232176 368714 232232
rect 368770 232176 371916 232232
rect 368709 232174 371916 232176
rect 368709 232171 368775 232174
rect 368801 231826 368867 231829
rect 368801 231824 371916 231826
rect 368801 231768 368806 231824
rect 368862 231768 371916 231824
rect 368801 231766 371916 231768
rect 368801 231763 368867 231766
rect 368893 231418 368959 231421
rect 368893 231416 371916 231418
rect 368893 231360 368898 231416
rect 368954 231360 371916 231416
rect 368893 231358 371916 231360
rect 368893 231355 368959 231358
rect 368801 231010 368867 231013
rect 368801 231008 371916 231010
rect 368801 230952 368806 231008
rect 368862 230952 371916 231008
rect 368801 230950 371916 230952
rect 368801 230947 368867 230950
rect 368709 230602 368775 230605
rect 368709 230600 371916 230602
rect 368709 230544 368714 230600
rect 368770 230544 371916 230600
rect 368709 230542 371916 230544
rect 368709 230539 368775 230542
rect 368893 230194 368959 230197
rect 368893 230192 371916 230194
rect 368893 230136 368898 230192
rect 368954 230136 371916 230192
rect 368893 230134 371916 230136
rect 368893 230131 368959 230134
rect 369537 229922 369603 229925
rect 369537 229920 371916 229922
rect 369537 229864 369542 229920
rect 369598 229864 371916 229920
rect 369537 229862 371916 229864
rect 369537 229859 369603 229862
rect 9896 229650 10376 229680
rect 13037 229650 13103 229653
rect 9896 229648 13103 229650
rect 9896 229592 13042 229648
rect 13098 229592 13103 229648
rect 9896 229590 13103 229592
rect 9896 229560 10376 229590
rect 13037 229587 13103 229590
rect 368709 229514 368775 229517
rect 368709 229512 371916 229514
rect 368709 229456 368714 229512
rect 368770 229456 371916 229512
rect 368709 229454 371916 229456
rect 368709 229451 368775 229454
rect 368801 229106 368867 229109
rect 368801 229104 371916 229106
rect 368801 229048 368806 229104
rect 368862 229048 371916 229104
rect 368801 229046 371916 229048
rect 368801 229043 368867 229046
rect 368709 228698 368775 228701
rect 368709 228696 371916 228698
rect 368709 228640 368714 228696
rect 368770 228640 371916 228696
rect 368709 228638 371916 228640
rect 368709 228635 368775 228638
rect 368709 228290 368775 228293
rect 368709 228288 371916 228290
rect 368709 228232 368714 228288
rect 368770 228232 371916 228288
rect 368709 228230 371916 228232
rect 368709 228227 368775 228230
rect 369537 227882 369603 227885
rect 428693 227882 428759 227885
rect 434416 227882 434896 227912
rect 369537 227880 371916 227882
rect 369537 227824 369542 227880
rect 369598 227824 371916 227880
rect 369537 227822 371916 227824
rect 428693 227880 434896 227882
rect 428693 227824 428698 227880
rect 428754 227824 434896 227880
rect 428693 227822 434896 227824
rect 369537 227819 369603 227822
rect 428693 227819 428759 227822
rect 434416 227792 434896 227822
rect 368801 227474 368867 227477
rect 368801 227472 371916 227474
rect 368801 227416 368806 227472
rect 368862 227416 371916 227472
rect 368801 227414 371916 227416
rect 368801 227411 368867 227414
rect 185854 227004 185860 227068
rect 185924 227066 185930 227068
rect 193030 227066 193036 227068
rect 185924 227006 193036 227066
rect 185924 227004 185930 227006
rect 193030 227004 193036 227006
rect 193100 227004 193106 227068
rect 368709 227066 368775 227069
rect 368709 227064 371916 227066
rect 368709 227008 368714 227064
rect 368770 227008 371916 227064
rect 368709 227006 371916 227008
rect 368709 227003 368775 227006
rect 55398 226868 55404 226932
rect 55468 226930 55474 226932
rect 55541 226930 55607 226933
rect 55468 226928 55607 226930
rect 55468 226872 55546 226928
rect 55602 226872 55607 226928
rect 55468 226870 55607 226872
rect 55468 226868 55474 226870
rect 55541 226867 55607 226870
rect 174078 226868 174084 226932
rect 174148 226930 174154 226932
rect 174148 226870 183714 226930
rect 174148 226868 174154 226870
rect 116118 226732 116124 226796
rect 116188 226794 116194 226796
rect 135438 226794 135444 226796
rect 116188 226734 135444 226794
rect 116188 226732 116194 226734
rect 135438 226732 135444 226734
rect 135508 226732 135514 226796
rect 154758 226596 154764 226660
rect 154828 226658 154834 226660
rect 164377 226658 164443 226661
rect 154828 226656 164443 226658
rect 154828 226600 164382 226656
rect 164438 226600 164443 226656
rect 154828 226598 164443 226600
rect 183654 226658 183714 226870
rect 185854 226658 185860 226660
rect 183654 226598 185860 226658
rect 154828 226596 154834 226598
rect 164377 226595 164443 226598
rect 185854 226596 185860 226598
rect 185924 226596 185930 226660
rect 369721 226658 369787 226661
rect 369721 226656 371916 226658
rect 369721 226600 369726 226656
rect 369782 226600 371916 226656
rect 369721 226598 371916 226600
rect 369721 226595 369787 226598
rect 92566 226460 92572 226524
rect 92636 226522 92642 226524
rect 109126 226522 109132 226524
rect 92636 226462 109132 226522
rect 92636 226460 92642 226462
rect 109126 226460 109132 226462
rect 109196 226460 109202 226524
rect 109494 226460 109500 226524
rect 109564 226522 109570 226524
rect 116118 226522 116124 226524
rect 109564 226462 116124 226522
rect 109564 226460 109570 226462
rect 116118 226460 116124 226462
rect 116188 226460 116194 226524
rect 135438 226460 135444 226524
rect 135508 226522 135514 226524
rect 174078 226522 174084 226524
rect 135508 226462 137714 226522
rect 135508 226460 135514 226462
rect 137237 226386 137303 226389
rect 134740 226384 137303 226386
rect 134740 226328 137242 226384
rect 137298 226328 137303 226384
rect 134740 226326 137303 226328
rect 137654 226386 137714 226462
rect 167278 226462 174084 226522
rect 154758 226386 154764 226388
rect 137654 226326 154764 226386
rect 137237 226323 137303 226326
rect 154758 226324 154764 226326
rect 154828 226324 154834 226388
rect 164377 226250 164443 226253
rect 167278 226250 167338 226462
rect 174078 226460 174084 226462
rect 174148 226460 174154 226524
rect 178678 226460 178684 226524
rect 178748 226522 178754 226524
rect 182910 226522 182916 226524
rect 178748 226462 182916 226522
rect 178748 226460 178754 226462
rect 182910 226460 182916 226462
rect 182980 226460 182986 226524
rect 193214 226460 193220 226524
rect 193284 226522 193290 226524
rect 369077 226522 369143 226525
rect 193284 226520 369143 226522
rect 193284 226464 369082 226520
rect 369138 226464 369143 226520
rect 193284 226462 369143 226464
rect 193284 226460 193290 226462
rect 369077 226459 369143 226462
rect 231169 226386 231235 226389
rect 322985 226386 323051 226389
rect 324733 226386 324799 226389
rect 228764 226384 231235 226386
rect 228764 226328 231174 226384
rect 231230 226328 231235 226384
rect 228764 226326 231235 226328
rect 322788 226384 324799 226386
rect 322788 226328 322990 226384
rect 323046 226328 324738 226384
rect 324794 226328 324799 226384
rect 322788 226326 324799 226328
rect 231169 226323 231235 226326
rect 322985 226323 323051 226326
rect 324733 226323 324799 226326
rect 368893 226386 368959 226389
rect 368893 226384 371916 226386
rect 368893 226328 368898 226384
rect 368954 226328 371916 226384
rect 368893 226326 371916 226328
rect 368893 226323 368959 226326
rect 164377 226248 167338 226250
rect 164377 226192 164382 226248
rect 164438 226192 167338 226248
rect 164377 226190 167338 226192
rect 164377 226187 164443 226190
rect 368801 225978 368867 225981
rect 368801 225976 371916 225978
rect 368801 225920 368806 225976
rect 368862 225920 371916 225976
rect 368801 225918 371916 225920
rect 368801 225915 368867 225918
rect 368709 225570 368775 225573
rect 368709 225568 371916 225570
rect 368709 225512 368714 225568
rect 368770 225512 371916 225568
rect 368709 225510 371916 225512
rect 368709 225507 368775 225510
rect 368801 225162 368867 225165
rect 368801 225160 371916 225162
rect 368801 225104 368806 225160
rect 368862 225104 371916 225160
rect 368801 225102 371916 225104
rect 368801 225099 368867 225102
rect 368709 224754 368775 224757
rect 368709 224752 371916 224754
rect 368709 224696 368714 224752
rect 368770 224696 371916 224752
rect 368709 224694 371916 224696
rect 368709 224691 368775 224694
rect 73798 224284 73804 224348
rect 73868 224346 73874 224348
rect 73941 224346 74007 224349
rect 73868 224344 74007 224346
rect 73868 224288 73946 224344
rect 74002 224288 74007 224344
rect 73868 224286 74007 224288
rect 73868 224284 73874 224286
rect 73941 224283 74007 224286
rect 368893 224346 368959 224349
rect 368893 224344 371916 224346
rect 368893 224288 368898 224344
rect 368954 224288 371916 224344
rect 368893 224286 371916 224288
rect 368893 224283 368959 224286
rect 73798 224148 73804 224212
rect 73868 224210 73874 224212
rect 74534 224210 74540 224212
rect 73868 224150 74540 224210
rect 73868 224148 73874 224150
rect 74534 224148 74540 224150
rect 74604 224148 74610 224212
rect 73798 224012 73804 224076
rect 73868 224074 73874 224076
rect 74534 224074 74540 224076
rect 73868 224014 74540 224074
rect 73868 224012 73874 224014
rect 74534 224012 74540 224014
rect 74604 224012 74610 224076
rect 73798 223876 73804 223940
rect 73868 223938 73874 223940
rect 73941 223938 74007 223941
rect 73868 223936 74007 223938
rect 73868 223880 73946 223936
rect 74002 223880 74007 223936
rect 73868 223878 74007 223880
rect 73868 223876 73874 223878
rect 73941 223875 74007 223878
rect 368801 223938 368867 223941
rect 368801 223936 371916 223938
rect 368801 223880 368806 223936
rect 368862 223880 371916 223936
rect 368801 223878 371916 223880
rect 368801 223875 368867 223878
rect 369813 223530 369879 223533
rect 369813 223528 371916 223530
rect 369813 223472 369818 223528
rect 369874 223472 371916 223528
rect 369813 223470 371916 223472
rect 369813 223467 369879 223470
rect 137329 223258 137395 223261
rect 230709 223258 230775 223261
rect 324641 223258 324707 223261
rect 134740 223256 137395 223258
rect 134740 223200 137334 223256
rect 137390 223200 137395 223256
rect 134740 223198 137395 223200
rect 228764 223256 230775 223258
rect 228764 223200 230714 223256
rect 230770 223200 230775 223256
rect 228764 223198 230775 223200
rect 322788 223256 324707 223258
rect 322788 223200 324646 223256
rect 324702 223200 324707 223256
rect 322788 223198 324707 223200
rect 137329 223195 137395 223198
rect 230709 223195 230775 223198
rect 324641 223195 324707 223198
rect 368709 223258 368775 223261
rect 368709 223256 371916 223258
rect 368709 223200 368714 223256
rect 368770 223200 371916 223256
rect 368709 223198 371916 223200
rect 368709 223195 368775 223198
rect 369077 222850 369143 222853
rect 369077 222848 371916 222850
rect 369077 222792 369082 222848
rect 369138 222792 371916 222848
rect 369077 222790 371916 222792
rect 369077 222787 369143 222790
rect 368801 222442 368867 222445
rect 368801 222440 371916 222442
rect 368801 222384 368806 222440
rect 368862 222384 371916 222440
rect 368801 222382 371916 222384
rect 368801 222379 368867 222382
rect 50573 222034 50639 222037
rect 55398 222034 55404 222036
rect 50573 222032 55404 222034
rect 50573 221976 50578 222032
rect 50634 221976 55404 222032
rect 50573 221974 55404 221976
rect 50573 221971 50639 221974
rect 55398 221972 55404 221974
rect 55468 221972 55474 222036
rect 369077 222034 369143 222037
rect 369077 222032 371916 222034
rect 369077 221976 369082 222032
rect 369138 221976 371916 222032
rect 369077 221974 371916 221976
rect 369077 221971 369143 221974
rect 38521 221762 38587 221765
rect 35718 221760 38587 221762
rect 35718 221704 38526 221760
rect 38582 221704 38587 221760
rect 35718 221702 38587 221704
rect 35718 221528 35778 221702
rect 38521 221699 38587 221702
rect 368709 221626 368775 221629
rect 406613 221626 406679 221629
rect 368709 221624 371916 221626
rect 368709 221568 368714 221624
rect 368770 221568 371916 221624
rect 368709 221566 371916 221568
rect 406613 221624 408930 221626
rect 406613 221568 406618 221624
rect 406674 221568 408930 221624
rect 406613 221566 408930 221568
rect 368709 221563 368775 221566
rect 406613 221563 406679 221566
rect 408870 221460 408930 221566
rect 53241 221354 53307 221357
rect 55582 221354 55588 221356
rect 53241 221352 55588 221354
rect 53241 221296 53246 221352
rect 53302 221296 55588 221352
rect 53241 221294 55588 221296
rect 53241 221291 53307 221294
rect 55582 221292 55588 221294
rect 55652 221354 55658 221356
rect 56318 221354 56324 221356
rect 55652 221294 56324 221354
rect 55652 221292 55658 221294
rect 56318 221292 56324 221294
rect 56388 221292 56394 221356
rect 368985 221218 369051 221221
rect 368985 221216 371916 221218
rect 368985 221160 368990 221216
rect 369046 221160 371916 221216
rect 368985 221158 371916 221160
rect 368985 221155 369051 221158
rect 70678 220402 70738 220916
rect 368801 220810 368867 220813
rect 368801 220808 371916 220810
rect 368801 220752 368806 220808
rect 368862 220752 371916 220808
rect 368801 220750 371916 220752
rect 368801 220747 368867 220750
rect 74217 220402 74283 220405
rect 70678 220400 74283 220402
rect 70678 220344 74222 220400
rect 74278 220344 74283 220400
rect 70678 220342 74283 220344
rect 74217 220339 74283 220342
rect 368709 220402 368775 220405
rect 368709 220400 371916 220402
rect 368709 220344 368714 220400
rect 368770 220344 371916 220400
rect 368709 220342 371916 220344
rect 368709 220339 368775 220342
rect 52045 220266 52111 220269
rect 355093 220266 355159 220269
rect 427405 220266 427471 220269
rect 52045 220264 55068 220266
rect 16165 219994 16231 219997
rect 20078 219994 20138 220236
rect 52045 220208 52050 220264
rect 52106 220208 55068 220264
rect 52045 220206 55068 220208
rect 352780 220264 355159 220266
rect 352780 220208 355098 220264
rect 355154 220208 355159 220264
rect 352780 220206 355159 220208
rect 424724 220264 427471 220266
rect 424724 220208 427410 220264
rect 427466 220208 427471 220264
rect 424724 220206 427471 220208
rect 52045 220203 52111 220206
rect 355093 220203 355159 220206
rect 427405 220203 427471 220206
rect 137145 220130 137211 220133
rect 230985 220130 231051 220133
rect 325745 220130 325811 220133
rect 134740 220128 137211 220130
rect 134740 220072 137150 220128
rect 137206 220072 137211 220128
rect 134740 220070 137211 220072
rect 228764 220128 231051 220130
rect 228764 220072 230990 220128
rect 231046 220072 231051 220128
rect 228764 220070 231051 220072
rect 322788 220128 325811 220130
rect 322788 220072 325750 220128
rect 325806 220072 325811 220128
rect 322788 220070 325811 220072
rect 137145 220067 137211 220070
rect 230985 220067 231051 220070
rect 325745 220067 325811 220070
rect 16165 219992 20138 219994
rect 16165 219936 16170 219992
rect 16226 219936 20138 219992
rect 16165 219934 20138 219936
rect 358037 219994 358103 219997
rect 358221 219994 358287 219997
rect 358037 219992 358287 219994
rect 358037 219936 358042 219992
rect 358098 219936 358226 219992
rect 358282 219936 358287 219992
rect 358037 219934 358287 219936
rect 16165 219931 16231 219934
rect 358037 219931 358103 219934
rect 358221 219931 358287 219934
rect 369261 219994 369327 219997
rect 369261 219992 371916 219994
rect 369261 219936 369266 219992
rect 369322 219936 371916 219992
rect 369261 219934 371916 219936
rect 369261 219931 369327 219934
rect 368709 219722 368775 219725
rect 368709 219720 371916 219722
rect 368709 219664 368714 219720
rect 368770 219664 371916 219720
rect 368709 219662 371916 219664
rect 368709 219659 368775 219662
rect 81669 219586 81735 219589
rect 178913 219586 178979 219589
rect 272937 219586 273003 219589
rect 81669 219584 85060 219586
rect 81669 219528 81674 219584
rect 81730 219528 85060 219584
rect 81669 219526 85060 219528
rect 178900 219584 178979 219586
rect 178900 219528 178918 219584
rect 178974 219528 178979 219584
rect 178900 219526 178979 219528
rect 272924 219584 273003 219586
rect 272924 219528 272942 219584
rect 272998 219528 273003 219584
rect 272924 219526 273003 219528
rect 81669 219523 81735 219526
rect 178913 219523 178979 219526
rect 272937 219523 273003 219526
rect 38061 219450 38127 219453
rect 35718 219448 38127 219450
rect 35718 219392 38066 219448
rect 38122 219392 38127 219448
rect 35718 219390 38127 219392
rect 35718 219080 35778 219390
rect 38061 219387 38127 219390
rect 368985 219314 369051 219317
rect 368985 219312 371916 219314
rect 368985 219256 368990 219312
rect 369046 219256 371916 219312
rect 368985 219254 371916 219256
rect 368985 219251 369051 219254
rect 368801 218906 368867 218909
rect 368801 218904 371916 218906
rect 368801 218848 368806 218904
rect 368862 218848 371916 218904
rect 368801 218846 371916 218848
rect 368801 218843 368867 218846
rect 405969 218770 406035 218773
rect 409054 218770 409114 219012
rect 405969 218768 409114 218770
rect 405969 218712 405974 218768
rect 406030 218712 409114 218768
rect 405969 218710 409114 218712
rect 405969 218707 406035 218710
rect 370089 218498 370155 218501
rect 370089 218496 371916 218498
rect 370089 218440 370094 218496
rect 370150 218440 371916 218496
rect 370089 218438 371916 218440
rect 370089 218435 370155 218438
rect 368709 218090 368775 218093
rect 368709 218088 371916 218090
rect 368709 218032 368714 218088
rect 368770 218032 371916 218088
rect 368709 218030 371916 218032
rect 368709 218027 368775 218030
rect 369077 217682 369143 217685
rect 369077 217680 371916 217682
rect 369077 217624 369082 217680
rect 369138 217624 371916 217680
rect 369077 217622 371916 217624
rect 369077 217619 369143 217622
rect 369077 217546 369143 217549
rect 370089 217546 370155 217549
rect 369077 217544 370155 217546
rect 369077 217488 369082 217544
rect 369138 217488 370094 217544
rect 370150 217488 370155 217544
rect 369077 217486 370155 217488
rect 369077 217483 369143 217486
rect 370089 217483 370155 217486
rect 75413 217410 75479 217413
rect 70862 217408 75479 217410
rect 70862 217352 75418 217408
rect 75474 217352 75479 217408
rect 70862 217350 75479 217352
rect 70862 217244 70922 217350
rect 75413 217347 75479 217350
rect 368801 217274 368867 217277
rect 368801 217272 371916 217274
rect 368801 217216 368806 217272
rect 368862 217216 371916 217272
rect 368801 217214 371916 217216
rect 368801 217211 368867 217214
rect 137053 217002 137119 217005
rect 230893 217002 230959 217005
rect 325837 217002 325903 217005
rect 134740 217000 137119 217002
rect 134740 216944 137058 217000
rect 137114 216944 137119 217000
rect 134740 216942 137119 216944
rect 228764 217000 230959 217002
rect 228764 216944 230898 217000
rect 230954 216944 230959 217000
rect 228764 216942 230959 216944
rect 322788 217000 325903 217002
rect 322788 216944 325842 217000
rect 325898 216944 325903 217000
rect 322788 216942 325903 216944
rect 137053 216939 137119 216942
rect 230893 216939 230959 216942
rect 325837 216939 325903 216942
rect 38521 216866 38587 216869
rect 35718 216864 38587 216866
rect 35718 216808 38526 216864
rect 38582 216808 38587 216864
rect 35718 216806 38587 216808
rect 35718 216496 35778 216806
rect 38521 216803 38587 216806
rect 369353 216866 369419 216869
rect 369353 216864 371916 216866
rect 369353 216808 369358 216864
rect 369414 216808 371916 216864
rect 369353 216806 371916 216808
rect 369353 216803 369419 216806
rect 231537 216594 231603 216597
rect 242710 216594 242716 216596
rect 231537 216592 242716 216594
rect 231537 216536 231542 216592
rect 231598 216536 242716 216592
rect 231537 216534 242716 216536
rect 231537 216531 231603 216534
rect 242710 216532 242716 216534
rect 242780 216532 242786 216596
rect 258902 216532 258908 216596
rect 258972 216594 258978 216596
rect 272702 216594 272708 216596
rect 258972 216534 272708 216594
rect 258972 216532 258978 216534
rect 272702 216532 272708 216534
rect 272772 216532 272778 216596
rect 322750 216532 322756 216596
rect 322820 216594 322826 216596
rect 336734 216594 336740 216596
rect 322820 216534 336740 216594
rect 322820 216532 322826 216534
rect 336734 216532 336740 216534
rect 336804 216532 336810 216596
rect 352742 216532 352748 216596
rect 352812 216594 352818 216596
rect 368985 216594 369051 216597
rect 352812 216592 369051 216594
rect 352812 216536 368990 216592
rect 369046 216536 369051 216592
rect 352812 216534 369051 216536
rect 352812 216532 352818 216534
rect 368985 216531 369051 216534
rect 358262 216396 358268 216460
rect 358332 216458 358338 216460
rect 358332 216398 371916 216458
rect 358332 216396 358338 216398
rect 9896 216186 10376 216216
rect 148326 216194 148908 216254
rect 242350 216194 242932 216254
rect 13313 216186 13379 216189
rect 9896 216184 13379 216186
rect 9896 216128 13318 216184
rect 13374 216128 13379 216184
rect 9896 216126 13379 216128
rect 9896 216096 10376 216126
rect 13313 216123 13379 216126
rect 145149 216186 145215 216189
rect 148326 216186 148386 216194
rect 145149 216184 148386 216186
rect 145149 216128 145154 216184
rect 145210 216128 148386 216184
rect 145149 216126 148386 216128
rect 240921 216186 240987 216189
rect 242350 216186 242410 216194
rect 240921 216184 242410 216186
rect 240921 216128 240926 216184
rect 240982 216128 242410 216184
rect 240921 216126 242410 216128
rect 334209 216186 334275 216189
rect 368709 216186 368775 216189
rect 334209 216184 336956 216186
rect 334209 216128 334214 216184
rect 334270 216128 336956 216184
rect 334209 216126 336956 216128
rect 368709 216184 371916 216186
rect 368709 216128 368714 216184
rect 368770 216128 371916 216184
rect 368709 216126 371916 216128
rect 145149 216123 145215 216126
rect 240921 216123 240987 216126
rect 334209 216123 334275 216126
rect 368709 216123 368775 216126
rect 356289 215914 356355 215917
rect 357526 215914 357532 215916
rect 356289 215912 357532 215914
rect 356289 215856 356294 215912
rect 356350 215856 357532 215912
rect 356289 215854 357532 215856
rect 356289 215851 356355 215854
rect 357526 215852 357532 215854
rect 357596 215852 357602 215916
rect 405918 215852 405924 215916
rect 405988 215914 405994 215916
rect 409054 215914 409114 216428
rect 405988 215854 409114 215914
rect 405988 215852 405994 215854
rect 368709 215778 368775 215781
rect 368709 215776 371916 215778
rect 368709 215720 368714 215776
rect 368770 215720 371916 215776
rect 368709 215718 371916 215720
rect 368709 215715 368775 215718
rect 369169 215370 369235 215373
rect 429705 215370 429771 215373
rect 434416 215370 434896 215400
rect 369169 215368 371916 215370
rect 369169 215312 369174 215368
rect 369230 215312 371916 215368
rect 369169 215310 371916 215312
rect 429705 215368 434896 215370
rect 429705 215312 429710 215368
rect 429766 215312 434896 215368
rect 429705 215310 434896 215312
rect 369169 215307 369235 215310
rect 429705 215307 429771 215310
rect 434416 215280 434896 215310
rect 51401 215234 51467 215237
rect 356197 215234 356263 215237
rect 428693 215234 428759 215237
rect 51401 215232 55068 215234
rect 16073 214554 16139 214557
rect 20078 214554 20138 215204
rect 51401 215176 51406 215232
rect 51462 215176 55068 215232
rect 51401 215174 55068 215176
rect 352780 215232 356263 215234
rect 352780 215176 356202 215232
rect 356258 215176 356263 215232
rect 352780 215174 356263 215176
rect 424724 215232 428759 215234
rect 424724 215176 428698 215232
rect 428754 215176 428759 215232
rect 424724 215174 428759 215176
rect 51401 215171 51467 215174
rect 356197 215171 356263 215174
rect 428693 215171 428759 215174
rect 368709 214962 368775 214965
rect 368709 214960 371916 214962
rect 368709 214904 368714 214960
rect 368770 214904 371916 214960
rect 368709 214902 371916 214904
rect 368709 214899 368775 214902
rect 16073 214552 20138 214554
rect 16073 214496 16078 214552
rect 16134 214496 20138 214552
rect 16073 214494 20138 214496
rect 368801 214554 368867 214557
rect 368801 214552 371916 214554
rect 368801 214496 368806 214552
rect 368862 214496 371916 214552
rect 368801 214494 371916 214496
rect 16073 214491 16139 214494
rect 368801 214491 368867 214494
rect 38521 214282 38587 214285
rect 35718 214280 38587 214282
rect 35718 214224 38526 214280
rect 38582 214224 38587 214280
rect 35718 214222 38587 214224
rect 35718 214048 35778 214222
rect 38521 214219 38587 214222
rect 368893 214146 368959 214149
rect 405969 214146 406035 214149
rect 368893 214144 371916 214146
rect 368893 214088 368898 214144
rect 368954 214088 371916 214144
rect 368893 214086 371916 214088
rect 405969 214144 408930 214146
rect 405969 214088 405974 214144
rect 406030 214088 408930 214144
rect 405969 214086 408930 214088
rect 368893 214083 368959 214086
rect 405969 214083 406035 214086
rect 408870 213980 408930 214086
rect 136869 213874 136935 213877
rect 231721 213874 231787 213877
rect 324917 213874 324983 213877
rect 134740 213872 136935 213874
rect 134740 213816 136874 213872
rect 136930 213816 136935 213872
rect 134740 213814 136935 213816
rect 228764 213872 231787 213874
rect 228764 213816 231726 213872
rect 231782 213816 231787 213872
rect 228764 213814 231787 213816
rect 322788 213872 324983 213874
rect 322788 213816 324922 213872
rect 324978 213816 324983 213872
rect 322788 213814 324983 213816
rect 136869 213811 136935 213814
rect 231721 213811 231787 213814
rect 324917 213811 324983 213814
rect 73430 213738 73436 213740
rect 70862 213678 73436 213738
rect 70862 213572 70922 213678
rect 73430 213676 73436 213678
rect 73500 213676 73506 213740
rect 368709 213738 368775 213741
rect 368709 213736 371916 213738
rect 368709 213680 368714 213736
rect 368770 213680 371916 213736
rect 368709 213678 371916 213680
rect 368709 213675 368775 213678
rect 367973 213330 368039 213333
rect 367973 213328 371916 213330
rect 367973 213272 367978 213328
rect 368034 213272 371916 213328
rect 367973 213270 371916 213272
rect 367973 213267 368039 213270
rect 368709 213058 368775 213061
rect 368709 213056 371916 213058
rect 368709 213000 368714 213056
rect 368770 213000 371916 213056
rect 368709 212998 371916 213000
rect 368709 212995 368775 212998
rect 167873 212786 167939 212789
rect 261713 212786 261779 212789
rect 164732 212784 167939 212786
rect 164732 212728 167878 212784
rect 167934 212728 167939 212784
rect 164732 212726 167939 212728
rect 258756 212784 261779 212786
rect 258756 212728 261718 212784
rect 261774 212728 261779 212784
rect 258756 212726 261779 212728
rect 167873 212723 167939 212726
rect 261713 212723 261779 212726
rect 358405 211698 358471 211701
rect 358589 211698 358655 211701
rect 358405 211696 358655 211698
rect 358405 211640 358410 211696
rect 358466 211640 358594 211696
rect 358650 211640 358655 211696
rect 358405 211638 358655 211640
rect 358405 211635 358471 211638
rect 358589 211635 358655 211638
rect 38705 211562 38771 211565
rect 35748 211560 38771 211562
rect 35748 211504 38710 211560
rect 38766 211504 38771 211560
rect 35748 211502 38771 211504
rect 38705 211499 38771 211502
rect 54069 211018 54135 211021
rect 54662 211018 54668 211020
rect 54069 211016 54668 211018
rect 54069 210960 54074 211016
rect 54130 210960 54668 211016
rect 54069 210958 54668 210960
rect 54069 210955 54135 210958
rect 54662 210956 54668 210958
rect 54732 210956 54738 211020
rect 405969 211018 406035 211021
rect 409054 211018 409114 211532
rect 405969 211016 409114 211018
rect 405969 210960 405974 211016
rect 406030 210960 409114 211016
rect 405969 210958 409114 210960
rect 405969 210955 406035 210958
rect 136961 210746 137027 210749
rect 231629 210746 231695 210749
rect 325653 210746 325719 210749
rect 134740 210744 137027 210746
rect 134740 210688 136966 210744
rect 137022 210688 137027 210744
rect 134740 210686 137027 210688
rect 228764 210744 231695 210746
rect 228764 210688 231634 210744
rect 231690 210688 231695 210744
rect 228764 210686 231695 210688
rect 322788 210744 325719 210746
rect 322788 210688 325658 210744
rect 325714 210688 325719 210744
rect 322788 210686 325719 210688
rect 136961 210683 137027 210686
rect 231629 210683 231695 210686
rect 325653 210683 325719 210686
rect 51401 210202 51467 210205
rect 74677 210202 74743 210205
rect 356197 210202 356263 210205
rect 427313 210202 427379 210205
rect 51401 210200 55068 210202
rect 17545 209658 17611 209661
rect 20078 209658 20138 210172
rect 51401 210144 51406 210200
rect 51462 210144 55068 210200
rect 51401 210142 55068 210144
rect 70862 210200 74743 210202
rect 70862 210144 74682 210200
rect 74738 210144 74743 210200
rect 70862 210142 74743 210144
rect 352780 210200 356263 210202
rect 352780 210144 356202 210200
rect 356258 210144 356263 210200
rect 352780 210142 356263 210144
rect 424724 210200 427379 210202
rect 424724 210144 427318 210200
rect 427374 210144 427379 210200
rect 424724 210142 427379 210144
rect 51401 210139 51467 210142
rect 70862 210066 70922 210142
rect 74677 210139 74743 210142
rect 356197 210139 356263 210142
rect 427313 210139 427379 210142
rect 70708 210036 70922 210066
rect 17545 209656 20138 209658
rect 17545 209600 17550 209656
rect 17606 209600 20138 209656
rect 17545 209598 20138 209600
rect 70678 210006 70892 210036
rect 17545 209595 17611 209598
rect 70678 209522 70738 210006
rect 70813 209522 70879 209525
rect 70678 209520 70879 209522
rect 70678 209464 70818 209520
rect 70874 209464 70879 209520
rect 70678 209462 70879 209464
rect 70813 209459 70879 209462
rect 405969 209522 406035 209525
rect 405969 209520 408930 209522
rect 405969 209464 405974 209520
rect 406030 209464 408930 209520
rect 405969 209462 408930 209464
rect 405969 209459 406035 209462
rect 38521 209250 38587 209253
rect 35718 209248 38587 209250
rect 35718 209192 38526 209248
rect 38582 209192 38587 209248
rect 35718 209190 38587 209192
rect 35718 209016 35778 209190
rect 38521 209187 38587 209190
rect 16257 208978 16323 208981
rect 17545 208978 17611 208981
rect 16257 208976 17611 208978
rect 16257 208920 16262 208976
rect 16318 208920 17550 208976
rect 17606 208920 17611 208976
rect 408870 208948 408930 209462
rect 16257 208918 17611 208920
rect 16257 208915 16323 208918
rect 17545 208915 17611 208918
rect 138157 208298 138223 208301
rect 147030 208298 147036 208300
rect 134710 208296 147036 208298
rect 134710 208240 138162 208296
rect 138218 208240 147036 208296
rect 134710 208238 147036 208240
rect 134710 207588 134770 208238
rect 138157 208235 138223 208238
rect 147030 208236 147036 208238
rect 147100 208236 147106 208300
rect 231445 207754 231511 207757
rect 242209 207754 242275 207757
rect 228734 207752 242275 207754
rect 228734 207696 231450 207752
rect 231506 207696 242214 207752
rect 242270 207696 242275 207752
rect 228734 207694 242275 207696
rect 228734 207588 228794 207694
rect 231445 207691 231511 207694
rect 242209 207691 242275 207694
rect 325469 207618 325535 207621
rect 322788 207616 325535 207618
rect 322788 207560 325474 207616
rect 325530 207560 325535 207616
rect 322788 207558 325535 207560
rect 325469 207555 325535 207558
rect 51401 206802 51467 206805
rect 52638 206802 52644 206804
rect 51401 206800 52644 206802
rect 51401 206744 51406 206800
rect 51462 206744 52644 206800
rect 51401 206742 52644 206744
rect 51401 206739 51467 206742
rect 52638 206740 52644 206742
rect 52708 206740 52714 206804
rect 405969 206802 406035 206805
rect 405969 206800 408930 206802
rect 405969 206744 405974 206800
rect 406030 206744 408930 206800
rect 405969 206742 408930 206744
rect 405969 206739 406035 206742
rect 38521 206666 38587 206669
rect 35718 206664 38587 206666
rect 35718 206608 38526 206664
rect 38582 206608 38587 206664
rect 35718 206606 38587 206608
rect 35718 206568 35778 206606
rect 38521 206603 38587 206606
rect 74125 206530 74191 206533
rect 70862 206528 74191 206530
rect 70862 206472 74130 206528
rect 74186 206472 74191 206528
rect 408870 206500 408930 206742
rect 70862 206470 74191 206472
rect 70862 206364 70922 206470
rect 74125 206467 74191 206470
rect 51401 205306 51467 205309
rect 356197 205306 356263 205309
rect 427497 205306 427563 205309
rect 51401 205304 55068 205306
rect 16349 204898 16415 204901
rect 20078 204898 20138 205276
rect 51401 205248 51406 205304
rect 51462 205248 55068 205304
rect 51401 205246 55068 205248
rect 352780 205304 356263 205306
rect 352780 205248 356202 205304
rect 356258 205248 356263 205304
rect 352780 205246 356263 205248
rect 424724 205304 427563 205306
rect 424724 205248 427502 205304
rect 427558 205248 427563 205304
rect 424724 205246 427563 205248
rect 51401 205243 51467 205246
rect 356197 205243 356263 205246
rect 427497 205243 427563 205246
rect 73849 205036 73915 205037
rect 73798 205034 73804 205036
rect 73758 204974 73804 205034
rect 73868 205032 73915 205036
rect 73910 204976 73915 205032
rect 73798 204972 73804 204974
rect 73868 204972 73915 204976
rect 73849 204971 73915 204972
rect 16349 204896 20138 204898
rect 16349 204840 16354 204896
rect 16410 204840 20138 204896
rect 16349 204838 20138 204840
rect 16349 204835 16415 204838
rect 73798 204836 73804 204900
rect 73868 204898 73874 204900
rect 74125 204898 74191 204901
rect 73868 204896 74191 204898
rect 73868 204840 74130 204896
rect 74186 204840 74191 204896
rect 73868 204838 74191 204840
rect 73868 204836 73874 204838
rect 74125 204835 74191 204838
rect 74401 204898 74467 204901
rect 74534 204898 74540 204900
rect 74401 204896 74540 204898
rect 74401 204840 74406 204896
rect 74462 204840 74540 204896
rect 74401 204838 74540 204840
rect 74401 204835 74467 204838
rect 74534 204836 74540 204838
rect 74604 204836 74610 204900
rect 134702 204836 134708 204900
rect 134772 204836 134778 204900
rect 70813 204762 70879 204765
rect 72142 204762 72148 204764
rect 70813 204760 72148 204762
rect 70813 204704 70818 204760
rect 70874 204704 72148 204760
rect 70813 204702 72148 204704
rect 70813 204699 70879 204702
rect 72142 204700 72148 204702
rect 72212 204700 72218 204764
rect 73849 204762 73915 204765
rect 73982 204762 73988 204764
rect 73849 204760 73988 204762
rect 73849 204704 73854 204760
rect 73910 204704 73988 204760
rect 73849 204702 73988 204704
rect 73849 204699 73915 204702
rect 73982 204700 73988 204702
rect 74052 204700 74058 204764
rect 74401 204762 74467 204765
rect 74534 204762 74540 204764
rect 74401 204760 74540 204762
rect 74401 204704 74406 204760
rect 74462 204704 74540 204760
rect 74401 204702 74540 204704
rect 74401 204699 74467 204702
rect 74534 204700 74540 204702
rect 74604 204700 74610 204764
rect 134710 204762 134770 204836
rect 136869 204762 136935 204765
rect 134710 204760 136935 204762
rect 134710 204704 136874 204760
rect 136930 204704 136935 204760
rect 134710 204702 136935 204704
rect 38521 204490 38587 204493
rect 35718 204488 38587 204490
rect 35718 204432 38526 204488
rect 38582 204432 38587 204488
rect 35718 204430 38587 204432
rect 35718 204120 35778 204430
rect 38521 204427 38587 204430
rect 73614 204428 73620 204492
rect 73684 204490 73690 204492
rect 84654 204490 84660 204492
rect 73684 204430 84660 204490
rect 73684 204428 73690 204430
rect 84654 204428 84660 204430
rect 84724 204428 84730 204492
rect 134710 204460 134770 204702
rect 136869 204699 136935 204702
rect 242209 204626 242275 204629
rect 242710 204626 242716 204628
rect 242209 204624 242716 204626
rect 242209 204568 242214 204624
rect 242270 204568 242716 204624
rect 242209 204566 242716 204568
rect 242209 204563 242275 204566
rect 242710 204564 242716 204566
rect 242780 204564 242786 204628
rect 406061 204626 406127 204629
rect 406061 204624 408930 204626
rect 406061 204568 406066 204624
rect 406122 204568 408930 204624
rect 406061 204566 408930 204568
rect 406061 204563 406127 204566
rect 325561 204490 325627 204493
rect 322788 204488 325627 204490
rect 322788 204460 325566 204488
rect 322758 204432 325566 204460
rect 325622 204432 325627 204488
rect 322758 204430 325627 204432
rect 228734 204354 228794 204392
rect 231629 204354 231695 204357
rect 228734 204352 231695 204354
rect 228734 204296 231634 204352
rect 231690 204296 231695 204352
rect 228734 204294 231695 204296
rect 231629 204291 231695 204294
rect 237374 204292 237380 204356
rect 237444 204354 237450 204356
rect 237517 204354 237583 204357
rect 239582 204354 239588 204356
rect 237444 204352 239588 204354
rect 237444 204296 237522 204352
rect 237578 204296 239588 204352
rect 237444 204294 239588 204296
rect 237444 204292 237450 204294
rect 237517 204291 237583 204294
rect 239582 204292 239588 204294
rect 239652 204292 239658 204356
rect 322758 204220 322818 204430
rect 325561 204427 325627 204430
rect 322750 204156 322756 204220
rect 322820 204156 322826 204220
rect 408870 204052 408930 204566
rect 73614 203476 73620 203540
rect 73684 203538 73690 203540
rect 74125 203538 74191 203541
rect 73684 203536 74191 203538
rect 73684 203480 74130 203536
rect 74186 203480 74191 203536
rect 73684 203478 74191 203480
rect 73684 203476 73690 203478
rect 74125 203475 74191 203478
rect 9896 202858 10376 202888
rect 148326 202866 148908 202926
rect 242350 202866 242932 202926
rect 13957 202858 14023 202861
rect 9896 202856 14023 202858
rect 9896 202800 13962 202856
rect 14018 202800 14023 202856
rect 9896 202798 14023 202800
rect 9896 202768 10376 202798
rect 13957 202795 14023 202798
rect 81669 202858 81735 202861
rect 145149 202858 145215 202861
rect 148326 202858 148386 202866
rect 178913 202858 178979 202861
rect 81669 202856 85060 202858
rect 81669 202800 81674 202856
rect 81730 202800 85060 202856
rect 81669 202798 85060 202800
rect 145149 202856 148386 202858
rect 145149 202800 145154 202856
rect 145210 202800 148386 202856
rect 145149 202798 148386 202800
rect 178900 202856 178979 202858
rect 178900 202800 178918 202856
rect 178974 202800 178979 202856
rect 178900 202798 178979 202800
rect 81669 202795 81735 202798
rect 145149 202795 145215 202798
rect 178913 202795 178979 202798
rect 240369 202858 240435 202861
rect 242350 202858 242410 202866
rect 272937 202858 273003 202861
rect 240369 202856 242410 202858
rect 240369 202800 240374 202856
rect 240430 202800 242410 202856
rect 240369 202798 242410 202800
rect 272924 202856 273003 202858
rect 272924 202800 272942 202856
rect 272998 202800 273003 202856
rect 272924 202798 273003 202800
rect 240369 202795 240435 202798
rect 272937 202795 273003 202798
rect 334209 202858 334275 202861
rect 430073 202858 430139 202861
rect 434416 202858 434896 202888
rect 334209 202856 336956 202858
rect 334209 202800 334214 202856
rect 334270 202800 336956 202856
rect 334209 202798 336956 202800
rect 430073 202856 434896 202858
rect 430073 202800 430078 202856
rect 430134 202800 434896 202856
rect 430073 202798 434896 202800
rect 334209 202795 334275 202798
rect 430073 202795 430139 202798
rect 434416 202768 434896 202798
rect 70678 202178 70738 202692
rect 73614 202178 73620 202180
rect 70678 202118 73620 202178
rect 73614 202116 73620 202118
rect 73684 202178 73690 202180
rect 74350 202178 74356 202180
rect 73684 202118 74356 202178
rect 73684 202116 73690 202118
rect 74350 202116 74356 202118
rect 74420 202116 74426 202180
rect 242577 202042 242643 202045
rect 242710 202042 242716 202044
rect 242577 202040 242716 202042
rect 242577 201984 242582 202040
rect 242638 201984 242716 202040
rect 242577 201982 242716 201984
rect 242577 201979 242643 201982
rect 242710 201980 242716 201982
rect 242780 201980 242786 202044
rect 38521 201498 38587 201501
rect 35748 201496 38587 201498
rect 35748 201440 38526 201496
rect 38582 201440 38587 201496
rect 35748 201438 38587 201440
rect 38521 201435 38587 201438
rect 405969 201362 406035 201365
rect 409054 201362 409114 201468
rect 405969 201360 409114 201362
rect 134710 200954 134770 201264
rect 228734 200956 228794 201264
rect 322758 200956 322818 201332
rect 405969 201304 405974 201360
rect 406030 201304 409114 201360
rect 405969 201302 409114 201304
rect 405969 201299 406035 201302
rect 136910 200954 136916 200956
rect 134710 200894 136916 200954
rect 136910 200892 136916 200894
rect 136980 200892 136986 200956
rect 228726 200954 228732 200956
rect 228604 200894 228732 200954
rect 228726 200892 228732 200894
rect 228796 200892 228802 200956
rect 322750 200892 322756 200956
rect 322820 200892 322826 200956
rect 228734 200682 228794 200892
rect 230801 200682 230867 200685
rect 228734 200680 230867 200682
rect 228734 200624 230806 200680
rect 230862 200624 230867 200680
rect 228734 200622 230867 200624
rect 230801 200619 230867 200622
rect 51217 200274 51283 200277
rect 356197 200274 356263 200277
rect 427129 200274 427195 200277
rect 51217 200272 55068 200274
rect 17637 199730 17703 199733
rect 20078 199730 20138 200244
rect 51217 200216 51222 200272
rect 51278 200216 55068 200272
rect 51217 200214 55068 200216
rect 352780 200272 356263 200274
rect 352780 200216 356202 200272
rect 356258 200216 356263 200272
rect 352780 200214 356263 200216
rect 424724 200272 427195 200274
rect 424724 200216 427134 200272
rect 427190 200216 427195 200272
rect 424724 200214 427195 200216
rect 51217 200211 51283 200214
rect 356197 200211 356263 200214
rect 427129 200211 427195 200214
rect 17637 199728 20138 199730
rect 17637 199672 17642 199728
rect 17698 199672 20138 199728
rect 17637 199670 20138 199672
rect 17637 199667 17703 199670
rect 38521 199186 38587 199189
rect 74534 199186 74540 199188
rect 35718 199184 38587 199186
rect 35718 199128 38526 199184
rect 38582 199128 38587 199184
rect 35718 199126 38587 199128
rect 35718 199088 35778 199126
rect 38521 199123 38587 199126
rect 70862 199126 74540 199186
rect 70862 199020 70922 199126
rect 74534 199124 74540 199126
rect 74604 199124 74610 199188
rect 405969 199186 406035 199189
rect 405969 199184 408930 199186
rect 405969 199128 405974 199184
rect 406030 199128 408930 199184
rect 405969 199126 408930 199128
rect 405969 199123 406035 199126
rect 408870 199020 408930 199126
rect 164878 198852 164884 198916
rect 164948 198914 164954 198916
rect 176654 198914 176660 198916
rect 164948 198854 176660 198914
rect 164948 198852 164954 198854
rect 176654 198852 176660 198854
rect 176724 198852 176730 198916
rect 322750 198716 322756 198780
rect 322820 198778 322826 198780
rect 324549 198778 324615 198781
rect 322820 198776 324615 198778
rect 322820 198720 324554 198776
rect 324610 198720 324615 198776
rect 322820 198718 324615 198720
rect 322820 198716 322826 198718
rect 136910 198234 136916 198236
rect 134740 198174 136916 198234
rect 136910 198172 136916 198174
rect 136980 198172 136986 198236
rect 322758 198204 322818 198716
rect 324549 198715 324615 198718
rect 228734 197554 228794 198136
rect 230709 197556 230775 197557
rect 230709 197554 230756 197556
rect 228734 197552 230756 197554
rect 230820 197554 230826 197556
rect 228734 197496 230714 197552
rect 228734 197494 230756 197496
rect 230709 197492 230756 197494
rect 230820 197494 230902 197554
rect 230820 197492 230826 197494
rect 261110 197492 261116 197556
rect 261180 197554 261186 197556
rect 270494 197554 270500 197556
rect 261180 197494 270500 197554
rect 261180 197492 261186 197494
rect 270494 197492 270500 197494
rect 270564 197492 270570 197556
rect 230709 197491 230775 197492
rect 38521 196466 38587 196469
rect 35748 196464 38587 196466
rect 35748 196408 38526 196464
rect 38582 196408 38587 196464
rect 35748 196406 38587 196408
rect 38521 196403 38587 196406
rect 405969 195922 406035 195925
rect 409054 195922 409114 196436
rect 405969 195920 409114 195922
rect 405969 195864 405974 195920
rect 406030 195864 409114 195920
rect 405969 195862 409114 195864
rect 405969 195859 406035 195862
rect 17453 195378 17519 195381
rect 17453 195376 19954 195378
rect 17453 195320 17458 195376
rect 17514 195320 19954 195376
rect 17453 195318 19954 195320
rect 17453 195315 17519 195318
rect 19894 195212 19954 195318
rect 51309 195242 51375 195245
rect 70678 195242 70738 195484
rect 74217 195244 74283 195245
rect 74166 195242 74172 195244
rect 51309 195240 55068 195242
rect 51309 195184 51314 195240
rect 51370 195184 55068 195240
rect 51309 195182 55068 195184
rect 70678 195182 74172 195242
rect 74236 195242 74283 195244
rect 74493 195244 74559 195245
rect 74493 195242 74540 195244
rect 74236 195240 74328 195242
rect 74278 195184 74328 195240
rect 51309 195179 51375 195182
rect 74166 195180 74172 195182
rect 74236 195182 74328 195184
rect 74448 195240 74540 195242
rect 74448 195184 74498 195240
rect 74448 195182 74540 195184
rect 74236 195180 74283 195182
rect 74217 195179 74283 195180
rect 74493 195180 74540 195182
rect 74604 195180 74610 195244
rect 356197 195242 356263 195245
rect 427589 195242 427655 195245
rect 352780 195240 356263 195242
rect 352780 195184 356202 195240
rect 356258 195184 356263 195240
rect 352780 195182 356263 195184
rect 424724 195240 427655 195242
rect 424724 195184 427594 195240
rect 427650 195184 427655 195240
rect 424724 195182 427655 195184
rect 74493 195179 74559 195180
rect 356197 195179 356263 195182
rect 427589 195179 427655 195182
rect 74217 195106 74283 195109
rect 74493 195108 74559 195109
rect 74350 195106 74356 195108
rect 74217 195104 74356 195106
rect 74217 195048 74222 195104
rect 74278 195048 74356 195104
rect 74217 195046 74356 195048
rect 74217 195043 74283 195046
rect 74350 195044 74356 195046
rect 74420 195044 74426 195108
rect 74493 195104 74540 195108
rect 74604 195106 74610 195108
rect 74493 195048 74498 195104
rect 74493 195044 74540 195048
rect 74604 195046 74650 195106
rect 74604 195044 74610 195046
rect 74493 195043 74559 195044
rect 134710 194698 134770 195008
rect 228734 194970 228794 195008
rect 230750 194970 230756 194972
rect 228734 194910 230756 194970
rect 230750 194908 230756 194910
rect 230820 194970 230826 194972
rect 230893 194970 230959 194973
rect 231077 194970 231143 194973
rect 230820 194968 231143 194970
rect 230820 194912 230898 194968
rect 230954 194912 231082 194968
rect 231138 194912 231143 194968
rect 230820 194910 231143 194912
rect 230820 194908 230826 194910
rect 230893 194907 230959 194910
rect 231077 194907 231143 194910
rect 138014 194698 138020 194700
rect 134710 194638 138020 194698
rect 138014 194636 138020 194638
rect 138084 194636 138090 194700
rect 38797 194562 38863 194565
rect 322758 194564 322818 195076
rect 35718 194560 38863 194562
rect 35718 194504 38802 194560
rect 38858 194504 38863 194560
rect 35718 194502 38863 194504
rect 35718 194056 35778 194502
rect 38797 194499 38863 194502
rect 322750 194500 322756 194564
rect 322820 194500 322826 194564
rect 406061 194562 406127 194565
rect 406061 194560 408930 194562
rect 406061 194504 406066 194560
rect 406122 194504 408930 194560
rect 406061 194502 408930 194504
rect 406061 194499 406127 194502
rect 408870 193988 408930 194502
rect 167965 192794 168031 192797
rect 262357 192794 262423 192797
rect 164732 192792 168031 192794
rect 164732 192736 167970 192792
rect 168026 192736 168031 192792
rect 164732 192734 168031 192736
rect 258756 192792 262423 192794
rect 258756 192736 262362 192792
rect 262418 192736 262423 192792
rect 258756 192734 262423 192736
rect 167965 192731 168031 192734
rect 262357 192731 262423 192734
rect 72326 192596 72332 192660
rect 72396 192658 72402 192660
rect 72396 192598 72762 192658
rect 72396 192596 72402 192598
rect 72702 192524 72762 192598
rect 242577 192524 242643 192525
rect 72694 192460 72700 192524
rect 72764 192460 72770 192524
rect 242526 192522 242532 192524
rect 242486 192462 242532 192522
rect 242596 192520 242643 192524
rect 242638 192464 242643 192520
rect 242526 192460 242532 192462
rect 242596 192460 242643 192464
rect 242577 192459 242643 192460
rect 137605 191978 137671 191981
rect 231537 191978 231603 191981
rect 325377 191978 325443 191981
rect 134740 191976 137671 191978
rect 134740 191920 137610 191976
rect 137666 191920 137671 191976
rect 134740 191918 137671 191920
rect 228764 191976 231603 191978
rect 228764 191920 231542 191976
rect 231598 191920 231603 191976
rect 228764 191918 231603 191920
rect 322788 191976 325443 191978
rect 322788 191920 325382 191976
rect 325438 191920 325443 191976
rect 322788 191918 325443 191920
rect 137605 191915 137671 191918
rect 231537 191915 231603 191918
rect 325377 191915 325443 191918
rect 38797 191570 38863 191573
rect 35748 191568 38863 191570
rect 35748 191512 38802 191568
rect 38858 191512 38863 191568
rect 35748 191510 38863 191512
rect 38797 191507 38863 191510
rect 70678 191298 70738 191812
rect 405969 191706 406035 191709
rect 405969 191704 408930 191706
rect 405969 191648 405974 191704
rect 406030 191648 408930 191704
rect 405969 191646 408930 191648
rect 405969 191643 406035 191646
rect 408870 191540 408930 191646
rect 352793 191436 352859 191437
rect 352742 191372 352748 191436
rect 352812 191434 352859 191436
rect 352812 191432 352904 191434
rect 352854 191376 352904 191432
rect 352812 191374 352904 191376
rect 352812 191372 352859 191374
rect 352793 191371 352859 191372
rect 73982 191298 73988 191300
rect 70678 191238 73988 191298
rect 73982 191236 73988 191238
rect 74052 191236 74058 191300
rect 434416 190346 434896 190376
rect 424694 190286 434896 190346
rect 424694 190248 424754 190286
rect 434416 190256 434896 190286
rect 51217 190210 51283 190213
rect 356197 190210 356263 190213
rect 51217 190208 55068 190210
rect 16441 189666 16507 189669
rect 20078 189666 20138 190180
rect 51217 190152 51222 190208
rect 51278 190152 55068 190208
rect 51217 190150 55068 190152
rect 352780 190208 356263 190210
rect 352780 190152 356202 190208
rect 356258 190152 356263 190208
rect 352780 190150 356263 190152
rect 51217 190147 51283 190150
rect 356197 190147 356263 190150
rect 16441 189664 20138 189666
rect 16441 189608 16446 189664
rect 16502 189608 20138 189664
rect 16441 189606 20138 189608
rect 16441 189603 16507 189606
rect 148326 189538 148908 189598
rect 242350 189538 242932 189598
rect 145609 189530 145675 189533
rect 148326 189530 148386 189538
rect 145609 189528 148386 189530
rect 145609 189472 145614 189528
rect 145670 189472 148386 189528
rect 145609 189470 148386 189472
rect 240369 189530 240435 189533
rect 242350 189530 242410 189538
rect 240369 189528 242410 189530
rect 240369 189472 240374 189528
rect 240430 189472 242410 189528
rect 240369 189470 242410 189472
rect 334209 189530 334275 189533
rect 405969 189530 406035 189533
rect 334209 189528 336956 189530
rect 334209 189472 334214 189528
rect 334270 189472 336956 189528
rect 334209 189470 336956 189472
rect 405969 189528 408930 189530
rect 405969 189472 405974 189528
rect 406030 189472 408930 189528
rect 405969 189470 408930 189472
rect 145609 189467 145675 189470
rect 240369 189467 240435 189470
rect 334209 189467 334275 189470
rect 405969 189467 406035 189470
rect 9896 189394 10376 189424
rect 13313 189394 13379 189397
rect 9896 189392 13379 189394
rect 9896 189336 13318 189392
rect 13374 189336 13379 189392
rect 9896 189334 13379 189336
rect 9896 189304 10376 189334
rect 13313 189331 13379 189334
rect 38061 189258 38127 189261
rect 35718 189256 38127 189258
rect 35718 189200 38066 189256
rect 38122 189200 38127 189256
rect 35718 189198 38127 189200
rect 35718 189024 35778 189198
rect 38061 189195 38127 189198
rect 408870 188956 408930 189470
rect 231997 188850 232063 188853
rect 324549 188850 324615 188853
rect 228764 188848 232063 188850
rect 228764 188792 232002 188848
rect 232058 188792 232063 188848
rect 228764 188790 232063 188792
rect 322788 188848 324615 188850
rect 322788 188792 324554 188848
rect 324610 188792 324615 188848
rect 322788 188790 324615 188792
rect 231997 188787 232063 188790
rect 324549 188787 324615 188790
rect 134710 188578 134770 188752
rect 137789 188578 137855 188581
rect 134710 188576 137855 188578
rect 134710 188520 137794 188576
rect 137850 188520 137855 188576
rect 134710 188518 137855 188520
rect 137789 188515 137855 188518
rect 70678 188034 70738 188140
rect 74125 188034 74191 188037
rect 70678 188032 74191 188034
rect 70678 187976 74130 188032
rect 74186 187976 74191 188032
rect 70678 187974 74191 187976
rect 74125 187971 74191 187974
rect 38061 186538 38127 186541
rect 35748 186536 38127 186538
rect 35748 186480 38066 186536
rect 38122 186480 38127 186536
rect 35748 186478 38127 186480
rect 38061 186475 38127 186478
rect 81669 186266 81735 186269
rect 178913 186266 178979 186269
rect 273121 186266 273187 186269
rect 81669 186264 85060 186266
rect 81669 186208 81674 186264
rect 81730 186208 85060 186264
rect 81669 186206 85060 186208
rect 178900 186264 178979 186266
rect 178900 186208 178918 186264
rect 178974 186208 178979 186264
rect 178900 186206 178979 186208
rect 273108 186264 273187 186266
rect 273108 186208 273126 186264
rect 273182 186208 273187 186264
rect 273108 186206 273187 186208
rect 81669 186203 81735 186206
rect 178913 186203 178979 186206
rect 273121 186203 273187 186206
rect 405969 186266 406035 186269
rect 409054 186266 409114 186508
rect 405969 186264 409114 186266
rect 405969 186208 405974 186264
rect 406030 186208 409114 186264
rect 405969 186206 409114 186208
rect 405969 186203 406035 186206
rect 74309 185722 74375 185725
rect 74534 185722 74540 185724
rect 74309 185720 74540 185722
rect 74309 185664 74314 185720
rect 74370 185664 74540 185720
rect 74309 185662 74540 185664
rect 74309 185659 74375 185662
rect 74534 185660 74540 185662
rect 74604 185660 74610 185724
rect 137329 185722 137395 185725
rect 231353 185722 231419 185725
rect 325285 185722 325351 185725
rect 134740 185720 137395 185722
rect 134740 185664 137334 185720
rect 137390 185664 137395 185720
rect 134740 185662 137395 185664
rect 228764 185720 231419 185722
rect 228764 185664 231358 185720
rect 231414 185664 231419 185720
rect 228764 185662 231419 185664
rect 322788 185720 325351 185722
rect 322788 185664 325290 185720
rect 325346 185664 325351 185720
rect 322788 185662 325351 185664
rect 137329 185659 137395 185662
rect 231353 185659 231419 185662
rect 325285 185659 325351 185662
rect 73941 185588 74007 185589
rect 73941 185584 73988 185588
rect 74052 185586 74058 185588
rect 74217 185586 74283 185589
rect 74534 185586 74540 185588
rect 73941 185528 73946 185584
rect 73941 185524 73988 185528
rect 74052 185526 74098 185586
rect 74217 185584 74540 185586
rect 74217 185528 74222 185584
rect 74278 185528 74540 185584
rect 74217 185526 74540 185528
rect 74052 185524 74058 185526
rect 73941 185523 74007 185524
rect 74217 185523 74283 185526
rect 74534 185524 74540 185526
rect 74604 185524 74610 185588
rect 17453 185450 17519 185453
rect 73941 185452 74007 185453
rect 73941 185450 73988 185452
rect 17453 185448 19954 185450
rect 17453 185392 17458 185448
rect 17514 185392 19954 185448
rect 17453 185390 19954 185392
rect 73896 185448 73988 185450
rect 73896 185392 73946 185448
rect 73896 185390 73988 185392
rect 17453 185387 17519 185390
rect 19894 185284 19954 185390
rect 73941 185388 73988 185390
rect 74052 185388 74058 185452
rect 427221 185450 427287 185453
rect 424694 185448 427287 185450
rect 424694 185392 427226 185448
rect 427282 185392 427287 185448
rect 424694 185390 427287 185392
rect 73941 185387 74007 185388
rect 424694 185352 424754 185390
rect 427221 185387 427287 185390
rect 51401 185314 51467 185317
rect 51401 185312 55068 185314
rect 51401 185256 51406 185312
rect 51462 185256 55068 185312
rect 51401 185254 55068 185256
rect 51401 185251 51467 185254
rect 71958 185252 71964 185316
rect 72028 185314 72034 185316
rect 72694 185314 72700 185316
rect 72028 185254 72700 185314
rect 72028 185252 72034 185254
rect 72694 185252 72700 185254
rect 72764 185252 72770 185316
rect 356197 185314 356263 185317
rect 352780 185312 356263 185314
rect 352780 185256 356202 185312
rect 356258 185256 356263 185312
rect 352780 185254 356263 185256
rect 356197 185251 356263 185254
rect 74033 185042 74099 185045
rect 70862 185040 74099 185042
rect 70862 184984 74038 185040
rect 74094 184984 74099 185040
rect 70862 184982 74099 184984
rect 70862 184604 70922 184982
rect 74033 184979 74099 184982
rect 38797 184090 38863 184093
rect 35748 184088 38863 184090
rect 35748 184032 38802 184088
rect 38858 184032 38863 184088
rect 35748 184030 38863 184032
rect 38797 184027 38863 184030
rect 351638 184028 351644 184092
rect 351708 184090 351714 184092
rect 352793 184090 352859 184093
rect 351708 184088 352859 184090
rect 351708 184032 352798 184088
rect 352854 184032 352859 184088
rect 351708 184030 352859 184032
rect 351708 184028 351714 184030
rect 352793 184027 352859 184030
rect 405969 183954 406035 183957
rect 409054 183954 409114 184060
rect 405969 183952 409114 183954
rect 405969 183896 405974 183952
rect 406030 183896 409114 183952
rect 405969 183894 409114 183896
rect 405969 183891 406035 183894
rect 242710 183076 242716 183140
rect 242780 183138 242786 183140
rect 248925 183138 248991 183141
rect 242780 183136 248991 183138
rect 242780 183080 248930 183136
rect 248986 183080 248991 183136
rect 242780 183078 248991 183080
rect 242780 183076 242786 183078
rect 248925 183075 248991 183078
rect 137605 182594 137671 182597
rect 231445 182594 231511 182597
rect 325469 182594 325535 182597
rect 134740 182592 137671 182594
rect 134740 182536 137610 182592
rect 137666 182536 137671 182592
rect 134740 182534 137671 182536
rect 228764 182592 231511 182594
rect 228764 182536 231450 182592
rect 231506 182536 231511 182592
rect 228764 182534 231511 182536
rect 322788 182592 325535 182594
rect 322788 182536 325474 182592
rect 325530 182536 325535 182592
rect 322788 182534 325535 182536
rect 137605 182531 137671 182534
rect 231445 182531 231511 182534
rect 325469 182531 325535 182534
rect 249017 182186 249083 182189
rect 271414 182186 271420 182188
rect 249017 182184 271420 182186
rect 249017 182128 249022 182184
rect 249078 182128 271420 182184
rect 249017 182126 271420 182128
rect 249017 182123 249083 182126
rect 271414 182124 271420 182126
rect 271484 182124 271490 182188
rect 322934 182124 322940 182188
rect 323004 182186 323010 182188
rect 352885 182186 352951 182189
rect 323004 182184 352951 182186
rect 323004 182128 352890 182184
rect 352946 182128 352951 182184
rect 323004 182126 352951 182128
rect 323004 182124 323010 182126
rect 352885 182123 352951 182126
rect 154717 182050 154783 182053
rect 174814 182050 174820 182052
rect 154717 182048 174820 182050
rect 154717 181992 154722 182048
rect 154778 181992 174820 182048
rect 154717 181990 174820 181992
rect 154717 181987 154783 181990
rect 174814 181988 174820 181990
rect 174884 181988 174890 182052
rect 228910 181988 228916 182052
rect 228980 182050 228986 182052
rect 271414 182050 271420 182052
rect 228980 181990 271420 182050
rect 228980 181988 228986 181990
rect 271414 181988 271420 181990
rect 271484 181988 271490 182052
rect 322934 181988 322940 182052
rect 323004 182050 323010 182052
rect 352977 182050 353043 182053
rect 323004 182048 353043 182050
rect 323004 181992 352982 182048
rect 353038 181992 353043 182048
rect 323004 181990 353043 181992
rect 323004 181988 323010 181990
rect 352977 181987 353043 181990
rect 147030 181172 147036 181236
rect 147100 181234 147106 181236
rect 155269 181234 155335 181237
rect 147100 181232 155335 181234
rect 147100 181176 155274 181232
rect 155330 181176 155335 181232
rect 147100 181174 155335 181176
rect 147100 181172 147106 181174
rect 155269 181171 155335 181174
rect 159041 181098 159107 181101
rect 169110 181098 169116 181100
rect 159041 181096 169116 181098
rect 159041 181040 159046 181096
rect 159102 181040 169116 181096
rect 159041 181038 169116 181040
rect 159041 181035 159107 181038
rect 169110 181036 169116 181038
rect 169180 181036 169186 181100
rect 158397 180962 158463 180965
rect 168558 180962 168564 180964
rect 158397 180960 168564 180962
rect 158397 180904 158402 180960
rect 158458 180904 168564 180960
rect 158397 180902 168564 180904
rect 158397 180899 158463 180902
rect 168558 180900 168564 180902
rect 168628 180900 168634 180964
rect 157201 180826 157267 180829
rect 167638 180826 167644 180828
rect 157201 180824 167644 180826
rect 157201 180768 157206 180824
rect 157262 180768 167644 180824
rect 157201 180766 167644 180768
rect 157201 180763 157267 180766
rect 167638 180764 167644 180766
rect 167708 180764 167714 180828
rect 253341 180826 253407 180829
rect 261662 180826 261668 180828
rect 253341 180824 261668 180826
rect 253341 180768 253346 180824
rect 253402 180768 261668 180824
rect 253341 180766 261668 180768
rect 253341 180763 253407 180766
rect 261662 180764 261668 180766
rect 261732 180764 261738 180828
rect 157753 180690 157819 180693
rect 169478 180690 169484 180692
rect 157753 180688 169484 180690
rect 157753 180632 157758 180688
rect 157814 180632 169484 180688
rect 157753 180630 169484 180632
rect 157753 180627 157819 180630
rect 169478 180628 169484 180630
rect 169548 180628 169554 180692
rect 242342 180628 242348 180692
rect 242412 180690 242418 180692
rect 251409 180690 251475 180693
rect 242412 180688 251475 180690
rect 242412 180632 251414 180688
rect 251470 180632 251475 180688
rect 242412 180630 251475 180632
rect 242412 180628 242418 180630
rect 251409 180627 251475 180630
rect 252697 180690 252763 180693
rect 262398 180690 262404 180692
rect 252697 180688 262404 180690
rect 252697 180632 252702 180688
rect 252758 180632 262404 180688
rect 252697 180630 262404 180632
rect 252697 180627 252763 180630
rect 262398 180628 262404 180630
rect 262468 180628 262474 180692
rect 147950 180492 147956 180556
rect 148020 180554 148026 180556
rect 155913 180554 155979 180557
rect 148020 180552 155979 180554
rect 148020 180496 155918 180552
rect 155974 180496 155979 180552
rect 148020 180494 155979 180496
rect 148020 180492 148026 180494
rect 155913 180491 155979 180494
rect 156557 180554 156623 180557
rect 167822 180554 167828 180556
rect 156557 180552 167828 180554
rect 156557 180496 156562 180552
rect 156618 180496 167828 180552
rect 156557 180494 167828 180496
rect 156557 180491 156623 180494
rect 167822 180492 167828 180494
rect 167892 180492 167898 180556
rect 251317 180554 251383 180557
rect 262950 180554 262956 180556
rect 251317 180552 262956 180554
rect 251317 180496 251322 180552
rect 251378 180496 262956 180552
rect 251317 180494 262956 180496
rect 251317 180491 251383 180494
rect 262950 180492 262956 180494
rect 263020 180492 263026 180556
rect 241790 180084 241796 180148
rect 241860 180146 241866 180148
rect 250213 180146 250279 180149
rect 241860 180144 250279 180146
rect 241860 180088 250218 180144
rect 250274 180088 250279 180144
rect 241860 180086 250279 180088
rect 241860 180084 241866 180086
rect 250213 180083 250279 180086
rect 242894 179948 242900 180012
rect 242964 180010 242970 180012
rect 249569 180010 249635 180013
rect 242964 180008 249635 180010
rect 242964 179952 249574 180008
rect 249630 179952 249635 180008
rect 242964 179950 249635 179952
rect 242964 179948 242970 179950
rect 249569 179947 249635 179950
rect 138893 179466 138959 179469
rect 230985 179466 231051 179469
rect 324549 179466 324615 179469
rect 134740 179464 138959 179466
rect 134740 179408 138898 179464
rect 138954 179408 138959 179464
rect 134740 179406 138959 179408
rect 228764 179464 231051 179466
rect 228764 179408 230990 179464
rect 231046 179408 231051 179464
rect 228764 179406 231051 179408
rect 322788 179464 324615 179466
rect 322788 179408 324554 179464
rect 324610 179408 324615 179464
rect 322788 179406 324615 179408
rect 138893 179403 138959 179406
rect 230985 179403 231051 179406
rect 324549 179403 324615 179406
rect 287422 179268 287428 179332
rect 287492 179330 287498 179332
rect 289446 179330 289452 179332
rect 287492 179270 289452 179330
rect 287492 179268 287498 179270
rect 289446 179268 289452 179270
rect 289516 179268 289522 179332
rect 310974 179268 310980 179332
rect 311044 179330 311050 179332
rect 317046 179330 317052 179332
rect 311044 179270 317052 179330
rect 311044 179268 311050 179270
rect 317046 179268 317052 179270
rect 317116 179268 317122 179332
rect 286134 179132 286140 179196
rect 286204 179194 286210 179196
rect 288526 179194 288532 179196
rect 286204 179134 288532 179194
rect 286204 179132 286210 179134
rect 288526 179132 288532 179134
rect 288596 179132 288602 179196
rect 309870 179132 309876 179196
rect 309940 179194 309946 179196
rect 311894 179194 311900 179196
rect 309940 179134 311900 179194
rect 309940 179132 309946 179134
rect 311894 179132 311900 179134
rect 311964 179132 311970 179196
rect 178269 178244 178335 178245
rect 178269 178242 178316 178244
rect 178188 178240 178316 178242
rect 178380 178242 178386 178244
rect 182133 178242 182199 178245
rect 178380 178240 182199 178242
rect 178188 178184 178274 178240
rect 178380 178184 182138 178240
rect 182194 178184 182199 178240
rect 178188 178182 178316 178184
rect 178269 178180 178316 178182
rect 178380 178182 182199 178184
rect 178380 178180 178386 178182
rect 178269 178179 178335 178180
rect 182133 178179 182199 178182
rect 73614 177908 73620 177972
rect 73684 177970 73690 177972
rect 75454 177970 75460 177972
rect 73684 177910 75460 177970
rect 73684 177908 73690 177910
rect 75454 177908 75460 177910
rect 75524 177908 75530 177972
rect 429889 177834 429955 177837
rect 434416 177834 434896 177864
rect 429889 177832 434896 177834
rect 429889 177776 429894 177832
rect 429950 177776 434896 177832
rect 429889 177774 434896 177776
rect 429889 177771 429955 177774
rect 434416 177744 434896 177774
rect 46893 176474 46959 176477
rect 71958 176474 71964 176476
rect 46893 176472 71964 176474
rect 46893 176416 46898 176472
rect 46954 176416 71964 176472
rect 46893 176414 71964 176416
rect 46893 176411 46959 176414
rect 71958 176412 71964 176414
rect 72028 176412 72034 176476
rect 9896 176066 10376 176096
rect 13405 176066 13471 176069
rect 9896 176064 13471 176066
rect 9896 176008 13410 176064
rect 13466 176008 13471 176064
rect 9896 176006 13471 176008
rect 9896 175976 10376 176006
rect 13405 176003 13471 176006
rect 45789 175930 45855 175933
rect 46893 175930 46959 175933
rect 45789 175928 46959 175930
rect 45789 175872 45794 175928
rect 45850 175872 46898 175928
rect 46954 175872 46959 175928
rect 45789 175870 46959 175872
rect 45789 175867 45855 175870
rect 46893 175867 46959 175870
rect 71958 175868 71964 175932
rect 72028 175930 72034 175932
rect 72326 175930 72332 175932
rect 72028 175870 72332 175930
rect 72028 175868 72034 175870
rect 72326 175868 72332 175870
rect 72396 175868 72402 175932
rect 182869 175796 182935 175797
rect 182869 175792 182916 175796
rect 182980 175794 182986 175796
rect 182869 175736 182874 175792
rect 182869 175732 182916 175736
rect 182980 175734 183026 175794
rect 182980 175732 182986 175734
rect 182869 175731 182935 175732
rect 218013 175522 218079 175525
rect 219710 175522 219716 175524
rect 218013 175520 219716 175522
rect 218013 175464 218018 175520
rect 218074 175464 219716 175520
rect 218013 175462 219716 175464
rect 218013 175459 218079 175462
rect 219710 175460 219716 175462
rect 219780 175460 219786 175524
rect 74166 173692 74172 173756
rect 74236 173754 74242 173756
rect 74309 173754 74375 173757
rect 74236 173752 74375 173754
rect 74236 173696 74314 173752
rect 74370 173696 74375 173752
rect 74236 173694 74375 173696
rect 74236 173692 74242 173694
rect 74309 173691 74375 173694
rect 368525 173074 368591 173077
rect 368709 173074 368775 173077
rect 368525 173072 368775 173074
rect 368525 173016 368530 173072
rect 368586 173016 368714 173072
rect 368770 173016 368775 173072
rect 368525 173014 368775 173016
rect 368525 173011 368591 173014
rect 368709 173011 368775 173014
rect 52638 172876 52644 172940
rect 52708 172938 52714 172940
rect 53517 172938 53583 172941
rect 52708 172936 53583 172938
rect 52708 172880 53522 172936
rect 53578 172880 53583 172936
rect 52708 172878 53583 172880
rect 52708 172876 52714 172878
rect 53517 172875 53583 172878
rect 54529 172938 54595 172941
rect 55541 172940 55607 172941
rect 54662 172938 54668 172940
rect 54529 172936 54668 172938
rect 54529 172880 54534 172936
rect 54590 172880 54668 172936
rect 54529 172878 54668 172880
rect 54529 172875 54595 172878
rect 54662 172876 54668 172878
rect 54732 172876 54738 172940
rect 55541 172938 55588 172940
rect 55496 172936 55588 172938
rect 55496 172880 55546 172936
rect 55496 172878 55588 172880
rect 55541 172876 55588 172878
rect 55652 172876 55658 172940
rect 55541 172875 55607 172876
rect 55398 172740 55404 172804
rect 55468 172802 55474 172804
rect 56553 172802 56619 172805
rect 55468 172800 56619 172802
rect 55468 172744 56558 172800
rect 56614 172744 56619 172800
rect 55468 172742 56619 172744
rect 55468 172740 55474 172742
rect 56553 172739 56619 172742
rect 350953 172666 351019 172669
rect 351638 172666 351644 172668
rect 350953 172664 351644 172666
rect 350953 172608 350958 172664
rect 351014 172608 351644 172664
rect 350953 172606 351644 172608
rect 350953 172603 351019 172606
rect 351638 172604 351644 172606
rect 351708 172604 351714 172668
rect 351822 172604 351828 172668
rect 351892 172666 351898 172668
rect 352057 172666 352123 172669
rect 351892 172664 352123 172666
rect 351892 172608 352062 172664
rect 352118 172608 352123 172664
rect 351892 172606 352123 172608
rect 351892 172604 351898 172606
rect 352057 172603 352123 172606
rect 75454 169748 75460 169812
rect 75524 169810 75530 169812
rect 76742 169810 76748 169812
rect 75524 169750 76748 169810
rect 75524 169748 75530 169750
rect 76742 169748 76748 169750
rect 76812 169748 76818 169812
rect 74166 169612 74172 169676
rect 74236 169674 74242 169676
rect 76374 169674 76380 169676
rect 74236 169614 76380 169674
rect 74236 169612 74242 169614
rect 76374 169612 76380 169614
rect 76444 169612 76450 169676
rect 71641 169538 71707 169541
rect 73430 169538 73436 169540
rect 71641 169536 73436 169538
rect 71641 169480 71646 169536
rect 71702 169480 73436 169536
rect 71641 169478 73436 169480
rect 71641 169475 71707 169478
rect 73430 169476 73436 169478
rect 73500 169476 73506 169540
rect 73798 169476 73804 169540
rect 73868 169538 73874 169540
rect 75454 169538 75460 169540
rect 73868 169478 75460 169538
rect 73868 169476 73874 169478
rect 75454 169476 75460 169478
rect 75524 169476 75530 169540
rect 74718 169340 74724 169404
rect 74788 169402 74794 169404
rect 75638 169402 75644 169404
rect 74788 169342 75644 169402
rect 74788 169340 74794 169342
rect 75638 169340 75644 169342
rect 75708 169340 75714 169404
rect 72326 169204 72332 169268
rect 72396 169266 72402 169268
rect 75822 169266 75828 169268
rect 72396 169206 75828 169266
rect 72396 169204 72402 169206
rect 75822 169204 75828 169206
rect 75892 169204 75898 169268
rect 144086 169204 144092 169268
rect 144156 169266 144162 169268
rect 147950 169266 147956 169268
rect 144156 169206 147956 169266
rect 144156 169204 144162 169206
rect 147950 169204 147956 169206
rect 148020 169204 148026 169268
rect 79737 169130 79803 169133
rect 76780 169128 79803 169130
rect 76780 169072 79742 169128
rect 79798 169072 79803 169128
rect 76780 169070 79803 169072
rect 79737 169067 79803 169070
rect 140549 169130 140615 169133
rect 173577 169130 173643 169133
rect 140549 169128 143020 169130
rect 140549 169072 140554 169128
rect 140610 169072 143020 169128
rect 140549 169070 143020 169072
rect 170804 169128 173643 169130
rect 170804 169072 173582 169128
rect 173638 169072 173643 169128
rect 170804 169070 173643 169072
rect 140549 169067 140615 169070
rect 173577 169067 173643 169070
rect 233469 169130 233535 169133
rect 267417 169130 267483 169133
rect 233469 169128 237044 169130
rect 233469 169072 233474 169128
rect 233530 169072 237044 169128
rect 233469 169070 237044 169072
rect 264828 169128 267483 169130
rect 264828 169072 267422 169128
rect 267478 169072 267483 169128
rect 264828 169070 267483 169072
rect 233469 169067 233535 169070
rect 267417 169067 267483 169070
rect 328413 169130 328479 169133
rect 328413 169128 331068 169130
rect 328413 169072 328418 169128
rect 328474 169072 331068 169128
rect 328413 169070 331068 169072
rect 328413 169067 328479 169070
rect 49193 168858 49259 168861
rect 49150 168856 49259 168858
rect 49150 168800 49198 168856
rect 49254 168800 49259 168856
rect 49150 168795 49259 168800
rect 49150 168284 49210 168795
rect 359049 168314 359115 168317
rect 359693 168314 359759 168317
rect 358852 168312 359759 168314
rect 358852 168256 359054 168312
rect 359110 168256 359698 168312
rect 359754 168256 359759 168312
rect 358852 168254 359759 168256
rect 359049 168251 359115 168254
rect 359693 168251 359759 168254
rect 140549 167770 140615 167773
rect 173393 167770 173459 167773
rect 140549 167768 143020 167770
rect 140549 167712 140554 167768
rect 140610 167712 143020 167768
rect 140549 167710 143020 167712
rect 170804 167768 173459 167770
rect 170804 167712 173398 167768
rect 173454 167712 173459 167768
rect 170804 167710 173459 167712
rect 140549 167707 140615 167710
rect 173393 167707 173459 167710
rect 233469 167770 233535 167773
rect 267693 167770 267759 167773
rect 233469 167768 237044 167770
rect 233469 167712 233474 167768
rect 233530 167712 237044 167768
rect 233469 167710 237044 167712
rect 264828 167768 267759 167770
rect 264828 167712 267698 167768
rect 267754 167712 267759 167768
rect 264828 167710 267759 167712
rect 233469 167707 233535 167710
rect 267693 167707 267759 167710
rect 327217 167770 327283 167773
rect 327217 167768 331068 167770
rect 327217 167712 327222 167768
rect 327278 167712 331068 167768
rect 327217 167710 331068 167712
rect 327217 167707 327283 167710
rect 77253 167702 77319 167705
rect 76780 167700 77319 167702
rect 76780 167644 77258 167700
rect 77314 167644 77319 167700
rect 76780 167642 77319 167644
rect 77253 167639 77319 167642
rect 236873 167090 236939 167093
rect 237006 167090 237012 167092
rect 236873 167088 237012 167090
rect 236873 167032 236878 167088
rect 236934 167032 237012 167088
rect 236873 167030 237012 167032
rect 236873 167027 236939 167030
rect 237006 167028 237012 167030
rect 237076 167028 237082 167092
rect 140549 166410 140615 166413
rect 173485 166410 173551 166413
rect 140549 166408 143020 166410
rect 140549 166352 140554 166408
rect 140610 166352 143020 166408
rect 140549 166350 143020 166352
rect 170804 166408 173551 166410
rect 170804 166352 173490 166408
rect 173546 166352 173551 166408
rect 170804 166350 173551 166352
rect 140549 166347 140615 166350
rect 173485 166347 173551 166350
rect 233469 166410 233535 166413
rect 267509 166410 267575 166413
rect 233469 166408 237044 166410
rect 233469 166352 233474 166408
rect 233530 166352 237044 166408
rect 233469 166350 237044 166352
rect 264828 166408 267575 166410
rect 264828 166352 267514 166408
rect 267570 166352 267575 166408
rect 264828 166350 267575 166352
rect 233469 166347 233535 166350
rect 267509 166347 267575 166350
rect 328413 166410 328479 166413
rect 328413 166408 331068 166410
rect 328413 166352 328418 166408
rect 328474 166352 331068 166408
rect 328413 166350 331068 166352
rect 328413 166347 328479 166350
rect 77253 166342 77319 166345
rect 76780 166340 77319 166342
rect 76780 166284 77258 166340
rect 77314 166284 77319 166340
rect 76780 166282 77319 166284
rect 77253 166279 77319 166282
rect 428785 165322 428851 165325
rect 434416 165322 434896 165352
rect 428785 165320 434896 165322
rect 428785 165264 428790 165320
rect 428846 165264 434896 165320
rect 428785 165262 434896 165264
rect 428785 165259 428851 165262
rect 434416 165232 434896 165262
rect 46893 165186 46959 165189
rect 360429 165186 360495 165189
rect 361257 165186 361323 165189
rect 46893 165184 48996 165186
rect 46893 165128 46898 165184
rect 46954 165128 48996 165184
rect 46893 165126 48996 165128
rect 358852 165184 361323 165186
rect 358852 165128 360434 165184
rect 360490 165128 361262 165184
rect 361318 165128 361323 165184
rect 358852 165126 361323 165128
rect 46893 165123 46959 165126
rect 360429 165123 360495 165126
rect 361257 165123 361323 165126
rect 79737 164914 79803 164917
rect 76780 164912 79803 164914
rect 76780 164856 79742 164912
rect 79798 164856 79803 164912
rect 76780 164854 79803 164856
rect 79737 164851 79803 164854
rect 139629 164914 139695 164917
rect 173301 164914 173367 164917
rect 139629 164912 143020 164914
rect 139629 164856 139634 164912
rect 139690 164856 143020 164912
rect 139629 164854 143020 164856
rect 170804 164912 173367 164914
rect 170804 164856 173306 164912
rect 173362 164856 173367 164912
rect 170804 164854 173367 164856
rect 139629 164851 139695 164854
rect 173301 164851 173367 164854
rect 233469 164914 233535 164917
rect 267141 164914 267207 164917
rect 233469 164912 237044 164914
rect 233469 164856 233474 164912
rect 233530 164856 237044 164912
rect 233469 164854 237044 164856
rect 264828 164912 267207 164914
rect 264828 164856 267146 164912
rect 267202 164856 267207 164912
rect 264828 164854 267207 164856
rect 233469 164851 233535 164854
rect 267141 164851 267207 164854
rect 328505 164914 328571 164917
rect 328505 164912 331068 164914
rect 328505 164856 328510 164912
rect 328566 164856 331068 164912
rect 328505 164854 331068 164856
rect 328505 164851 328571 164854
rect 87189 164098 87255 164101
rect 87189 164096 90058 164098
rect 87189 164040 87194 164096
rect 87250 164040 90058 164096
rect 87189 164038 90058 164040
rect 87189 164035 87255 164038
rect 77253 163486 77319 163489
rect 76780 163484 77319 163486
rect 76780 163428 77258 163484
rect 77314 163428 77319 163484
rect 89998 163456 90058 164038
rect 139629 163554 139695 163557
rect 174037 163554 174103 163557
rect 139629 163552 143020 163554
rect 139629 163496 139634 163552
rect 139690 163496 143020 163552
rect 139629 163494 143020 163496
rect 170804 163552 174103 163554
rect 170804 163496 174042 163552
rect 174098 163496 174103 163552
rect 170804 163494 174103 163496
rect 139629 163491 139695 163494
rect 174037 163491 174103 163494
rect 233469 163554 233535 163557
rect 267877 163554 267943 163557
rect 233469 163552 237044 163554
rect 233469 163496 233474 163552
rect 233530 163496 237044 163552
rect 233469 163494 237044 163496
rect 264828 163552 267943 163554
rect 264828 163496 267882 163552
rect 267938 163496 267943 163552
rect 264828 163494 267943 163496
rect 233469 163491 233535 163494
rect 267877 163491 267943 163494
rect 76780 163426 77319 163428
rect 77253 163423 77319 163426
rect 330486 163426 331068 163486
rect 131349 163418 131415 163421
rect 129772 163416 131415 163418
rect 129772 163360 131354 163416
rect 131410 163360 131415 163416
rect 129772 163358 131415 163360
rect 131349 163355 131415 163358
rect 182317 163418 182383 163421
rect 226293 163418 226359 163421
rect 182317 163416 184052 163418
rect 182317 163360 182322 163416
rect 182378 163360 184052 163416
rect 182317 163358 184052 163360
rect 223796 163416 226359 163418
rect 223796 163360 226298 163416
rect 226354 163360 226359 163416
rect 223796 163358 226359 163360
rect 182317 163355 182383 163358
rect 226293 163355 226359 163358
rect 274501 163418 274567 163421
rect 321605 163418 321671 163421
rect 274501 163416 278076 163418
rect 274501 163360 274506 163416
rect 274562 163360 278076 163416
rect 274501 163358 278076 163360
rect 317820 163416 321671 163418
rect 317820 163360 321610 163416
rect 321666 163360 321671 163416
rect 317820 163358 321671 163360
rect 274501 163355 274567 163358
rect 321605 163355 321671 163358
rect 327217 163418 327283 163421
rect 330486 163418 330546 163426
rect 327217 163416 330546 163418
rect 327217 163360 327222 163416
rect 327278 163360 330546 163416
rect 327217 163358 330546 163360
rect 327217 163355 327283 163358
rect 87189 163146 87255 163149
rect 87189 163144 90058 163146
rect 87189 163088 87194 163144
rect 87250 163088 90058 163144
rect 87189 163086 90058 163088
rect 87189 163083 87255 163086
rect 9896 162738 10376 162768
rect 12853 162738 12919 162741
rect 9896 162736 12919 162738
rect 9896 162680 12858 162736
rect 12914 162680 12919 162736
rect 9896 162678 12919 162680
rect 9896 162648 10376 162678
rect 12853 162675 12919 162678
rect 48958 162540 48964 162604
rect 49028 162540 49034 162604
rect 46617 162058 46683 162061
rect 48966 162058 49026 162540
rect 89998 162504 90058 163086
rect 131993 162466 132059 162469
rect 129772 162464 132059 162466
rect 129772 162408 131998 162464
rect 132054 162408 132059 162464
rect 129772 162406 132059 162408
rect 131993 162403 132059 162406
rect 181765 162466 181831 162469
rect 226293 162466 226359 162469
rect 181765 162464 184052 162466
rect 181765 162408 181770 162464
rect 181826 162408 184052 162464
rect 181765 162406 184052 162408
rect 223796 162464 226359 162466
rect 223796 162408 226298 162464
rect 226354 162408 226359 162464
rect 223796 162406 226359 162408
rect 181765 162403 181831 162406
rect 226293 162403 226359 162406
rect 274869 162466 274935 162469
rect 320961 162466 321027 162469
rect 274869 162464 278076 162466
rect 274869 162408 274874 162464
rect 274930 162408 278076 162464
rect 274869 162406 278076 162408
rect 317820 162464 321027 162466
rect 317820 162408 320966 162464
rect 321022 162408 321027 162464
rect 317820 162406 321027 162408
rect 274869 162403 274935 162406
rect 320961 162403 321027 162406
rect 139629 162194 139695 162197
rect 173669 162194 173735 162197
rect 139629 162192 143020 162194
rect 139629 162136 139634 162192
rect 139690 162136 143020 162192
rect 139629 162134 143020 162136
rect 170804 162192 173735 162194
rect 170804 162136 173674 162192
rect 173730 162136 173735 162192
rect 170804 162134 173735 162136
rect 139629 162131 139695 162134
rect 173669 162131 173735 162134
rect 233469 162194 233535 162197
rect 267049 162194 267115 162197
rect 233469 162192 237044 162194
rect 233469 162136 233474 162192
rect 233530 162136 237044 162192
rect 233469 162134 237044 162136
rect 264828 162192 267115 162194
rect 264828 162136 267054 162192
rect 267110 162136 267115 162192
rect 264828 162134 267115 162136
rect 233469 162131 233535 162134
rect 267049 162131 267115 162134
rect 328413 162194 328479 162197
rect 328413 162192 331068 162194
rect 328413 162136 328418 162192
rect 328474 162136 331068 162192
rect 328413 162134 331068 162136
rect 328413 162131 328479 162134
rect 77161 162126 77227 162129
rect 76780 162124 77227 162126
rect 76780 162068 77166 162124
rect 77222 162068 77227 162124
rect 76780 162066 77227 162068
rect 77161 162063 77227 162066
rect 360521 162058 360587 162061
rect 46617 162056 49026 162058
rect 46617 162000 46622 162056
rect 46678 162028 49026 162056
rect 358852 162056 360587 162058
rect 46678 162000 48996 162028
rect 46617 161998 48996 162000
rect 358852 162000 360526 162056
rect 360582 162000 360587 162056
rect 358852 161998 360587 162000
rect 46617 161995 46683 161998
rect 360521 161995 360587 161998
rect 87281 161922 87347 161925
rect 321789 161922 321855 161925
rect 87281 161920 90058 161922
rect 87281 161864 87286 161920
rect 87342 161864 90058 161920
rect 87281 161862 90058 161864
rect 87281 161859 87347 161862
rect 89998 161688 90058 161862
rect 317790 161920 321855 161922
rect 317790 161864 321794 161920
rect 321850 161864 321855 161920
rect 317790 161862 321855 161864
rect 131533 161650 131599 161653
rect 129772 161648 131599 161650
rect 129772 161592 131538 161648
rect 131594 161592 131599 161648
rect 129772 161590 131599 161592
rect 131533 161587 131599 161590
rect 182317 161650 182383 161653
rect 226385 161650 226451 161653
rect 182317 161648 184052 161650
rect 182317 161592 182322 161648
rect 182378 161592 184052 161648
rect 182317 161590 184052 161592
rect 223796 161648 226451 161650
rect 223796 161592 226390 161648
rect 226446 161592 226451 161648
rect 223796 161590 226451 161592
rect 182317 161587 182383 161590
rect 226385 161587 226451 161590
rect 274869 161650 274935 161653
rect 274869 161648 278076 161650
rect 274869 161592 274874 161648
rect 274930 161592 278076 161648
rect 317790 161620 317850 161862
rect 321789 161859 321855 161862
rect 274869 161590 278076 161592
rect 274869 161587 274935 161590
rect 87189 161378 87255 161381
rect 87189 161376 90058 161378
rect 87189 161320 87194 161376
rect 87250 161320 90058 161376
rect 87189 161318 90058 161320
rect 87189 161315 87255 161318
rect 89998 160736 90058 161318
rect 131349 160698 131415 160701
rect 129772 160696 131415 160698
rect 129772 160640 131354 160696
rect 131410 160640 131415 160696
rect 129772 160638 131415 160640
rect 131349 160635 131415 160638
rect 139629 160698 139695 160701
rect 173945 160698 174011 160701
rect 139629 160696 143020 160698
rect 139629 160640 139634 160696
rect 139690 160640 143020 160696
rect 139629 160638 143020 160640
rect 170804 160696 174011 160698
rect 170804 160640 173950 160696
rect 174006 160640 174011 160696
rect 170804 160638 174011 160640
rect 139629 160635 139695 160638
rect 173945 160635 174011 160638
rect 181673 160698 181739 160701
rect 225649 160698 225715 160701
rect 181673 160696 184052 160698
rect 181673 160640 181678 160696
rect 181734 160640 184052 160696
rect 181673 160638 184052 160640
rect 223796 160696 225715 160698
rect 223796 160640 225654 160696
rect 225710 160640 225715 160696
rect 223796 160638 225715 160640
rect 181673 160635 181739 160638
rect 225649 160635 225715 160638
rect 233469 160698 233535 160701
rect 266589 160698 266655 160701
rect 233469 160696 237044 160698
rect 233469 160640 233474 160696
rect 233530 160640 237044 160696
rect 233469 160638 237044 160640
rect 264828 160696 266655 160698
rect 264828 160640 266594 160696
rect 266650 160640 266655 160696
rect 264828 160638 266655 160640
rect 233469 160635 233535 160638
rect 266589 160635 266655 160638
rect 274869 160698 274935 160701
rect 320777 160698 320843 160701
rect 274869 160696 278076 160698
rect 274869 160640 274874 160696
rect 274930 160640 278076 160696
rect 274869 160638 278076 160640
rect 317820 160696 320843 160698
rect 317820 160640 320782 160696
rect 320838 160640 320843 160696
rect 317820 160638 320843 160640
rect 274869 160635 274935 160638
rect 320777 160635 320843 160638
rect 327309 160698 327375 160701
rect 327309 160696 331068 160698
rect 327309 160640 327314 160696
rect 327370 160640 331068 160696
rect 327309 160638 331068 160640
rect 327309 160635 327375 160638
rect 76750 160018 76810 160600
rect 87189 160426 87255 160429
rect 87189 160424 90058 160426
rect 87189 160368 87194 160424
rect 87250 160368 90058 160424
rect 87189 160366 90058 160368
rect 87189 160363 87255 160366
rect 81669 160018 81735 160021
rect 76750 160016 81735 160018
rect 76750 159960 81674 160016
rect 81730 159960 81735 160016
rect 76750 159958 81735 159960
rect 81669 159955 81735 159958
rect 89998 159920 90058 160366
rect 131809 159882 131875 159885
rect 129772 159880 131875 159882
rect 129772 159824 131814 159880
rect 131870 159824 131875 159880
rect 129772 159822 131875 159824
rect 131809 159819 131875 159822
rect 182317 159882 182383 159885
rect 226293 159882 226359 159885
rect 182317 159880 184052 159882
rect 182317 159824 182322 159880
rect 182378 159824 184052 159880
rect 182317 159822 184052 159824
rect 223796 159880 226359 159882
rect 223796 159824 226298 159880
rect 226354 159824 226359 159880
rect 223796 159822 226359 159824
rect 182317 159819 182383 159822
rect 226293 159819 226359 159822
rect 275697 159882 275763 159885
rect 321697 159882 321763 159885
rect 275697 159880 278076 159882
rect 275697 159824 275702 159880
rect 275758 159824 278076 159880
rect 275697 159822 278076 159824
rect 317820 159880 321763 159882
rect 317820 159824 321702 159880
rect 321758 159824 321763 159880
rect 317820 159822 321763 159824
rect 275697 159819 275763 159822
rect 321697 159819 321763 159822
rect 79277 159338 79343 159341
rect 76780 159336 79343 159338
rect 76780 159280 79282 159336
rect 79338 159280 79343 159336
rect 76780 159278 79343 159280
rect 79277 159275 79343 159278
rect 139629 159338 139695 159341
rect 173945 159338 174011 159341
rect 139629 159336 143020 159338
rect 139629 159280 139634 159336
rect 139690 159280 143020 159336
rect 139629 159278 143020 159280
rect 170804 159336 174011 159338
rect 170804 159280 173950 159336
rect 174006 159280 174011 159336
rect 170804 159278 174011 159280
rect 139629 159275 139695 159278
rect 173945 159275 174011 159278
rect 233469 159338 233535 159341
rect 266589 159338 266655 159341
rect 233469 159336 237044 159338
rect 233469 159280 233474 159336
rect 233530 159280 237044 159336
rect 233469 159278 237044 159280
rect 264828 159336 266655 159338
rect 264828 159280 266594 159336
rect 266650 159280 266655 159336
rect 264828 159278 266655 159280
rect 233469 159275 233535 159278
rect 266589 159275 266655 159278
rect 327217 159338 327283 159341
rect 327217 159336 331068 159338
rect 327217 159280 327222 159336
rect 327278 159280 331068 159336
rect 327217 159278 331068 159280
rect 327217 159275 327283 159278
rect 46525 158930 46591 158933
rect 87189 158930 87255 158933
rect 131349 158930 131415 158933
rect 226385 158930 226451 158933
rect 46525 158928 49180 158930
rect 46525 158872 46530 158928
rect 46586 158900 49180 158928
rect 87189 158928 90028 158930
rect 46586 158872 49210 158900
rect 46525 158870 49210 158872
rect 46525 158867 46591 158870
rect 49150 158388 49210 158870
rect 87189 158872 87194 158928
rect 87250 158872 90028 158928
rect 87189 158870 90028 158872
rect 129772 158928 131415 158930
rect 129772 158872 131354 158928
rect 131410 158872 131415 158928
rect 223796 158928 226451 158930
rect 129772 158870 131415 158872
rect 87189 158867 87255 158870
rect 131349 158867 131415 158870
rect 87281 158658 87347 158661
rect 87281 158656 90058 158658
rect 87281 158600 87286 158656
rect 87342 158600 90058 158656
rect 87281 158598 90058 158600
rect 87281 158595 87347 158598
rect 49142 158324 49148 158388
rect 49212 158324 49218 158388
rect 89998 158152 90058 158598
rect 180293 158386 180359 158389
rect 184022 158386 184082 158900
rect 223796 158872 226390 158928
rect 226446 158872 226451 158928
rect 223796 158870 226451 158872
rect 226385 158867 226451 158870
rect 274133 158930 274199 158933
rect 321053 158930 321119 158933
rect 360613 158930 360679 158933
rect 361257 158930 361323 158933
rect 274133 158928 278076 158930
rect 274133 158872 274138 158928
rect 274194 158872 278076 158928
rect 274133 158870 278076 158872
rect 317820 158928 321119 158930
rect 317820 158872 321058 158928
rect 321114 158872 321119 158928
rect 317820 158870 321119 158872
rect 358852 158928 361323 158930
rect 358852 158872 360618 158928
rect 360674 158872 361262 158928
rect 361318 158872 361323 158928
rect 358852 158870 361323 158872
rect 274133 158867 274199 158870
rect 321053 158867 321119 158870
rect 360613 158867 360679 158870
rect 361257 158867 361323 158870
rect 180293 158384 184082 158386
rect 180293 158328 180298 158384
rect 180354 158328 184082 158384
rect 180293 158326 184082 158328
rect 180293 158323 180359 158326
rect 132269 158114 132335 158117
rect 129772 158112 132335 158114
rect 129772 158056 132274 158112
rect 132330 158056 132335 158112
rect 129772 158054 132335 158056
rect 132269 158051 132335 158054
rect 182317 158114 182383 158117
rect 226293 158114 226359 158117
rect 182317 158112 184052 158114
rect 182317 158056 182322 158112
rect 182378 158056 184052 158112
rect 182317 158054 184052 158056
rect 223796 158112 226359 158114
rect 223796 158056 226298 158112
rect 226354 158056 226359 158112
rect 223796 158054 226359 158056
rect 182317 158051 182383 158054
rect 226293 158051 226359 158054
rect 275513 158114 275579 158117
rect 321605 158114 321671 158117
rect 275513 158112 278076 158114
rect 275513 158056 275518 158112
rect 275574 158056 278076 158112
rect 275513 158054 278076 158056
rect 317820 158112 321671 158114
rect 317820 158056 321610 158112
rect 321666 158056 321671 158112
rect 317820 158054 321671 158056
rect 275513 158051 275579 158054
rect 321605 158051 321671 158054
rect 79737 157978 79803 157981
rect 76780 157976 79803 157978
rect 76780 157920 79742 157976
rect 79798 157920 79803 157976
rect 76780 157918 79803 157920
rect 79737 157915 79803 157918
rect 139629 157978 139695 157981
rect 173761 157978 173827 157981
rect 139629 157976 143020 157978
rect 139629 157920 139634 157976
rect 139690 157920 143020 157976
rect 139629 157918 143020 157920
rect 170804 157976 173827 157978
rect 170804 157920 173766 157976
rect 173822 157920 173827 157976
rect 170804 157918 173827 157920
rect 139629 157915 139695 157918
rect 173761 157915 173827 157918
rect 233469 157978 233535 157981
rect 266589 157978 266655 157981
rect 233469 157976 237044 157978
rect 233469 157920 233474 157976
rect 233530 157920 237044 157976
rect 233469 157918 237044 157920
rect 264828 157976 266655 157978
rect 264828 157920 266594 157976
rect 266650 157920 266655 157976
rect 264828 157918 266655 157920
rect 233469 157915 233535 157918
rect 266589 157915 266655 157918
rect 327217 157978 327283 157981
rect 327217 157976 331068 157978
rect 327217 157920 327222 157976
rect 327278 157920 331068 157976
rect 327217 157918 331068 157920
rect 327217 157915 327283 157918
rect 87189 157842 87255 157845
rect 87189 157840 90058 157842
rect 87189 157784 87194 157840
rect 87250 157784 90058 157840
rect 87189 157782 90058 157784
rect 87189 157779 87255 157782
rect 76558 157508 76564 157572
rect 76628 157508 76634 157572
rect 76566 157162 76626 157508
rect 89998 157200 90058 157782
rect 76742 157162 76748 157164
rect 76566 157102 76748 157162
rect 76742 157100 76748 157102
rect 76812 157100 76818 157164
rect 132453 157162 132519 157165
rect 129772 157160 132519 157162
rect 129772 157104 132458 157160
rect 132514 157104 132519 157160
rect 129772 157102 132519 157104
rect 132453 157099 132519 157102
rect 181765 157162 181831 157165
rect 226385 157162 226451 157165
rect 181765 157160 184052 157162
rect 181765 157104 181770 157160
rect 181826 157104 184052 157160
rect 181765 157102 184052 157104
rect 223796 157160 226451 157162
rect 223796 157104 226390 157160
rect 226446 157104 226451 157160
rect 223796 157102 226451 157104
rect 181765 157099 181831 157102
rect 226385 157099 226451 157102
rect 275605 157162 275671 157165
rect 321605 157162 321671 157165
rect 275605 157160 278076 157162
rect 275605 157104 275610 157160
rect 275666 157104 278076 157160
rect 275605 157102 278076 157104
rect 317820 157160 321671 157162
rect 317820 157104 321610 157160
rect 321666 157104 321671 157160
rect 317820 157102 321671 157104
rect 275605 157099 275671 157102
rect 321605 157099 321671 157102
rect 140365 156618 140431 156621
rect 172841 156618 172907 156621
rect 140365 156616 143020 156618
rect 140365 156560 140370 156616
rect 140426 156560 143020 156616
rect 140365 156558 143020 156560
rect 170804 156616 172907 156618
rect 170804 156560 172846 156616
rect 172902 156560 172907 156616
rect 170804 156558 172907 156560
rect 140365 156555 140431 156558
rect 172841 156555 172907 156558
rect 233469 156618 233535 156621
rect 267325 156618 267391 156621
rect 233469 156616 237044 156618
rect 233469 156560 233474 156616
rect 233530 156560 237044 156616
rect 233469 156558 237044 156560
rect 264828 156616 267391 156618
rect 264828 156560 267330 156616
rect 267386 156560 267391 156616
rect 264828 156558 267391 156560
rect 233469 156555 233535 156558
rect 267325 156555 267391 156558
rect 327217 156618 327283 156621
rect 327217 156616 331068 156618
rect 327217 156560 327222 156616
rect 327278 156560 331068 156616
rect 327217 156558 331068 156560
rect 327217 156555 327283 156558
rect 77253 156550 77319 156553
rect 76780 156548 77319 156550
rect 76780 156492 77258 156548
rect 77314 156492 77319 156548
rect 76780 156490 77319 156492
rect 77253 156487 77319 156490
rect 87189 156346 87255 156349
rect 132361 156346 132427 156349
rect 87189 156344 90028 156346
rect 87189 156288 87194 156344
rect 87250 156288 90028 156344
rect 87189 156286 90028 156288
rect 129772 156344 132427 156346
rect 129772 156288 132366 156344
rect 132422 156288 132427 156344
rect 129772 156286 132427 156288
rect 87189 156283 87255 156286
rect 132361 156283 132427 156286
rect 182225 156346 182291 156349
rect 226477 156346 226543 156349
rect 182225 156344 184052 156346
rect 182225 156288 182230 156344
rect 182286 156288 184052 156344
rect 182225 156286 184052 156288
rect 223796 156344 226543 156346
rect 223796 156288 226482 156344
rect 226538 156288 226543 156344
rect 223796 156286 226543 156288
rect 182225 156283 182291 156286
rect 226477 156283 226543 156286
rect 274961 156346 275027 156349
rect 321605 156346 321671 156349
rect 274961 156344 278076 156346
rect 274961 156288 274966 156344
rect 275022 156288 278076 156344
rect 274961 156286 278076 156288
rect 317820 156344 321671 156346
rect 317820 156288 321610 156344
rect 321666 156288 321671 156344
rect 317820 156286 321671 156288
rect 274961 156283 275027 156286
rect 321605 156283 321671 156286
rect 132177 156074 132243 156077
rect 129742 156072 132243 156074
rect 129742 156016 132182 156072
rect 132238 156016 132243 156072
rect 129742 156014 132243 156016
rect 46433 155802 46499 155805
rect 46433 155800 49180 155802
rect 46433 155744 46438 155800
rect 46494 155772 49180 155800
rect 46494 155744 49210 155772
rect 46433 155742 49210 155744
rect 46433 155739 46499 155742
rect 49150 155396 49210 155742
rect 129742 155432 129802 156014
rect 132177 156011 132243 156014
rect 182317 156074 182383 156077
rect 274869 156074 274935 156077
rect 182317 156072 184082 156074
rect 182317 156016 182322 156072
rect 182378 156016 184082 156072
rect 182317 156014 184082 156016
rect 182317 156011 182383 156014
rect 184022 155432 184082 156014
rect 274869 156072 278106 156074
rect 274869 156016 274874 156072
rect 274930 156016 278106 156072
rect 274869 156014 278106 156016
rect 274869 156011 274935 156014
rect 278046 155432 278106 156014
rect 360705 155802 360771 155805
rect 361165 155802 361231 155805
rect 358852 155800 361231 155802
rect 358852 155744 360710 155800
rect 360766 155744 361170 155800
rect 361226 155744 361231 155800
rect 358852 155742 361231 155744
rect 360705 155739 360771 155742
rect 361165 155739 361231 155742
rect 49142 155332 49148 155396
rect 49212 155332 49218 155396
rect 87189 155394 87255 155397
rect 225833 155394 225899 155397
rect 321605 155394 321671 155397
rect 87189 155392 90028 155394
rect 87189 155336 87194 155392
rect 87250 155336 90028 155392
rect 87189 155334 90028 155336
rect 223796 155392 225899 155394
rect 223796 155336 225838 155392
rect 225894 155336 225899 155392
rect 223796 155334 225899 155336
rect 317820 155392 321671 155394
rect 317820 155336 321610 155392
rect 321666 155336 321671 155392
rect 317820 155334 321671 155336
rect 87189 155331 87255 155334
rect 225833 155331 225899 155334
rect 321605 155331 321671 155334
rect 79737 155122 79803 155125
rect 131993 155122 132059 155125
rect 76780 155120 79803 155122
rect 76780 155064 79742 155120
rect 79798 155064 79803 155120
rect 76780 155062 79803 155064
rect 79737 155059 79803 155062
rect 129742 155120 132059 155122
rect 129742 155064 131998 155120
rect 132054 155064 132059 155120
rect 129742 155062 132059 155064
rect 129742 154480 129802 155062
rect 131993 155059 132059 155062
rect 140549 155122 140615 155125
rect 174037 155122 174103 155125
rect 140549 155120 143020 155122
rect 140549 155064 140554 155120
rect 140610 155064 143020 155120
rect 140549 155062 143020 155064
rect 170804 155120 174103 155122
rect 170804 155064 174042 155120
rect 174098 155064 174103 155120
rect 170804 155062 174103 155064
rect 140549 155059 140615 155062
rect 174037 155059 174103 155062
rect 232825 155122 232891 155125
rect 266589 155122 266655 155125
rect 232825 155120 237044 155122
rect 232825 155064 232830 155120
rect 232886 155064 237044 155120
rect 232825 155062 237044 155064
rect 264828 155120 266655 155122
rect 264828 155064 266594 155120
rect 266650 155064 266655 155120
rect 264828 155062 266655 155064
rect 232825 155059 232891 155062
rect 266589 155059 266655 155062
rect 328413 155122 328479 155125
rect 328413 155120 331068 155122
rect 328413 155064 328418 155120
rect 328474 155064 331068 155120
rect 328413 155062 331068 155064
rect 328413 155059 328479 155062
rect 274869 154986 274935 154989
rect 274869 154984 278106 154986
rect 274869 154928 274874 154984
rect 274930 154928 278106 154984
rect 274869 154926 278106 154928
rect 274869 154923 274935 154926
rect 181121 154714 181187 154717
rect 181121 154712 184082 154714
rect 181121 154656 181126 154712
rect 181182 154656 184082 154712
rect 181121 154654 184082 154656
rect 181121 154651 181187 154654
rect 184022 154480 184082 154654
rect 278046 154480 278106 154926
rect 87189 154442 87255 154445
rect 226017 154442 226083 154445
rect 320869 154442 320935 154445
rect 87189 154440 90028 154442
rect 87189 154384 87194 154440
rect 87250 154384 90028 154440
rect 87189 154382 90028 154384
rect 223796 154440 226083 154442
rect 223796 154384 226022 154440
rect 226078 154384 226083 154440
rect 223796 154382 226083 154384
rect 317820 154440 320935 154442
rect 317820 154384 320874 154440
rect 320930 154384 320935 154440
rect 317820 154382 320935 154384
rect 87189 154379 87255 154382
rect 226017 154379 226083 154382
rect 320869 154379 320935 154382
rect 79737 153762 79803 153765
rect 76780 153760 79803 153762
rect 76780 153704 79742 153760
rect 79798 153704 79803 153760
rect 76780 153702 79803 153704
rect 79737 153699 79803 153702
rect 139721 153762 139787 153765
rect 172933 153762 172999 153765
rect 139721 153760 143020 153762
rect 139721 153704 139726 153760
rect 139782 153704 143020 153760
rect 139721 153702 143020 153704
rect 170804 153760 172999 153762
rect 170804 153704 172938 153760
rect 172994 153704 172999 153760
rect 170804 153702 172999 153704
rect 139721 153699 139787 153702
rect 172933 153699 172999 153702
rect 234021 153762 234087 153765
rect 266865 153762 266931 153765
rect 234021 153760 237044 153762
rect 234021 153704 234026 153760
rect 234082 153704 237044 153760
rect 234021 153702 237044 153704
rect 264828 153760 266931 153762
rect 264828 153704 266870 153760
rect 266926 153704 266931 153760
rect 264828 153702 266931 153704
rect 234021 153699 234087 153702
rect 266865 153699 266931 153702
rect 328413 153762 328479 153765
rect 328413 153760 331068 153762
rect 328413 153704 328418 153760
rect 328474 153704 331068 153760
rect 328413 153702 331068 153704
rect 328413 153699 328479 153702
rect 87189 153626 87255 153629
rect 132085 153626 132151 153629
rect 87189 153624 90028 153626
rect 87189 153568 87194 153624
rect 87250 153568 90028 153624
rect 87189 153566 90028 153568
rect 129772 153624 132151 153626
rect 129772 153568 132090 153624
rect 132146 153568 132151 153624
rect 129772 153566 132151 153568
rect 87189 153563 87255 153566
rect 132085 153563 132151 153566
rect 181949 153626 182015 153629
rect 225925 153626 225991 153629
rect 181949 153624 184052 153626
rect 181949 153568 181954 153624
rect 182010 153568 184052 153624
rect 181949 153566 184052 153568
rect 223796 153624 225991 153626
rect 223796 153568 225930 153624
rect 225986 153568 225991 153624
rect 223796 153566 225991 153568
rect 181949 153563 182015 153566
rect 225925 153563 225991 153566
rect 274869 153626 274935 153629
rect 321605 153626 321671 153629
rect 274869 153624 278076 153626
rect 274869 153568 274874 153624
rect 274930 153568 278076 153624
rect 274869 153566 278076 153568
rect 317820 153624 321671 153626
rect 317820 153568 321610 153624
rect 321666 153568 321671 153624
rect 317820 153566 321671 153568
rect 274869 153563 274935 153566
rect 321605 153563 321671 153566
rect 132545 153354 132611 153357
rect 129742 153352 132611 153354
rect 129742 153296 132550 153352
rect 132606 153296 132611 153352
rect 129742 153294 132611 153296
rect 49142 152884 49148 152948
rect 49212 152884 49218 152948
rect 49150 152644 49210 152884
rect 129742 152712 129802 153294
rect 132545 153291 132611 153294
rect 274961 153354 275027 153357
rect 274961 153352 278106 153354
rect 274961 153296 274966 153352
rect 275022 153296 278106 153352
rect 274961 153294 278106 153296
rect 274961 153291 275027 153294
rect 181397 153218 181463 153221
rect 181397 153216 184082 153218
rect 181397 153160 181402 153216
rect 181458 153160 184082 153216
rect 181397 153158 184082 153160
rect 181397 153155 181463 153158
rect 184022 152712 184082 153158
rect 278046 152712 278106 153294
rect 429429 152810 429495 152813
rect 434416 152810 434896 152840
rect 429429 152808 434896 152810
rect 429429 152752 429434 152808
rect 429490 152752 434896 152808
rect 429429 152750 434896 152752
rect 429429 152747 429495 152750
rect 434416 152720 434896 152750
rect 87189 152674 87255 152677
rect 225741 152674 225807 152677
rect 320501 152674 320567 152677
rect 360797 152674 360863 152677
rect 87189 152672 90028 152674
rect 87189 152616 87194 152672
rect 87250 152616 90028 152672
rect 87189 152614 90028 152616
rect 223796 152672 225807 152674
rect 223796 152616 225746 152672
rect 225802 152616 225807 152672
rect 223796 152614 225807 152616
rect 317820 152672 320567 152674
rect 317820 152616 320506 152672
rect 320562 152616 320567 152672
rect 317820 152614 320567 152616
rect 358852 152672 360863 152674
rect 358852 152616 360802 152672
rect 360858 152616 360863 152672
rect 358852 152614 360863 152616
rect 87189 152611 87255 152614
rect 225741 152611 225807 152614
rect 320501 152611 320567 152614
rect 360797 152611 360863 152614
rect 79737 152402 79803 152405
rect 76780 152400 79803 152402
rect 76780 152344 79742 152400
rect 79798 152344 79803 152400
rect 76780 152342 79803 152344
rect 79737 152339 79803 152342
rect 139629 152402 139695 152405
rect 173209 152402 173275 152405
rect 139629 152400 143020 152402
rect 139629 152344 139634 152400
rect 139690 152344 143020 152400
rect 139629 152342 143020 152344
rect 170804 152400 173275 152402
rect 170804 152344 173214 152400
rect 173270 152344 173275 152400
rect 170804 152342 173275 152344
rect 139629 152339 139695 152342
rect 173209 152339 173275 152342
rect 232917 152402 232983 152405
rect 266957 152402 267023 152405
rect 232917 152400 237044 152402
rect 232917 152344 232922 152400
rect 232978 152344 237044 152400
rect 232917 152342 237044 152344
rect 264828 152400 267023 152402
rect 264828 152344 266962 152400
rect 267018 152344 267023 152400
rect 264828 152342 267023 152344
rect 232917 152339 232983 152342
rect 266957 152339 267023 152342
rect 328413 152402 328479 152405
rect 328413 152400 331068 152402
rect 328413 152344 328418 152400
rect 328474 152344 331068 152400
rect 328413 152342 331068 152344
rect 328413 152339 328479 152342
rect 132637 152266 132703 152269
rect 129742 152264 132703 152266
rect 129742 152208 132642 152264
rect 132698 152208 132703 152264
rect 129742 152206 132703 152208
rect 129742 151896 129802 152206
rect 132637 152203 132703 152206
rect 182317 152130 182383 152133
rect 274869 152130 274935 152133
rect 182317 152128 184082 152130
rect 182317 152072 182322 152128
rect 182378 152072 184082 152128
rect 182317 152070 184082 152072
rect 182317 152067 182383 152070
rect 184022 151896 184082 152070
rect 274869 152128 278106 152130
rect 274869 152072 274874 152128
rect 274930 152072 278106 152128
rect 274869 152070 278106 152072
rect 274869 152067 274935 152070
rect 278046 151896 278106 152070
rect 87465 151858 87531 151861
rect 226109 151858 226175 151861
rect 320777 151858 320843 151861
rect 87465 151856 90028 151858
rect 87465 151800 87470 151856
rect 87526 151800 90028 151856
rect 87465 151798 90028 151800
rect 223796 151856 226175 151858
rect 223796 151800 226114 151856
rect 226170 151800 226175 151856
rect 223796 151798 226175 151800
rect 317820 151856 320843 151858
rect 317820 151800 320782 151856
rect 320838 151800 320843 151856
rect 317820 151798 320843 151800
rect 87465 151795 87531 151798
rect 226109 151795 226175 151798
rect 320777 151795 320843 151798
rect 87005 150906 87071 150909
rect 131901 150906 131967 150909
rect 87005 150904 90028 150906
rect 87005 150848 87010 150904
rect 87066 150848 90028 150904
rect 87005 150846 90028 150848
rect 129772 150904 131967 150906
rect 129772 150848 131906 150904
rect 131962 150848 131967 150904
rect 129772 150846 131967 150848
rect 87005 150843 87071 150846
rect 131901 150843 131967 150846
rect 140457 150906 140523 150909
rect 174037 150906 174103 150909
rect 140457 150904 143020 150906
rect 140457 150848 140462 150904
rect 140518 150848 143020 150904
rect 140457 150846 143020 150848
rect 170804 150904 174103 150906
rect 170804 150848 174042 150904
rect 174098 150848 174103 150904
rect 170804 150846 174103 150848
rect 140457 150843 140523 150846
rect 174037 150843 174103 150846
rect 182317 150906 182383 150909
rect 226201 150906 226267 150909
rect 182317 150904 184052 150906
rect 182317 150848 182322 150904
rect 182378 150848 184052 150904
rect 182317 150846 184052 150848
rect 223796 150904 226267 150906
rect 223796 150848 226206 150904
rect 226262 150848 226267 150904
rect 223796 150846 226267 150848
rect 182317 150843 182383 150846
rect 226201 150843 226267 150846
rect 233469 150906 233535 150909
rect 266589 150906 266655 150909
rect 233469 150904 237044 150906
rect 233469 150848 233474 150904
rect 233530 150848 237044 150904
rect 233469 150846 237044 150848
rect 264828 150904 266655 150906
rect 264828 150848 266594 150904
rect 266650 150848 266655 150904
rect 264828 150846 266655 150848
rect 233469 150843 233535 150846
rect 266589 150843 266655 150846
rect 274869 150906 274935 150909
rect 321053 150906 321119 150909
rect 274869 150904 278076 150906
rect 274869 150848 274874 150904
rect 274930 150848 278076 150904
rect 274869 150846 278076 150848
rect 317820 150904 321119 150906
rect 317820 150848 321058 150904
rect 321114 150848 321119 150904
rect 317820 150846 321119 150848
rect 274869 150843 274935 150846
rect 321053 150843 321119 150846
rect 328413 150906 328479 150909
rect 328413 150904 331068 150906
rect 328413 150848 328418 150904
rect 328474 150848 331068 150904
rect 328413 150846 331068 150848
rect 328413 150843 328479 150846
rect 77253 150838 77319 150841
rect 76780 150836 77319 150838
rect 76780 150780 77258 150836
rect 77314 150780 77319 150836
rect 76780 150778 77319 150780
rect 77253 150775 77319 150778
rect 182225 150634 182291 150637
rect 274317 150634 274383 150637
rect 182225 150632 184082 150634
rect 182225 150576 182230 150632
rect 182286 150576 184082 150632
rect 182225 150574 184082 150576
rect 182225 150571 182291 150574
rect 131717 150498 131783 150501
rect 129742 150496 131783 150498
rect 129742 150440 131722 150496
rect 131778 150440 131783 150496
rect 129742 150438 131783 150440
rect 129742 150128 129802 150438
rect 131717 150435 131783 150438
rect 184022 150128 184082 150574
rect 274317 150632 278106 150634
rect 274317 150576 274322 150632
rect 274378 150576 278106 150632
rect 274317 150574 278106 150576
rect 274317 150571 274383 150574
rect 278046 150128 278106 150574
rect 87189 150090 87255 150093
rect 225557 150090 225623 150093
rect 321605 150090 321671 150093
rect 87189 150088 90028 150090
rect 87189 150032 87194 150088
rect 87250 150032 90028 150088
rect 87189 150030 90028 150032
rect 223796 150088 225623 150090
rect 223796 150032 225562 150088
rect 225618 150032 225623 150088
rect 223796 150030 225623 150032
rect 317820 150088 321671 150090
rect 317820 150032 321610 150088
rect 321666 150032 321671 150088
rect 317820 150030 321671 150032
rect 87189 150027 87255 150030
rect 225557 150027 225623 150030
rect 321605 150027 321671 150030
rect 139629 149546 139695 149549
rect 174037 149546 174103 149549
rect 139629 149544 143020 149546
rect 9896 149274 10376 149304
rect 12853 149274 12919 149277
rect 9896 149272 12919 149274
rect 9896 149216 12858 149272
rect 12914 149216 12919 149272
rect 9896 149214 12919 149216
rect 9896 149184 10376 149214
rect 12853 149211 12919 149214
rect 49150 149004 49210 149516
rect 139629 149488 139634 149544
rect 139690 149488 143020 149544
rect 139629 149486 143020 149488
rect 170804 149544 174103 149546
rect 170804 149488 174042 149544
rect 174098 149488 174103 149544
rect 170804 149486 174103 149488
rect 139629 149483 139695 149486
rect 174037 149483 174103 149486
rect 232733 149546 232799 149549
rect 266589 149546 266655 149549
rect 232733 149544 237044 149546
rect 232733 149488 232738 149544
rect 232794 149488 237044 149544
rect 232733 149486 237044 149488
rect 264828 149544 266655 149546
rect 264828 149488 266594 149544
rect 266650 149488 266655 149544
rect 264828 149486 266655 149488
rect 232733 149483 232799 149486
rect 266589 149483 266655 149486
rect 274225 149546 274291 149549
rect 328413 149546 328479 149549
rect 360981 149546 361047 149549
rect 274225 149544 278106 149546
rect 274225 149488 274230 149544
rect 274286 149488 278106 149544
rect 274225 149486 278106 149488
rect 274225 149483 274291 149486
rect 49142 148940 49148 149004
rect 49212 148940 49218 149004
rect 76750 149002 76810 149448
rect 278046 149176 278106 149486
rect 328413 149544 331068 149546
rect 328413 149488 328418 149544
rect 328474 149488 331068 149544
rect 328413 149486 331068 149488
rect 358852 149544 361047 149546
rect 358852 149488 360986 149544
rect 361042 149488 361047 149544
rect 358852 149486 361047 149488
rect 328413 149483 328479 149486
rect 360981 149483 361047 149486
rect 87189 149138 87255 149141
rect 131349 149138 131415 149141
rect 225281 149138 225347 149141
rect 321605 149138 321671 149141
rect 87189 149136 90028 149138
rect 87189 149080 87194 149136
rect 87250 149080 90028 149136
rect 87189 149078 90028 149080
rect 129772 149136 131415 149138
rect 129772 149080 131354 149136
rect 131410 149080 131415 149136
rect 223796 149136 225347 149138
rect 129772 149078 131415 149080
rect 87189 149075 87255 149078
rect 131349 149075 131415 149078
rect 78909 149002 78975 149005
rect 76750 149000 78975 149002
rect 76750 148944 78914 149000
rect 78970 148944 78975 149000
rect 76750 148942 78975 148944
rect 78909 148939 78975 148942
rect 131625 148866 131691 148869
rect 129742 148864 131691 148866
rect 129742 148808 131630 148864
rect 131686 148808 131691 148864
rect 129742 148806 131691 148808
rect 76558 148532 76564 148596
rect 76628 148594 76634 148596
rect 76977 148594 77043 148597
rect 76628 148592 77043 148594
rect 76628 148536 76982 148592
rect 77038 148536 77043 148592
rect 76628 148534 77043 148536
rect 76628 148532 76634 148534
rect 76977 148531 77043 148534
rect 129742 148360 129802 148806
rect 131625 148803 131691 148806
rect 180385 148594 180451 148597
rect 184022 148594 184082 149108
rect 223796 149080 225286 149136
rect 225342 149080 225347 149136
rect 223796 149078 225347 149080
rect 317820 149136 321671 149138
rect 317820 149080 321610 149136
rect 321666 149080 321671 149136
rect 317820 149078 321671 149080
rect 225281 149075 225347 149078
rect 321605 149075 321671 149078
rect 274409 148866 274475 148869
rect 274409 148864 278106 148866
rect 274409 148808 274414 148864
rect 274470 148808 278106 148864
rect 274409 148806 278106 148808
rect 274409 148803 274475 148806
rect 180385 148592 184082 148594
rect 180385 148536 180390 148592
rect 180446 148536 184082 148592
rect 180385 148534 184082 148536
rect 180385 148531 180451 148534
rect 278046 148360 278106 148806
rect 87097 148322 87163 148325
rect 182317 148322 182383 148325
rect 225189 148322 225255 148325
rect 321697 148322 321763 148325
rect 87097 148320 90028 148322
rect 87097 148264 87102 148320
rect 87158 148264 90028 148320
rect 87097 148262 90028 148264
rect 182317 148320 184052 148322
rect 182317 148264 182322 148320
rect 182378 148264 184052 148320
rect 182317 148262 184052 148264
rect 223796 148320 225255 148322
rect 223796 148264 225194 148320
rect 225250 148264 225255 148320
rect 223796 148262 225255 148264
rect 317820 148320 321763 148322
rect 317820 148264 321702 148320
rect 321758 148264 321763 148320
rect 317820 148262 321763 148264
rect 87097 148259 87163 148262
rect 182317 148259 182383 148262
rect 225189 148259 225255 148262
rect 321697 148259 321763 148262
rect 138893 148186 138959 148189
rect 174037 148186 174103 148189
rect 138893 148184 143020 148186
rect 138893 148128 138898 148184
rect 138954 148128 143020 148184
rect 138893 148126 143020 148128
rect 170804 148184 174103 148186
rect 170804 148128 174042 148184
rect 174098 148128 174103 148184
rect 170804 148126 174103 148128
rect 138893 148123 138959 148126
rect 174037 148123 174103 148126
rect 233469 148186 233535 148189
rect 266589 148186 266655 148189
rect 233469 148184 237044 148186
rect 233469 148128 233474 148184
rect 233530 148128 237044 148184
rect 233469 148126 237044 148128
rect 264828 148184 266655 148186
rect 264828 148128 266594 148184
rect 266650 148128 266655 148184
rect 264828 148126 266655 148128
rect 233469 148123 233535 148126
rect 266589 148123 266655 148126
rect 328413 148186 328479 148189
rect 328413 148184 331068 148186
rect 328413 148128 328418 148184
rect 328474 148128 331068 148184
rect 328413 148126 331068 148128
rect 328413 148123 328479 148126
rect 76750 147914 76810 148088
rect 78909 147914 78975 147917
rect 76750 147912 78975 147914
rect 76750 147856 78914 147912
rect 78970 147856 78975 147912
rect 76750 147854 78975 147856
rect 78909 147851 78975 147854
rect 236822 147852 236828 147916
rect 236892 147914 236898 147916
rect 237190 147914 237196 147916
rect 236892 147854 237196 147914
rect 236892 147852 236898 147854
rect 237190 147852 237196 147854
rect 237260 147852 237266 147916
rect 80105 146690 80171 146693
rect 76780 146688 80171 146690
rect 76780 146632 80110 146688
rect 80166 146632 80171 146688
rect 76780 146630 80171 146632
rect 80105 146627 80171 146630
rect 140549 146690 140615 146693
rect 173853 146690 173919 146693
rect 140549 146688 143020 146690
rect 140549 146632 140554 146688
rect 140610 146632 143020 146688
rect 140549 146630 143020 146632
rect 170804 146688 173919 146690
rect 170804 146632 173858 146688
rect 173914 146632 173919 146688
rect 170804 146630 173919 146632
rect 140549 146627 140615 146630
rect 173853 146627 173919 146630
rect 233469 146690 233535 146693
rect 267877 146690 267943 146693
rect 233469 146688 237044 146690
rect 233469 146632 233474 146688
rect 233530 146632 237044 146688
rect 233469 146630 237044 146632
rect 264828 146688 267943 146690
rect 264828 146632 267882 146688
rect 267938 146632 267943 146688
rect 264828 146630 267943 146632
rect 233469 146627 233535 146630
rect 267877 146627 267943 146630
rect 327217 146690 327283 146693
rect 327217 146688 331068 146690
rect 327217 146632 327222 146688
rect 327278 146632 331068 146688
rect 327217 146630 331068 146632
rect 327217 146627 327283 146630
rect 360889 146418 360955 146421
rect 358852 146416 360955 146418
rect 49150 145876 49210 146388
rect 358852 146360 360894 146416
rect 360950 146360 360955 146416
rect 358852 146358 360955 146360
rect 360889 146355 360955 146358
rect 49142 145812 49148 145876
rect 49212 145812 49218 145876
rect 76558 145812 76564 145876
rect 76628 145874 76634 145876
rect 76885 145874 76951 145877
rect 76628 145872 76951 145874
rect 76628 145816 76890 145872
rect 76946 145816 76951 145872
rect 76628 145814 76951 145816
rect 76628 145812 76634 145814
rect 76885 145811 76951 145814
rect 79369 145330 79435 145333
rect 76780 145328 79435 145330
rect 76780 145272 79374 145328
rect 79430 145272 79435 145328
rect 76780 145270 79435 145272
rect 79369 145267 79435 145270
rect 140549 145330 140615 145333
rect 173761 145330 173827 145333
rect 140549 145328 143020 145330
rect 140549 145272 140554 145328
rect 140610 145272 143020 145328
rect 140549 145270 143020 145272
rect 170804 145328 173827 145330
rect 170804 145272 173766 145328
rect 173822 145272 173827 145328
rect 170804 145270 173827 145272
rect 140549 145267 140615 145270
rect 173761 145267 173827 145270
rect 233469 145330 233535 145333
rect 266773 145330 266839 145333
rect 233469 145328 237044 145330
rect 233469 145272 233474 145328
rect 233530 145272 237044 145328
rect 233469 145270 237044 145272
rect 264828 145328 266839 145330
rect 264828 145272 266778 145328
rect 266834 145272 266839 145328
rect 264828 145270 266839 145272
rect 233469 145267 233535 145270
rect 266773 145267 266839 145270
rect 327861 145330 327927 145333
rect 327861 145328 331068 145330
rect 327861 145272 327866 145328
rect 327922 145272 331068 145328
rect 327861 145270 331068 145272
rect 327861 145267 327927 145270
rect 176286 145132 176292 145196
rect 176356 145194 176362 145196
rect 187142 145194 187148 145196
rect 176356 145134 187148 145194
rect 176356 145132 176362 145134
rect 187142 145132 187148 145134
rect 187212 145132 187218 145196
rect 192897 144650 192963 144653
rect 197630 144650 197636 144652
rect 192897 144648 197636 144650
rect 192897 144592 192902 144648
rect 192958 144592 197636 144648
rect 192897 144590 197636 144592
rect 192897 144587 192963 144590
rect 197630 144588 197636 144590
rect 197700 144588 197706 144652
rect 196158 144452 196164 144516
rect 196228 144514 196234 144516
rect 203753 144514 203819 144517
rect 196228 144512 203819 144514
rect 196228 144456 203758 144512
rect 203814 144456 203819 144512
rect 196228 144454 203819 144456
rect 196228 144452 196234 144454
rect 203753 144451 203819 144454
rect 289998 144452 290004 144516
rect 290068 144514 290074 144516
rect 290509 144514 290575 144517
rect 290068 144512 290575 144514
rect 290068 144456 290514 144512
rect 290570 144456 290575 144512
rect 290068 144454 290575 144456
rect 290068 144452 290074 144454
rect 290509 144451 290575 144454
rect 98270 144180 98276 144244
rect 98340 144242 98346 144244
rect 98873 144242 98939 144245
rect 142246 144242 142252 144244
rect 98340 144240 142252 144242
rect 98340 144184 98878 144240
rect 98934 144184 142252 144240
rect 98340 144182 142252 144184
rect 98340 144180 98346 144182
rect 98873 144179 98939 144182
rect 142246 144180 142252 144182
rect 142316 144180 142322 144244
rect 76977 144108 77043 144109
rect 76926 144044 76932 144108
rect 76996 144106 77043 144108
rect 95285 144106 95351 144109
rect 142062 144106 142068 144108
rect 76996 144104 77088 144106
rect 77038 144048 77088 144104
rect 76996 144046 77088 144048
rect 95285 144104 142068 144106
rect 95285 144048 95290 144104
rect 95346 144048 142068 144104
rect 95285 144046 142068 144048
rect 76996 144044 77043 144046
rect 76977 144043 77043 144044
rect 95285 144043 95351 144046
rect 142062 144044 142068 144046
rect 142132 144044 142138 144108
rect 196485 144106 196551 144109
rect 196853 144106 196919 144109
rect 236086 144106 236092 144108
rect 196485 144104 236092 144106
rect 196485 144048 196490 144104
rect 196546 144048 196858 144104
rect 196914 144048 236092 144104
rect 196485 144046 236092 144048
rect 196485 144043 196551 144046
rect 196853 144043 196919 144046
rect 236086 144044 236092 144046
rect 236156 144044 236162 144108
rect 140549 143970 140615 143973
rect 173945 143970 174011 143973
rect 197681 143972 197747 143973
rect 140549 143968 143020 143970
rect 140549 143912 140554 143968
rect 140610 143912 143020 143968
rect 140549 143910 143020 143912
rect 170804 143968 174011 143970
rect 170804 143912 173950 143968
rect 174006 143912 174011 143968
rect 170804 143910 174011 143912
rect 140549 143907 140615 143910
rect 173945 143907 174011 143910
rect 197630 143908 197636 143972
rect 197700 143970 197747 143972
rect 233469 143970 233535 143973
rect 267785 143970 267851 143973
rect 197700 143968 197792 143970
rect 197742 143912 197792 143968
rect 197700 143910 197792 143912
rect 233469 143968 237044 143970
rect 233469 143912 233474 143968
rect 233530 143912 237044 143968
rect 233469 143910 237044 143912
rect 264828 143968 267851 143970
rect 264828 143912 267790 143968
rect 267846 143912 267851 143968
rect 264828 143910 267851 143912
rect 197700 143908 197747 143910
rect 197681 143907 197747 143908
rect 233469 143907 233535 143910
rect 267785 143907 267851 143910
rect 327309 143970 327375 143973
rect 327309 143968 331068 143970
rect 327309 143912 327314 143968
rect 327370 143912 331068 143968
rect 327309 143910 331068 143912
rect 327309 143907 327375 143910
rect 76750 143562 76810 143872
rect 78909 143562 78975 143565
rect 76750 143560 78975 143562
rect 76750 143504 78914 143560
rect 78970 143504 78975 143560
rect 76750 143502 78975 143504
rect 78909 143499 78975 143502
rect 47077 143426 47143 143429
rect 361073 143426 361139 143429
rect 47077 143424 48996 143426
rect 47077 143368 47082 143424
rect 47138 143368 48996 143424
rect 47077 143366 48996 143368
rect 358852 143424 361139 143426
rect 358852 143368 361078 143424
rect 361134 143368 361139 143424
rect 358852 143366 361139 143368
rect 47077 143363 47143 143366
rect 361073 143363 361139 143366
rect 109729 143290 109795 143293
rect 110414 143290 110420 143292
rect 109729 143288 110420 143290
rect 109729 143232 109734 143288
rect 109790 143232 110420 143288
rect 109729 143230 110420 143232
rect 109729 143227 109795 143230
rect 110414 143228 110420 143230
rect 110484 143290 110490 143292
rect 136910 143290 136916 143292
rect 110484 143230 136916 143290
rect 110484 143228 110490 143230
rect 136910 143228 136916 143230
rect 136980 143290 136986 143292
rect 137145 143290 137211 143293
rect 136980 143288 137211 143290
rect 136980 143232 137150 143288
rect 137206 143232 137211 143288
rect 136980 143230 137211 143232
rect 136980 143228 136986 143230
rect 137145 143227 137211 143230
rect 210142 143092 210148 143156
rect 210212 143154 210218 143156
rect 211021 143154 211087 143157
rect 294281 143156 294347 143157
rect 210212 143152 211087 143154
rect 210212 143096 211026 143152
rect 211082 143096 211087 143152
rect 210212 143094 211087 143096
rect 210212 143092 210218 143094
rect 211021 143091 211087 143094
rect 294230 143092 294236 143156
rect 294300 143154 294347 143156
rect 294300 143152 294392 143154
rect 294342 143096 294392 143152
rect 294300 143094 294392 143096
rect 294300 143092 294347 143094
rect 294281 143091 294347 143092
rect 88569 142882 88635 142885
rect 89622 142882 89628 142884
rect 88569 142880 89628 142882
rect 88569 142824 88574 142880
rect 88630 142824 89628 142880
rect 88569 142822 89628 142824
rect 88569 142819 88635 142822
rect 89622 142820 89628 142822
rect 89692 142820 89698 142884
rect 140273 142610 140339 142613
rect 173577 142610 173643 142613
rect 267233 142610 267299 142613
rect 140273 142608 143020 142610
rect 140273 142552 140278 142608
rect 140334 142552 143020 142608
rect 140273 142550 143020 142552
rect 170804 142608 173643 142610
rect 170804 142552 173582 142608
rect 173638 142552 173643 142608
rect 170804 142550 173643 142552
rect 264828 142608 267299 142610
rect 264828 142552 267238 142608
rect 267294 142552 267299 142608
rect 264828 142550 267299 142552
rect 140273 142547 140339 142550
rect 173577 142547 173643 142550
rect 267233 142547 267299 142550
rect 73798 142412 73804 142476
rect 73868 142474 73874 142476
rect 74350 142474 74356 142476
rect 73868 142414 74356 142474
rect 73868 142412 73874 142414
rect 74350 142412 74356 142414
rect 74420 142474 74426 142476
rect 74902 142474 74908 142476
rect 74420 142414 74908 142474
rect 74420 142412 74426 142414
rect 74902 142412 74908 142414
rect 74972 142412 74978 142476
rect 73941 142202 74007 142205
rect 74534 142202 74540 142204
rect 73941 142200 74540 142202
rect 73941 142144 73946 142200
rect 74002 142144 74540 142200
rect 73941 142142 74540 142144
rect 73941 142139 74007 142142
rect 74534 142140 74540 142142
rect 74604 142140 74610 142204
rect 75413 142202 75479 142205
rect 75638 142202 75644 142204
rect 75413 142200 75644 142202
rect 75413 142144 75418 142200
rect 75474 142144 75644 142200
rect 75413 142142 75644 142144
rect 75413 142139 75479 142142
rect 75638 142140 75644 142142
rect 75708 142140 75714 142204
rect 73982 142004 73988 142068
rect 74052 142066 74058 142068
rect 74534 142066 74540 142068
rect 74052 142006 74540 142066
rect 74052 142004 74058 142006
rect 74534 142004 74540 142006
rect 74604 142004 74610 142068
rect 75270 142004 75276 142068
rect 75340 142066 75346 142068
rect 76057 142066 76123 142069
rect 75340 142064 76123 142066
rect 75340 142008 76062 142064
rect 76118 142008 76123 142064
rect 75340 142006 76123 142008
rect 75340 142004 75346 142006
rect 74542 141930 74602 142004
rect 76057 142003 76123 142006
rect 76006 141930 76012 141932
rect 74542 141870 76012 141930
rect 76006 141868 76012 141870
rect 76076 141868 76082 141932
rect 76750 141930 76810 142512
rect 142430 142276 142436 142340
rect 142500 142338 142506 142340
rect 151814 142338 151820 142340
rect 142500 142278 151820 142338
rect 142500 142276 142506 142278
rect 150672 142205 150732 142278
rect 151814 142276 151820 142278
rect 151884 142276 151890 142340
rect 142246 142140 142252 142204
rect 142316 142202 142322 142204
rect 144086 142202 144092 142204
rect 142316 142142 144092 142202
rect 142316 142140 142322 142142
rect 144086 142140 144092 142142
rect 144156 142202 144162 142204
rect 147909 142202 147975 142205
rect 144156 142200 147975 142202
rect 144156 142144 147914 142200
rect 147970 142144 147975 142200
rect 144156 142142 147975 142144
rect 144156 142140 144162 142142
rect 147909 142139 147975 142142
rect 150669 142200 150735 142205
rect 150669 142144 150674 142200
rect 150730 142144 150735 142200
rect 150669 142139 150735 142144
rect 167638 142140 167644 142204
rect 167708 142202 167714 142204
rect 167965 142202 168031 142205
rect 167708 142200 168031 142202
rect 167708 142144 167970 142200
rect 168026 142144 168031 142200
rect 167708 142142 168031 142144
rect 167708 142140 167714 142142
rect 167965 142139 168031 142142
rect 142062 142004 142068 142068
rect 142132 142066 142138 142068
rect 146805 142066 146871 142069
rect 142132 142064 146871 142066
rect 142132 142008 146810 142064
rect 146866 142008 146871 142064
rect 142132 142006 146871 142008
rect 142132 142004 142138 142006
rect 146805 142003 146871 142006
rect 219669 142068 219735 142069
rect 219669 142064 219716 142068
rect 219780 142066 219786 142068
rect 233469 142066 233535 142069
rect 237014 142066 237074 142512
rect 238294 142412 238300 142476
rect 238364 142474 238370 142476
rect 242526 142474 242532 142476
rect 238364 142414 242532 142474
rect 238364 142412 238370 142414
rect 242526 142412 242532 142414
rect 242596 142412 242602 142476
rect 238110 142140 238116 142204
rect 238180 142202 238186 142204
rect 242025 142202 242091 142205
rect 238180 142200 242091 142202
rect 238180 142144 242030 142200
rect 242086 142144 242091 142200
rect 238180 142142 242091 142144
rect 238180 142140 238186 142142
rect 242025 142139 242091 142142
rect 261662 142140 261668 142204
rect 261732 142202 261738 142204
rect 261897 142202 261963 142205
rect 261732 142200 261963 142202
rect 261732 142144 261902 142200
rect 261958 142144 261963 142200
rect 261732 142142 261963 142144
rect 261732 142140 261738 142142
rect 261897 142139 261963 142142
rect 219669 142008 219674 142064
rect 219669 142004 219716 142008
rect 219780 142006 219826 142066
rect 233469 142064 237074 142066
rect 233469 142008 233474 142064
rect 233530 142008 237074 142064
rect 233469 142006 237074 142008
rect 219780 142004 219786 142006
rect 219669 142003 219735 142004
rect 233469 142003 233535 142006
rect 78909 141930 78975 141933
rect 76750 141928 78975 141930
rect 76750 141872 78914 141928
rect 78970 141872 78975 141928
rect 76750 141870 78975 141872
rect 78909 141867 78975 141870
rect 105078 141868 105084 141932
rect 105148 141930 105154 141932
rect 106141 141930 106207 141933
rect 136869 141930 136935 141933
rect 105148 141928 136935 141930
rect 105148 141872 106146 141928
rect 106202 141872 136874 141928
rect 136930 141872 136935 141928
rect 105148 141870 136935 141872
rect 105148 141868 105154 141870
rect 106141 141867 106207 141870
rect 136869 141867 136935 141870
rect 200165 141930 200231 141933
rect 230750 141930 230756 141932
rect 200165 141928 230756 141930
rect 200165 141872 200170 141928
rect 200226 141872 230756 141928
rect 200165 141870 230756 141872
rect 200165 141867 200231 141870
rect 230750 141868 230756 141870
rect 230820 141868 230826 141932
rect 327309 141930 327375 141933
rect 331038 141930 331098 142512
rect 327309 141928 331098 141930
rect 327309 141872 327314 141928
rect 327370 141872 331098 141928
rect 327309 141870 331098 141872
rect 327309 141867 327375 141870
rect 74350 141732 74356 141796
rect 74420 141794 74426 141796
rect 76926 141794 76932 141796
rect 74420 141734 76932 141794
rect 74420 141732 74426 141734
rect 76926 141732 76932 141734
rect 76996 141794 77002 141796
rect 78214 141794 78220 141796
rect 76996 141734 78220 141794
rect 76996 141732 77002 141734
rect 78214 141732 78220 141734
rect 78284 141732 78290 141796
rect 167822 141732 167828 141796
rect 167892 141794 167898 141796
rect 168374 141794 168380 141796
rect 167892 141734 168380 141794
rect 167892 141732 167898 141734
rect 168374 141732 168380 141734
rect 168444 141794 168450 141796
rect 168517 141794 168583 141797
rect 168444 141792 168583 141794
rect 168444 141736 168522 141792
rect 168578 141736 168583 141792
rect 168444 141734 168583 141736
rect 168444 141732 168450 141734
rect 168517 141731 168583 141734
rect 237742 141732 237748 141796
rect 237812 141794 237818 141796
rect 241974 141794 241980 141796
rect 237812 141734 241980 141794
rect 237812 141732 237818 141734
rect 241974 141732 241980 141734
rect 242044 141794 242050 141796
rect 243221 141794 243287 141797
rect 256694 141794 256700 141796
rect 242044 141792 256700 141794
rect 242044 141736 243226 141792
rect 243282 141736 256700 141792
rect 242044 141734 256700 141736
rect 242044 141732 242050 141734
rect 243221 141731 243287 141734
rect 256694 141732 256700 141734
rect 256764 141732 256770 141796
rect 137329 141114 137395 141117
rect 149105 141116 149171 141117
rect 207249 141116 207315 141117
rect 137462 141114 137468 141116
rect 137329 141112 137468 141114
rect 137329 141056 137334 141112
rect 137390 141056 137468 141112
rect 137329 141054 137468 141056
rect 137329 141051 137395 141054
rect 137462 141052 137468 141054
rect 137532 141052 137538 141116
rect 149054 141052 149060 141116
rect 149124 141114 149171 141116
rect 149124 141112 149216 141114
rect 149166 141056 149216 141112
rect 149124 141054 149216 141056
rect 149124 141052 149171 141054
rect 207198 141052 207204 141116
rect 207268 141114 207315 141116
rect 207268 141112 207360 141114
rect 207310 141056 207360 141112
rect 207268 141054 207360 141056
rect 207268 141052 207315 141054
rect 296990 141052 296996 141116
rect 297060 141114 297066 141116
rect 301089 141114 301155 141117
rect 297060 141112 301155 141114
rect 297060 141056 301094 141112
rect 301150 141056 301155 141112
rect 297060 141054 301155 141056
rect 297060 141052 297066 141054
rect 149105 141051 149171 141052
rect 207249 141051 207315 141052
rect 301089 141051 301155 141054
rect 152049 140436 152115 140437
rect 151998 140372 152004 140436
rect 152068 140434 152115 140436
rect 152068 140432 152160 140434
rect 152110 140376 152160 140432
rect 152068 140374 152160 140376
rect 152068 140372 152115 140374
rect 152049 140371 152115 140372
rect 137237 140300 137303 140301
rect 137237 140296 137284 140300
rect 137348 140298 137354 140300
rect 429521 140298 429587 140301
rect 434416 140298 434896 140328
rect 137237 140240 137242 140296
rect 137237 140236 137284 140240
rect 137348 140238 137394 140298
rect 429521 140296 434896 140298
rect 429521 140240 429526 140296
rect 429582 140240 434896 140296
rect 429521 140238 434896 140240
rect 137348 140236 137354 140238
rect 137237 140235 137303 140236
rect 429521 140235 429587 140238
rect 434416 140208 434896 140238
rect 230750 139964 230756 140028
rect 230820 140026 230826 140028
rect 230985 140026 231051 140029
rect 230820 140024 231051 140026
rect 230820 139968 230990 140024
rect 231046 139968 231051 140024
rect 230820 139966 231051 139968
rect 230820 139964 230826 139966
rect 230985 139963 231051 139966
rect 147449 139890 147515 139893
rect 147766 139890 147772 139892
rect 147449 139888 147772 139890
rect 147449 139832 147454 139888
rect 147510 139832 147772 139888
rect 147449 139830 147772 139832
rect 147449 139827 147515 139830
rect 147766 139828 147772 139830
rect 147836 139828 147842 139892
rect 148185 139890 148251 139893
rect 148502 139890 148508 139892
rect 148185 139888 148508 139890
rect 148185 139832 148190 139888
rect 148246 139832 148508 139888
rect 148185 139830 148508 139832
rect 148185 139827 148251 139830
rect 148502 139828 148508 139830
rect 148572 139828 148578 139892
rect 152693 139890 152759 139893
rect 169110 139890 169116 139892
rect 152693 139888 169116 139890
rect 152693 139832 152698 139888
rect 152754 139832 169116 139888
rect 152693 139830 169116 139832
rect 152693 139827 152759 139830
rect 169110 139828 169116 139830
rect 169180 139828 169186 139892
rect 243078 139828 243084 139892
rect 243148 139890 243154 139892
rect 244049 139890 244115 139893
rect 262950 139890 262956 139892
rect 243148 139888 262956 139890
rect 243148 139832 244054 139888
rect 244110 139832 262956 139888
rect 243148 139830 262956 139832
rect 243148 139828 243154 139830
rect 244049 139827 244115 139830
rect 262950 139828 262956 139830
rect 263020 139828 263026 139892
rect 231445 139754 231511 139757
rect 241749 139754 241815 139757
rect 242526 139754 242532 139756
rect 231445 139752 242532 139754
rect 231445 139696 231450 139752
rect 231506 139696 241754 139752
rect 241810 139696 242532 139752
rect 231445 139694 242532 139696
rect 231445 139691 231511 139694
rect 241749 139691 241815 139694
rect 242526 139692 242532 139694
rect 242596 139692 242602 139756
rect 246349 139754 246415 139757
rect 251358 139754 251364 139756
rect 246349 139752 251364 139754
rect 246349 139696 246354 139752
rect 246410 139696 251364 139752
rect 246349 139694 251364 139696
rect 246349 139691 246415 139694
rect 251358 139692 251364 139694
rect 251428 139692 251434 139756
rect 52638 139556 52644 139620
rect 52708 139618 52714 139620
rect 53517 139618 53583 139621
rect 52708 139616 53583 139618
rect 52708 139560 53522 139616
rect 53578 139560 53583 139616
rect 52708 139558 53583 139560
rect 52708 139556 52714 139558
rect 53517 139555 53583 139558
rect 54529 139618 54595 139621
rect 54846 139618 54852 139620
rect 54529 139616 54852 139618
rect 54529 139560 54534 139616
rect 54590 139560 54852 139616
rect 54529 139558 54852 139560
rect 54529 139555 54595 139558
rect 54846 139556 54852 139558
rect 54916 139556 54922 139620
rect 350953 139618 351019 139621
rect 351638 139618 351644 139620
rect 350953 139616 351644 139618
rect 350953 139560 350958 139616
rect 351014 139560 351644 139616
rect 350953 139558 351644 139560
rect 350953 139555 351019 139558
rect 351638 139556 351644 139558
rect 351708 139556 351714 139620
rect 351822 139556 351828 139620
rect 351892 139618 351898 139620
rect 352057 139618 352123 139621
rect 351892 139616 352123 139618
rect 351892 139560 352062 139616
rect 352118 139560 352123 139616
rect 351892 139558 352123 139560
rect 351892 139556 351898 139558
rect 352057 139555 352123 139558
rect 73430 139420 73436 139484
rect 73500 139482 73506 139484
rect 74217 139482 74283 139485
rect 75137 139482 75203 139485
rect 73500 139480 75203 139482
rect 73500 139424 74222 139480
rect 74278 139424 75142 139480
rect 75198 139424 75203 139480
rect 73500 139422 75203 139424
rect 73500 139420 73506 139422
rect 74217 139419 74283 139422
rect 75137 139419 75203 139422
rect 252237 138530 252303 138533
rect 252646 138530 252652 138532
rect 252237 138528 252652 138530
rect 252237 138472 252242 138528
rect 252298 138472 252652 138528
rect 252237 138470 252652 138472
rect 252237 138467 252303 138470
rect 252646 138468 252652 138470
rect 252716 138468 252722 138532
rect 283149 138530 283215 138533
rect 284437 138530 284503 138533
rect 252838 138528 284503 138530
rect 252838 138472 283154 138528
rect 283210 138472 284442 138528
rect 284498 138472 284503 138528
rect 252838 138470 284503 138472
rect 249661 138396 249727 138397
rect 249661 138392 249708 138396
rect 249772 138394 249778 138396
rect 252838 138394 252898 138470
rect 283149 138467 283215 138470
rect 284437 138467 284503 138470
rect 249661 138336 249666 138392
rect 249661 138332 249708 138336
rect 249772 138334 252898 138394
rect 249772 138332 249778 138334
rect 249661 138331 249727 138332
rect 252646 137788 252652 137852
rect 252716 137850 252722 137852
rect 296949 137850 297015 137853
rect 298094 137850 298100 137852
rect 252716 137848 298100 137850
rect 252716 137792 296954 137848
rect 297010 137792 298100 137848
rect 252716 137790 298100 137792
rect 252716 137788 252722 137790
rect 296949 137787 297015 137790
rect 298094 137788 298100 137790
rect 298164 137788 298170 137852
rect 73614 137108 73620 137172
rect 73684 137170 73690 137172
rect 76057 137170 76123 137173
rect 73684 137168 76123 137170
rect 73684 137112 76062 137168
rect 76118 137112 76123 137168
rect 73684 137110 76123 137112
rect 73684 137108 73690 137110
rect 76057 137107 76123 137110
rect 9896 135946 10376 135976
rect 12853 135946 12919 135949
rect 9896 135944 12919 135946
rect 9896 135888 12858 135944
rect 12914 135888 12919 135944
rect 9896 135886 12919 135888
rect 9896 135856 10376 135886
rect 12853 135883 12919 135886
rect 249109 135810 249175 135813
rect 285909 135810 285975 135813
rect 286737 135810 286803 135813
rect 249109 135808 286803 135810
rect 249109 135752 249114 135808
rect 249170 135752 285914 135808
rect 285970 135752 286742 135808
rect 286798 135752 286803 135808
rect 249109 135750 286803 135752
rect 249109 135747 249175 135750
rect 285909 135747 285975 135750
rect 286737 135747 286803 135750
rect 197681 135130 197747 135133
rect 198550 135130 198556 135132
rect 197681 135128 198556 135130
rect 197681 135072 197686 135128
rect 197742 135072 198556 135128
rect 197681 135070 198556 135072
rect 197681 135067 197747 135070
rect 198550 135068 198556 135070
rect 198620 135068 198626 135132
rect 55214 134388 55220 134452
rect 55284 134450 55290 134452
rect 55541 134450 55607 134453
rect 249109 134452 249175 134453
rect 249109 134450 249156 134452
rect 55284 134448 55607 134450
rect 55284 134392 55546 134448
rect 55602 134392 55607 134448
rect 55284 134390 55607 134392
rect 249064 134448 249156 134450
rect 249064 134392 249114 134448
rect 249064 134390 249156 134392
rect 55284 134388 55290 134390
rect 55541 134387 55607 134390
rect 249109 134388 249156 134390
rect 249220 134388 249226 134452
rect 249109 134387 249175 134388
rect 351822 134252 351828 134316
rect 351892 134252 351898 134316
rect 351830 134178 351890 134252
rect 352558 134178 352564 134180
rect 351830 134118 352564 134178
rect 352558 134116 352564 134118
rect 352628 134116 352634 134180
rect 136869 132954 136935 132957
rect 231353 132954 231419 132957
rect 134710 132952 136935 132954
rect 134710 132896 136874 132952
rect 136930 132896 136935 132952
rect 134710 132894 136935 132896
rect 55398 132348 55404 132412
rect 55468 132410 55474 132412
rect 56093 132410 56159 132413
rect 55468 132408 56159 132410
rect 55468 132352 56098 132408
rect 56154 132352 56159 132408
rect 55468 132350 56159 132352
rect 55468 132348 55474 132350
rect 56093 132347 56159 132350
rect 134710 132312 134770 132894
rect 136869 132891 136935 132894
rect 228734 132952 231419 132954
rect 228734 132896 231358 132952
rect 231414 132896 231419 132952
rect 228734 132894 231419 132896
rect 178678 132484 178684 132548
rect 178748 132546 178754 132548
rect 182910 132546 182916 132548
rect 178748 132486 182916 132546
rect 178748 132484 178754 132486
rect 182910 132484 182916 132486
rect 182980 132484 182986 132548
rect 198550 132484 198556 132548
rect 198620 132546 198626 132548
rect 199286 132546 199292 132548
rect 198620 132486 199292 132546
rect 198620 132484 198626 132486
rect 199286 132484 199292 132486
rect 199356 132484 199362 132548
rect 228734 132312 228794 132894
rect 231353 132891 231419 132894
rect 298094 132484 298100 132548
rect 298164 132546 298170 132548
rect 324641 132546 324707 132549
rect 298164 132544 324707 132546
rect 298164 132488 324646 132544
rect 324702 132488 324707 132544
rect 298164 132486 324707 132488
rect 298164 132484 298170 132486
rect 324641 132483 324707 132486
rect 324549 132410 324615 132413
rect 322758 132408 324615 132410
rect 322758 132352 324554 132408
rect 324610 132352 324615 132408
rect 322758 132350 324615 132352
rect 322758 132312 322818 132350
rect 324549 132347 324615 132350
rect 246206 130172 246212 130236
rect 246276 130234 246282 130236
rect 246441 130234 246507 130237
rect 246276 130232 246507 130234
rect 246276 130176 246446 130232
rect 246502 130176 246507 130232
rect 246276 130174 246507 130176
rect 246276 130172 246282 130174
rect 246441 130171 246507 130174
rect 137237 129826 137303 129829
rect 231077 129826 231143 129829
rect 325101 129826 325167 129829
rect 134710 129824 137303 129826
rect 134710 129768 137242 129824
rect 137298 129768 137303 129824
rect 134710 129766 137303 129768
rect 134710 129184 134770 129766
rect 137237 129763 137303 129766
rect 228734 129824 231143 129826
rect 228734 129768 231082 129824
rect 231138 129768 231143 129824
rect 228734 129766 231143 129768
rect 228734 129184 228794 129766
rect 231077 129763 231143 129766
rect 322758 129824 325167 129826
rect 322758 129768 325106 129824
rect 325162 129768 325167 129824
rect 322758 129766 325167 129768
rect 242025 129556 242091 129557
rect 241974 129554 241980 129556
rect 241934 129494 241980 129554
rect 242044 129552 242091 129556
rect 242086 129496 242091 129552
rect 241974 129492 241980 129494
rect 242044 129492 242091 129496
rect 242025 129491 242091 129492
rect 322758 129184 322818 129766
rect 325101 129763 325167 129766
rect 428693 127786 428759 127789
rect 434416 127786 434896 127816
rect 428693 127784 434896 127786
rect 428693 127728 428698 127784
rect 428754 127728 434896 127784
rect 428693 127726 434896 127728
rect 428693 127723 428759 127726
rect 434416 127696 434896 127726
rect 38797 127514 38863 127517
rect 84705 127516 84771 127517
rect 84654 127514 84660 127516
rect 35748 127512 38863 127514
rect 35748 127456 38802 127512
rect 38858 127456 38863 127512
rect 35748 127454 38863 127456
rect 84614 127454 84660 127514
rect 84724 127512 84771 127516
rect 84766 127456 84771 127512
rect 38797 127451 38863 127454
rect 84654 127452 84660 127454
rect 84724 127452 84771 127456
rect 252646 127452 252652 127516
rect 252716 127514 252722 127516
rect 259638 127514 259644 127516
rect 252716 127454 259644 127514
rect 252716 127452 252722 127454
rect 259638 127452 259644 127454
rect 259708 127452 259714 127516
rect 84705 127451 84771 127452
rect 48457 127242 48523 127245
rect 55398 127242 55404 127244
rect 48457 127240 55404 127242
rect 48457 127184 48462 127240
rect 48518 127184 55404 127240
rect 48457 127182 55404 127184
rect 48457 127179 48523 127182
rect 55398 127180 55404 127182
rect 55468 127180 55474 127244
rect 405969 126970 406035 126973
rect 409054 126970 409114 127484
rect 405969 126968 409114 126970
rect 70678 126426 70738 126940
rect 405969 126912 405974 126968
rect 406030 126912 409114 126968
rect 405969 126910 409114 126912
rect 405969 126907 406035 126910
rect 248598 126772 248604 126836
rect 248668 126834 248674 126836
rect 249702 126834 249708 126836
rect 248668 126774 249708 126834
rect 248668 126772 248674 126774
rect 249702 126772 249708 126774
rect 249772 126772 249778 126836
rect 74309 126426 74375 126429
rect 70678 126424 74375 126426
rect 70678 126368 74314 126424
rect 74370 126368 74375 126424
rect 70678 126366 74375 126368
rect 74309 126363 74375 126366
rect 52597 126290 52663 126293
rect 356197 126290 356263 126293
rect 427313 126290 427379 126293
rect 52597 126288 55068 126290
rect 16073 126154 16139 126157
rect 19894 126154 19954 126260
rect 52597 126232 52602 126288
rect 52658 126232 55068 126288
rect 52597 126230 55068 126232
rect 352780 126288 356263 126290
rect 352780 126232 356202 126288
rect 356258 126232 356263 126288
rect 352780 126230 356263 126232
rect 424724 126288 427379 126290
rect 424724 126232 427318 126288
rect 427374 126232 427379 126288
rect 424724 126230 427379 126232
rect 52597 126227 52663 126230
rect 356197 126227 356263 126230
rect 427313 126227 427379 126230
rect 16073 126152 19954 126154
rect 16073 126096 16078 126152
rect 16134 126096 19954 126152
rect 16073 126094 19954 126096
rect 16073 126091 16139 126094
rect 134710 126018 134770 126052
rect 137053 126018 137119 126021
rect 134710 126016 137119 126018
rect 134710 125960 137058 126016
rect 137114 125960 137119 126016
rect 134710 125958 137119 125960
rect 228734 126018 228794 126052
rect 231445 126018 231511 126021
rect 228734 126016 231511 126018
rect 228734 125960 231450 126016
rect 231506 125960 231511 126016
rect 228734 125958 231511 125960
rect 322758 126018 322818 126056
rect 324641 126018 324707 126021
rect 322758 126016 324707 126018
rect 322758 125960 324646 126016
rect 324702 125960 324707 126016
rect 322758 125958 324707 125960
rect 137053 125955 137119 125958
rect 231445 125955 231511 125958
rect 324641 125955 324707 125958
rect 38245 125610 38311 125613
rect 35718 125608 38311 125610
rect 35718 125552 38250 125608
rect 38306 125552 38311 125608
rect 35718 125550 38311 125552
rect 35718 125104 35778 125550
rect 38245 125547 38311 125550
rect 405969 125610 406035 125613
rect 405969 125608 408930 125610
rect 405969 125552 405974 125608
rect 406030 125552 408930 125608
rect 405969 125550 408930 125552
rect 405969 125547 406035 125550
rect 84478 125478 85060 125538
rect 178318 125482 178900 125542
rect 272342 125482 272924 125542
rect 82681 125474 82747 125477
rect 84478 125474 84538 125478
rect 82681 125472 84538 125474
rect 82681 125416 82686 125472
rect 82742 125416 84538 125472
rect 82681 125414 84538 125416
rect 175509 125474 175575 125477
rect 178318 125474 178378 125482
rect 175509 125472 178378 125474
rect 175509 125416 175514 125472
rect 175570 125416 178378 125472
rect 175509 125414 178378 125416
rect 270361 125474 270427 125477
rect 272342 125474 272402 125482
rect 270361 125472 272402 125474
rect 270361 125416 270366 125472
rect 270422 125416 272402 125472
rect 270361 125414 272402 125416
rect 82681 125411 82747 125414
rect 175509 125411 175575 125414
rect 270361 125411 270427 125414
rect 408870 125036 408930 125550
rect 73246 124732 73252 124796
rect 73316 124732 73322 124796
rect 242025 124794 242091 124797
rect 242158 124794 242164 124796
rect 242025 124792 242164 124794
rect 242025 124736 242030 124792
rect 242086 124736 242164 124792
rect 242025 124734 242164 124736
rect 73254 124660 73314 124732
rect 242025 124731 242091 124734
rect 242158 124732 242164 124734
rect 242228 124732 242234 124796
rect 358313 124794 358379 124797
rect 358497 124794 358563 124797
rect 358313 124792 358563 124794
rect 358313 124736 358318 124792
rect 358374 124736 358502 124792
rect 358558 124736 358563 124792
rect 358313 124734 358563 124736
rect 358313 124731 358379 124734
rect 358497 124731 358563 124734
rect 73246 124596 73252 124660
rect 73316 124596 73322 124660
rect 136961 123298 137027 123301
rect 230985 123298 231051 123301
rect 324733 123298 324799 123301
rect 134710 123296 137027 123298
rect 38797 122754 38863 122757
rect 35534 122752 38863 122754
rect 35534 122696 38802 122752
rect 38858 122696 38863 122752
rect 35534 122694 38863 122696
rect 70678 122754 70738 123268
rect 134710 123240 136966 123296
rect 137022 123240 137027 123296
rect 134710 123238 137027 123240
rect 134710 122928 134770 123238
rect 136961 123235 137027 123238
rect 228734 123296 231051 123298
rect 228734 123240 230990 123296
rect 231046 123240 231051 123296
rect 228734 123238 231051 123240
rect 228734 122928 228794 123238
rect 230985 123235 231051 123238
rect 322758 123296 324799 123298
rect 322758 123240 324738 123296
rect 324794 123240 324799 123296
rect 322758 123238 324799 123240
rect 322758 122928 322818 123238
rect 324733 123235 324799 123238
rect 75413 122754 75479 122757
rect 70678 122752 75479 122754
rect 70678 122696 75418 122752
rect 75474 122696 75479 122752
rect 70678 122694 75479 122696
rect 9896 122618 10376 122648
rect 12669 122618 12735 122621
rect 9896 122616 12735 122618
rect 9896 122560 12674 122616
rect 12730 122560 12735 122616
rect 9896 122558 12735 122560
rect 9896 122528 10376 122558
rect 12669 122555 12735 122558
rect 35534 122520 35594 122694
rect 38797 122691 38863 122694
rect 75413 122691 75479 122694
rect 405969 122618 406035 122621
rect 405969 122616 408930 122618
rect 405969 122560 405974 122616
rect 406030 122560 408930 122616
rect 405969 122558 408930 122560
rect 405969 122555 406035 122558
rect 408870 122452 408930 122558
rect 144229 122346 144295 122349
rect 148686 122346 148692 122348
rect 144229 122344 148692 122346
rect 144229 122288 144234 122344
rect 144290 122288 148692 122344
rect 144229 122286 148692 122288
rect 144229 122283 144295 122286
rect 148686 122284 148692 122286
rect 148756 122284 148762 122348
rect 148870 122148 148876 122212
rect 148940 122148 148946 122212
rect 240369 122210 240435 122213
rect 334209 122210 334275 122213
rect 240369 122208 242932 122210
rect 240369 122152 240374 122208
rect 240430 122152 242932 122208
rect 240369 122150 242932 122152
rect 334209 122208 336956 122210
rect 334209 122152 334214 122208
rect 334270 122152 336956 122208
rect 334209 122150 336956 122152
rect 240369 122147 240435 122150
rect 334209 122147 334275 122150
rect 54069 122074 54135 122077
rect 54662 122074 54668 122076
rect 54069 122072 54668 122074
rect 54069 122016 54074 122072
rect 54130 122016 54668 122072
rect 54069 122014 54668 122016
rect 54069 122011 54135 122014
rect 54662 122012 54668 122014
rect 54732 122074 54738 122076
rect 55030 122074 55036 122076
rect 54732 122014 55036 122074
rect 54732 122012 54738 122014
rect 55030 122012 55036 122014
rect 55100 122012 55106 122076
rect 52597 121258 52663 121261
rect 356197 121258 356263 121261
rect 427497 121258 427563 121261
rect 52597 121256 55068 121258
rect 16165 120714 16231 120717
rect 19894 120714 19954 121228
rect 52597 121200 52602 121256
rect 52658 121200 55068 121256
rect 52597 121198 55068 121200
rect 352780 121256 356263 121258
rect 352780 121200 356202 121256
rect 356258 121200 356263 121256
rect 352780 121198 356263 121200
rect 424724 121256 427563 121258
rect 424724 121200 427502 121256
rect 427558 121200 427563 121256
rect 424724 121198 427563 121200
rect 52597 121195 52663 121198
rect 356197 121195 356263 121198
rect 427497 121195 427563 121198
rect 16165 120712 19954 120714
rect 16165 120656 16170 120712
rect 16226 120656 19954 120712
rect 16165 120654 19954 120656
rect 16165 120651 16231 120654
rect 73389 120578 73455 120581
rect 74217 120578 74283 120581
rect 73389 120576 74283 120578
rect 73389 120520 73394 120576
rect 73450 120520 74222 120576
rect 74278 120520 74283 120576
rect 73389 120518 74283 120520
rect 73389 120515 73455 120518
rect 74217 120515 74283 120518
rect 405969 120578 406035 120581
rect 405969 120576 408930 120578
rect 405969 120520 405974 120576
rect 406030 120520 408930 120576
rect 405969 120518 408930 120520
rect 405969 120515 406035 120518
rect 136869 120442 136935 120445
rect 134710 120440 136935 120442
rect 134710 120384 136874 120440
rect 136930 120384 136935 120440
rect 134710 120382 136935 120384
rect 38797 120306 38863 120309
rect 35718 120304 38863 120306
rect 35718 120248 38802 120304
rect 38858 120248 38863 120304
rect 35718 120246 38863 120248
rect 35718 120072 35778 120246
rect 38797 120243 38863 120246
rect 134710 119800 134770 120382
rect 136869 120379 136935 120382
rect 408870 120004 408930 120518
rect 324549 119898 324615 119901
rect 322758 119896 324615 119898
rect 322758 119840 324554 119896
rect 324610 119840 324615 119896
rect 322758 119838 324615 119840
rect 322758 119800 322818 119838
rect 324549 119835 324615 119838
rect 73389 119762 73455 119765
rect 70862 119760 73455 119762
rect 70862 119704 73394 119760
rect 73450 119704 73455 119760
rect 70862 119702 73455 119704
rect 70862 119596 70922 119702
rect 73389 119699 73455 119702
rect 228734 119354 228794 119796
rect 231854 119354 231860 119356
rect 228734 119294 231860 119354
rect 231854 119292 231860 119294
rect 231924 119292 231930 119356
rect 167873 118810 167939 118813
rect 262357 118810 262423 118813
rect 164732 118808 167939 118810
rect 164732 118752 167878 118808
rect 167934 118752 167939 118808
rect 164732 118750 167939 118752
rect 258756 118808 262423 118810
rect 258756 118752 262362 118808
rect 262418 118752 262423 118808
rect 258756 118750 262423 118752
rect 167873 118747 167939 118750
rect 262357 118747 262423 118750
rect 73798 117660 73804 117724
rect 73868 117722 73874 117724
rect 74350 117722 74356 117724
rect 73868 117662 74356 117722
rect 73868 117660 73874 117662
rect 74350 117660 74356 117662
rect 74420 117660 74426 117724
rect 38245 117586 38311 117589
rect 35748 117584 38311 117586
rect 35748 117528 38250 117584
rect 38306 117528 38311 117584
rect 35748 117526 38311 117528
rect 38245 117523 38311 117526
rect 405969 117450 406035 117453
rect 409054 117450 409114 117556
rect 405969 117448 409114 117450
rect 405969 117392 405974 117448
rect 406030 117392 409114 117448
rect 405969 117390 409114 117392
rect 405969 117387 406035 117390
rect 324549 117314 324615 117317
rect 322758 117312 324615 117314
rect 322758 117256 324554 117312
rect 324610 117256 324615 117312
rect 322758 117254 324615 117256
rect 54069 117178 54135 117181
rect 54846 117178 54852 117180
rect 54069 117176 54852 117178
rect 54069 117120 54074 117176
rect 54130 117120 54852 117176
rect 54069 117118 54852 117120
rect 54069 117115 54135 117118
rect 54846 117116 54852 117118
rect 54916 117116 54922 117180
rect 322758 116672 322818 117254
rect 324549 117251 324615 117254
rect 134710 116634 134770 116668
rect 136910 116634 136916 116636
rect 134710 116574 136916 116634
rect 136910 116572 136916 116574
rect 136980 116572 136986 116636
rect 228734 116634 228794 116668
rect 229278 116634 229284 116636
rect 228734 116574 229284 116634
rect 229278 116572 229284 116574
rect 229348 116634 229354 116636
rect 238846 116634 238852 116636
rect 229348 116574 238852 116634
rect 229348 116572 229354 116574
rect 238846 116572 238852 116574
rect 238916 116572 238922 116636
rect 52137 116226 52203 116229
rect 74125 116226 74191 116229
rect 356197 116226 356263 116229
rect 428693 116226 428759 116229
rect 52137 116224 55068 116226
rect 16257 115138 16323 115141
rect 19894 115138 19954 116196
rect 52137 116168 52142 116224
rect 52198 116168 55068 116224
rect 52137 116166 55068 116168
rect 70862 116224 74191 116226
rect 70862 116168 74130 116224
rect 74186 116168 74191 116224
rect 70862 116166 74191 116168
rect 352780 116224 356263 116226
rect 352780 116168 356202 116224
rect 356258 116168 356263 116224
rect 352780 116166 356263 116168
rect 424724 116224 428759 116226
rect 424724 116168 428698 116224
rect 428754 116168 428759 116224
rect 424724 116166 428759 116168
rect 52137 116163 52203 116166
rect 70862 116060 70922 116166
rect 74125 116163 74191 116166
rect 356197 116163 356263 116166
rect 428693 116163 428759 116166
rect 429429 115274 429495 115277
rect 434416 115274 434896 115304
rect 429429 115272 434896 115274
rect 429429 115216 429434 115272
rect 429490 115216 434896 115272
rect 429429 115214 434896 115216
rect 429429 115211 429495 115214
rect 434416 115184 434896 115214
rect 16257 115136 19954 115138
rect 16257 115080 16262 115136
rect 16318 115080 19954 115136
rect 16257 115078 19954 115080
rect 73481 115138 73547 115141
rect 74125 115138 74191 115141
rect 73481 115136 74191 115138
rect 73481 115080 73486 115136
rect 73542 115080 74130 115136
rect 74186 115080 74191 115136
rect 73481 115078 74191 115080
rect 16257 115075 16323 115078
rect 73481 115075 73547 115078
rect 74125 115075 74191 115078
rect 38797 115002 38863 115005
rect 35748 115000 38863 115002
rect 35748 114944 38802 115000
rect 38858 114944 38863 115000
rect 35748 114942 38863 114944
rect 38797 114939 38863 114942
rect 405969 114866 406035 114869
rect 409054 114866 409114 114972
rect 405969 114864 409114 114866
rect 405969 114808 405974 114864
rect 406030 114808 409114 114864
rect 405969 114806 409114 114808
rect 405969 114803 406035 114806
rect 325469 113642 325535 113645
rect 322758 113640 325535 113642
rect 322758 113584 325474 113640
rect 325530 113584 325535 113640
rect 322758 113582 325535 113584
rect 322758 113544 322818 113582
rect 325469 113579 325535 113582
rect 134710 113234 134770 113540
rect 136869 113234 136935 113237
rect 134710 113232 136935 113234
rect 134710 113176 136874 113232
rect 136930 113176 136935 113232
rect 134710 113174 136935 113176
rect 136869 113171 136935 113174
rect 146621 113236 146687 113237
rect 146621 113232 146668 113236
rect 146732 113234 146738 113236
rect 147766 113234 147772 113236
rect 146621 113176 146626 113232
rect 146621 113172 146668 113176
rect 146732 113174 147772 113234
rect 146732 113172 146738 113174
rect 147766 113172 147772 113174
rect 147836 113172 147842 113236
rect 146621 113171 146687 113172
rect 51861 113098 51927 113101
rect 52638 113098 52644 113100
rect 51861 113096 52644 113098
rect 51861 113040 51866 113096
rect 51922 113040 52644 113096
rect 51861 113038 52644 113040
rect 51861 113035 51927 113038
rect 52638 113036 52644 113038
rect 52708 113036 52714 113100
rect 228734 112962 228794 113540
rect 230750 112962 230756 112964
rect 228734 112902 230756 112962
rect 230750 112900 230756 112902
rect 230820 112900 230826 112964
rect 38797 112826 38863 112829
rect 73573 112826 73639 112829
rect 74534 112826 74540 112828
rect 35534 112824 38863 112826
rect 35534 112768 38802 112824
rect 38858 112768 38863 112824
rect 35534 112766 38863 112768
rect 35534 112592 35594 112766
rect 38797 112763 38863 112766
rect 70862 112824 74540 112826
rect 70862 112768 73578 112824
rect 73634 112768 74540 112824
rect 70862 112766 74540 112768
rect 70862 112388 70922 112766
rect 73573 112763 73639 112766
rect 74534 112764 74540 112766
rect 74604 112764 74610 112828
rect 405969 112690 406035 112693
rect 405969 112688 408930 112690
rect 405969 112632 405974 112688
rect 406030 112632 408930 112688
rect 405969 112630 408930 112632
rect 405969 112627 406035 112630
rect 408870 112524 408930 112630
rect 52597 111330 52663 111333
rect 356197 111330 356263 111333
rect 427589 111330 427655 111333
rect 52597 111328 55068 111330
rect 16349 111058 16415 111061
rect 19894 111058 19954 111300
rect 52597 111272 52602 111328
rect 52658 111272 55068 111328
rect 52597 111270 55068 111272
rect 352780 111328 356263 111330
rect 352780 111272 356202 111328
rect 356258 111272 356263 111328
rect 352780 111270 356263 111272
rect 424724 111328 427655 111330
rect 424724 111272 427594 111328
rect 427650 111272 427655 111328
rect 424724 111270 427655 111272
rect 52597 111267 52663 111270
rect 356197 111267 356263 111270
rect 427589 111267 427655 111270
rect 16349 111056 19954 111058
rect 16349 111000 16354 111056
rect 16410 111000 19954 111056
rect 16349 110998 19954 111000
rect 16349 110995 16415 110998
rect 325377 110922 325443 110925
rect 322758 110920 325443 110922
rect 322758 110864 325382 110920
rect 325438 110864 325443 110920
rect 322758 110862 325443 110864
rect 136869 110786 136935 110789
rect 134710 110784 136935 110786
rect 134710 110728 136874 110784
rect 136930 110728 136935 110784
rect 134710 110726 136935 110728
rect 38245 110514 38311 110517
rect 35718 110512 38311 110514
rect 35718 110456 38250 110512
rect 38306 110456 38311 110512
rect 35718 110454 38311 110456
rect 35718 110144 35778 110454
rect 38245 110451 38311 110454
rect 84705 109836 84771 109837
rect 134710 109836 134770 110726
rect 136869 110723 136935 110726
rect 228734 109970 228794 110412
rect 241974 110180 241980 110244
rect 242044 110242 242050 110244
rect 242526 110242 242532 110244
rect 242044 110182 242532 110242
rect 242044 110180 242050 110182
rect 242526 110180 242532 110182
rect 242596 110180 242602 110244
rect 231997 109970 232063 109973
rect 228734 109968 232063 109970
rect 228734 109912 232002 109968
rect 232058 109912 232063 109968
rect 228734 109910 232063 109912
rect 231997 109907 232063 109910
rect 240093 109836 240159 109837
rect 322758 109836 322818 110862
rect 325377 110859 325443 110862
rect 406061 110650 406127 110653
rect 406061 110648 408930 110650
rect 406061 110592 406066 110648
rect 406122 110592 408930 110648
rect 406061 110590 408930 110592
rect 406061 110587 406127 110590
rect 408870 110076 408930 110590
rect 84654 109834 84660 109836
rect 84614 109774 84660 109834
rect 84724 109832 84771 109836
rect 84766 109776 84771 109832
rect 84654 109772 84660 109774
rect 84724 109772 84771 109776
rect 134702 109772 134708 109836
rect 134772 109772 134778 109836
rect 240093 109834 240140 109836
rect 240048 109832 240140 109834
rect 240048 109776 240098 109832
rect 240048 109774 240140 109776
rect 240093 109772 240140 109774
rect 240204 109772 240210 109836
rect 322750 109772 322756 109836
rect 322820 109772 322826 109836
rect 84705 109771 84771 109772
rect 240093 109771 240159 109772
rect 73665 109562 73731 109565
rect 73798 109562 73804 109564
rect 73665 109560 73804 109562
rect 73665 109504 73670 109560
rect 73726 109504 73804 109560
rect 73665 109502 73804 109504
rect 73665 109499 73731 109502
rect 73798 109500 73804 109502
rect 73868 109500 73874 109564
rect 9896 109154 10376 109184
rect 13405 109154 13471 109157
rect 9896 109152 13471 109154
rect 9896 109096 13410 109152
rect 13466 109096 13471 109152
rect 9896 109094 13471 109096
rect 9896 109064 10376 109094
rect 13405 109091 13471 109094
rect 73665 108882 73731 108885
rect 70862 108880 73731 108882
rect 70862 108824 73670 108880
rect 73726 108824 73731 108880
rect 70862 108822 73731 108824
rect 70862 108716 70922 108822
rect 73665 108819 73731 108822
rect 82589 108882 82655 108885
rect 143953 108882 144019 108885
rect 148686 108882 148692 108884
rect 82589 108880 84538 108882
rect 82589 108824 82594 108880
rect 82650 108824 84538 108880
rect 82589 108822 84538 108824
rect 82589 108819 82655 108822
rect 84478 108814 84538 108822
rect 143953 108880 148692 108882
rect 143953 108824 143958 108880
rect 144014 108824 148692 108880
rect 143953 108822 148692 108824
rect 143953 108819 144019 108822
rect 148686 108820 148692 108822
rect 148756 108820 148762 108884
rect 148870 108820 148876 108884
rect 148940 108820 148946 108884
rect 176245 108882 176311 108885
rect 240829 108882 240895 108885
rect 269993 108882 270059 108885
rect 334209 108882 334275 108885
rect 176245 108880 178378 108882
rect 176245 108824 176250 108880
rect 176306 108824 178378 108880
rect 176245 108822 178378 108824
rect 176245 108819 176311 108822
rect 178318 108814 178378 108822
rect 240829 108880 242932 108882
rect 240829 108824 240834 108880
rect 240890 108824 242932 108880
rect 240829 108822 242932 108824
rect 269993 108880 272402 108882
rect 269993 108824 269998 108880
rect 270054 108824 272402 108880
rect 269993 108822 272402 108824
rect 240829 108819 240895 108822
rect 269993 108819 270059 108822
rect 272342 108814 272402 108822
rect 334209 108880 336956 108882
rect 334209 108824 334214 108880
rect 334270 108824 336956 108880
rect 334209 108822 336956 108824
rect 334209 108819 334275 108822
rect 84478 108754 85060 108814
rect 178318 108754 178900 108814
rect 272342 108754 272924 108814
rect 230801 107932 230867 107933
rect 230750 107930 230756 107932
rect 228734 107870 230756 107930
rect 230820 107930 230867 107932
rect 230820 107928 230948 107930
rect 230862 107872 230948 107928
rect 38797 107522 38863 107525
rect 35748 107520 38863 107522
rect 35748 107464 38802 107520
rect 38858 107464 38863 107520
rect 35748 107462 38863 107464
rect 38797 107459 38863 107462
rect 228734 107288 228794 107870
rect 230750 107868 230756 107870
rect 230820 107870 230948 107872
rect 230820 107868 230867 107870
rect 230801 107867 230867 107868
rect 405969 107658 406035 107661
rect 405969 107656 408930 107658
rect 405969 107600 405974 107656
rect 406030 107600 408930 107656
rect 405969 107598 408930 107600
rect 405969 107595 406035 107598
rect 408870 107492 408930 107598
rect 134710 106842 134770 107284
rect 137462 106842 137468 106844
rect 134710 106782 137468 106842
rect 137462 106780 137468 106782
rect 137532 106780 137538 106844
rect 322758 106842 322818 107288
rect 324590 106842 324596 106844
rect 322758 106782 324596 106842
rect 324590 106780 324596 106782
rect 324660 106780 324666 106844
rect 18097 106298 18163 106301
rect 52597 106298 52663 106301
rect 356197 106298 356263 106301
rect 427589 106298 427655 106301
rect 18097 106296 19924 106298
rect 18097 106240 18102 106296
rect 18158 106240 19924 106296
rect 18097 106238 19924 106240
rect 52597 106296 55068 106298
rect 52597 106240 52602 106296
rect 52658 106240 55068 106296
rect 52597 106238 55068 106240
rect 352780 106296 356263 106298
rect 352780 106240 356202 106296
rect 356258 106240 356263 106296
rect 352780 106238 356263 106240
rect 424724 106296 427655 106298
rect 424724 106240 427594 106296
rect 427650 106240 427655 106296
rect 424724 106238 427655 106240
rect 18097 106235 18163 106238
rect 52597 106235 52663 106238
rect 356197 106235 356263 106238
rect 427589 106235 427655 106238
rect 38797 105346 38863 105349
rect 35534 105344 38863 105346
rect 35534 105288 38802 105344
rect 38858 105288 38863 105344
rect 35534 105286 38863 105288
rect 35534 105112 35594 105286
rect 38797 105283 38863 105286
rect 405969 105346 406035 105349
rect 405969 105344 408930 105346
rect 405969 105288 405974 105344
rect 406030 105288 408930 105344
rect 405969 105286 408930 105288
rect 405969 105283 406035 105286
rect 74033 105210 74099 105213
rect 70862 105208 74099 105210
rect 70862 105152 74038 105208
rect 74094 105152 74099 105208
rect 70862 105150 74099 105152
rect 70862 105044 70922 105150
rect 74033 105147 74099 105150
rect 408870 105044 408930 105286
rect 138014 104394 138020 104396
rect 134710 104334 138020 104394
rect 134710 104160 134770 104334
rect 138014 104332 138020 104334
rect 138084 104332 138090 104396
rect 230709 104394 230775 104397
rect 231854 104394 231860 104396
rect 228734 104392 231860 104394
rect 228734 104336 230714 104392
rect 230770 104336 231860 104392
rect 228734 104334 231860 104336
rect 228734 103988 228794 104334
rect 230709 104331 230775 104334
rect 231854 104332 231860 104334
rect 231924 104332 231930 104396
rect 322758 103988 322818 104160
rect 228726 103924 228732 103988
rect 228796 103924 228802 103988
rect 322750 103924 322756 103988
rect 322820 103924 322826 103988
rect 261110 102972 261116 103036
rect 261180 103034 261186 103036
rect 270494 103034 270500 103036
rect 261180 102974 270500 103034
rect 261180 102972 261186 102974
rect 270494 102972 270500 102974
rect 270564 102972 270570 103036
rect 429429 102762 429495 102765
rect 434416 102762 434896 102792
rect 429429 102760 434896 102762
rect 429429 102704 429434 102760
rect 429490 102704 434896 102760
rect 429429 102702 434896 102704
rect 429429 102699 429495 102702
rect 434416 102672 434896 102702
rect 38613 102490 38679 102493
rect 35748 102488 38679 102490
rect 35748 102432 38618 102488
rect 38674 102432 38679 102488
rect 35748 102430 38679 102432
rect 38613 102427 38679 102430
rect 171318 102292 171324 102356
rect 171388 102354 171394 102356
rect 177022 102354 177028 102356
rect 171388 102294 177028 102354
rect 171388 102292 171394 102294
rect 177022 102292 177028 102294
rect 177092 102292 177098 102356
rect 405969 102218 406035 102221
rect 409054 102218 409114 102460
rect 405969 102216 409114 102218
rect 405969 102160 405974 102216
rect 406030 102160 409114 102216
rect 405969 102158 409114 102160
rect 405969 102155 406035 102158
rect 74166 102082 74172 102084
rect 70862 102022 74172 102082
rect 70862 101508 70922 102022
rect 74166 102020 74172 102022
rect 74236 102020 74242 102084
rect 17453 101266 17519 101269
rect 52597 101266 52663 101269
rect 356197 101266 356263 101269
rect 427405 101266 427471 101269
rect 17453 101264 19924 101266
rect 17453 101208 17458 101264
rect 17514 101208 19924 101264
rect 17453 101206 19924 101208
rect 52597 101264 55068 101266
rect 52597 101208 52602 101264
rect 52658 101208 55068 101264
rect 52597 101206 55068 101208
rect 352780 101264 356263 101266
rect 352780 101208 356202 101264
rect 356258 101208 356263 101264
rect 352780 101206 356263 101208
rect 424724 101264 427471 101266
rect 424724 101208 427410 101264
rect 427466 101208 427471 101264
rect 424724 101206 427471 101208
rect 17453 101203 17519 101206
rect 52597 101203 52663 101206
rect 356197 101203 356263 101206
rect 427405 101203 427471 101206
rect 38797 100314 38863 100317
rect 35718 100312 38863 100314
rect 35718 100256 38802 100312
rect 38858 100256 38863 100312
rect 35718 100254 38863 100256
rect 134710 100314 134770 101028
rect 164878 100660 164884 100724
rect 164948 100722 164954 100724
rect 178678 100722 178684 100724
rect 164948 100662 178684 100722
rect 164948 100660 164954 100662
rect 178678 100660 178684 100662
rect 178748 100660 178754 100724
rect 134710 100254 136978 100314
rect 35718 100080 35778 100254
rect 38797 100251 38863 100254
rect 136918 99906 136978 100254
rect 164929 100042 164995 100045
rect 228734 100044 228794 101028
rect 242025 100724 242091 100725
rect 241974 100660 241980 100724
rect 242044 100722 242091 100724
rect 242044 100720 242136 100722
rect 242086 100664 242136 100720
rect 242044 100662 242136 100664
rect 242044 100660 242091 100662
rect 258718 100660 258724 100724
rect 258788 100722 258794 100724
rect 272702 100722 272708 100724
rect 258788 100662 272708 100722
rect 258788 100660 258794 100662
rect 272702 100660 272708 100662
rect 272772 100660 272778 100724
rect 242025 100659 242091 100660
rect 322758 100452 322818 101032
rect 405969 100586 406035 100589
rect 405969 100584 408930 100586
rect 405969 100528 405974 100584
rect 406030 100528 408930 100584
rect 405969 100526 408930 100528
rect 405969 100523 406035 100526
rect 322750 100388 322756 100452
rect 322820 100388 322826 100452
rect 178678 100042 178684 100044
rect 164929 100040 178684 100042
rect 164929 99984 164934 100040
rect 164990 99984 178684 100040
rect 164929 99982 178684 99984
rect 164929 99979 164995 99982
rect 178678 99980 178684 99982
rect 178748 99980 178754 100044
rect 228726 99980 228732 100044
rect 228796 100042 228802 100044
rect 230893 100042 230959 100045
rect 228796 100040 231922 100042
rect 228796 99984 230898 100040
rect 230954 99984 231922 100040
rect 228796 99982 231922 99984
rect 228796 99980 228802 99982
rect 230893 99979 230959 99982
rect 145742 99906 145748 99908
rect 136918 99846 145748 99906
rect 145742 99844 145748 99846
rect 145812 99844 145818 99908
rect 231862 99906 231922 99982
rect 258718 99980 258724 100044
rect 258788 100042 258794 100044
rect 272702 100042 272708 100044
rect 258788 99982 272708 100042
rect 258788 99980 258794 99982
rect 272702 99980 272708 99982
rect 272772 99980 272778 100044
rect 408870 100012 408930 100526
rect 242710 99906 242716 99908
rect 231862 99846 242716 99906
rect 242710 99844 242716 99846
rect 242780 99844 242786 99908
rect 167873 98818 167939 98821
rect 261161 98818 261227 98821
rect 164732 98816 167939 98818
rect 164732 98760 167878 98816
rect 167934 98760 167939 98816
rect 164732 98758 167939 98760
rect 258756 98816 261227 98818
rect 258756 98760 261166 98816
rect 261222 98760 261227 98816
rect 258756 98758 261227 98760
rect 167873 98755 167939 98758
rect 261161 98755 261227 98758
rect 164929 98684 164995 98685
rect 164878 98682 164884 98684
rect 164838 98622 164884 98682
rect 164948 98680 164995 98684
rect 164990 98624 164995 98680
rect 164878 98620 164884 98622
rect 164948 98620 164995 98624
rect 164929 98619 164995 98620
rect 137513 98546 137579 98549
rect 231353 98546 231419 98549
rect 325193 98546 325259 98549
rect 134710 98544 137579 98546
rect 134710 98488 137518 98544
rect 137574 98488 137579 98544
rect 134710 98486 137579 98488
rect 73614 98274 73620 98276
rect 70862 98214 73620 98274
rect 38797 97866 38863 97869
rect 35534 97864 38863 97866
rect 35534 97808 38802 97864
rect 38858 97808 38863 97864
rect 70862 97836 70922 98214
rect 73614 98212 73620 98214
rect 73684 98212 73690 98276
rect 134710 97904 134770 98486
rect 137513 98483 137579 98486
rect 228734 98544 231419 98546
rect 228734 98488 231358 98544
rect 231414 98488 231419 98544
rect 228734 98486 231419 98488
rect 228734 97904 228794 98486
rect 231353 98483 231419 98486
rect 322758 98544 325259 98546
rect 322758 98488 325198 98544
rect 325254 98488 325259 98544
rect 322758 98486 325259 98488
rect 322758 97904 322818 98486
rect 325193 98483 325259 98486
rect 352793 97868 352859 97869
rect 35534 97806 38863 97808
rect 35534 97632 35594 97806
rect 38797 97803 38863 97806
rect 352742 97804 352748 97868
rect 352812 97866 352859 97868
rect 352812 97864 352904 97866
rect 352854 97808 352904 97864
rect 352812 97806 352904 97808
rect 352812 97804 352859 97806
rect 352793 97803 352859 97804
rect 405969 97730 406035 97733
rect 405969 97728 408930 97730
rect 405969 97672 405974 97728
rect 406030 97672 408930 97728
rect 405969 97670 408930 97672
rect 405969 97667 406035 97670
rect 408870 97564 408930 97670
rect 18097 96234 18163 96237
rect 52597 96234 52663 96237
rect 356197 96234 356263 96237
rect 427221 96234 427287 96237
rect 18097 96232 19924 96234
rect 18097 96176 18102 96232
rect 18158 96176 19924 96232
rect 18097 96174 19924 96176
rect 52597 96232 55068 96234
rect 52597 96176 52602 96232
rect 52658 96176 55068 96232
rect 52597 96174 55068 96176
rect 352780 96232 356263 96234
rect 352780 96176 356202 96232
rect 356258 96176 356263 96232
rect 352780 96174 356263 96176
rect 424724 96232 427287 96234
rect 424724 96176 427226 96232
rect 427282 96176 427287 96232
rect 424724 96174 427287 96176
rect 18097 96171 18163 96174
rect 52597 96171 52663 96174
rect 356197 96171 356263 96174
rect 427221 96171 427287 96174
rect 9896 95826 10376 95856
rect 13129 95826 13195 95829
rect 242025 95828 242091 95829
rect 241974 95826 241980 95828
rect 9896 95824 13195 95826
rect 9896 95768 13134 95824
rect 13190 95768 13195 95824
rect 9896 95766 13195 95768
rect 241934 95766 241980 95826
rect 242044 95824 242091 95828
rect 242086 95768 242091 95824
rect 9896 95736 10376 95766
rect 13129 95763 13195 95766
rect 241974 95764 241980 95766
rect 242044 95764 242091 95768
rect 242025 95763 242091 95764
rect 148870 95492 148876 95556
rect 148940 95492 148946 95556
rect 240369 95554 240435 95557
rect 334209 95554 334275 95557
rect 405969 95554 406035 95557
rect 240369 95552 242932 95554
rect 240369 95496 240374 95552
rect 240430 95496 242932 95552
rect 240369 95494 242932 95496
rect 334209 95552 336956 95554
rect 334209 95496 334214 95552
rect 334270 95496 336956 95552
rect 334209 95494 336956 95496
rect 405969 95552 408930 95554
rect 405969 95496 405974 95552
rect 406030 95496 408930 95552
rect 405969 95494 408930 95496
rect 240369 95491 240435 95494
rect 334209 95491 334275 95494
rect 405969 95491 406035 95494
rect 38061 95418 38127 95421
rect 35718 95416 38127 95418
rect 35718 95360 38066 95416
rect 38122 95360 38127 95416
rect 35718 95358 38127 95360
rect 35718 95048 35778 95358
rect 38061 95355 38127 95358
rect 231997 95010 232063 95013
rect 324549 95010 324615 95013
rect 228734 95008 232063 95010
rect 228734 94952 232002 95008
rect 232058 94952 232063 95008
rect 228734 94950 232063 94952
rect 228734 94776 228794 94950
rect 231997 94947 232063 94950
rect 322758 95008 324615 95010
rect 322758 94952 324554 95008
rect 324610 94952 324615 95008
rect 408870 94980 408930 95494
rect 322758 94950 324615 94952
rect 322758 94776 322818 94950
rect 324549 94947 324615 94950
rect 134710 94602 134770 94772
rect 138157 94602 138223 94605
rect 134710 94600 138223 94602
rect 134710 94544 138162 94600
rect 138218 94544 138223 94600
rect 134710 94542 138223 94544
rect 138157 94539 138223 94542
rect 70678 93922 70738 94164
rect 74534 93922 74540 93924
rect 70678 93862 74540 93922
rect 74534 93860 74540 93862
rect 74604 93860 74610 93924
rect 84654 93452 84660 93516
rect 84724 93514 84730 93516
rect 84797 93514 84863 93517
rect 84724 93512 84863 93514
rect 84724 93456 84802 93512
rect 84858 93456 84863 93512
rect 84724 93454 84863 93456
rect 84724 93452 84730 93454
rect 84797 93451 84863 93454
rect 37601 92562 37667 92565
rect 35748 92560 37667 92562
rect 35748 92504 37606 92560
rect 37662 92504 37667 92560
rect 35748 92502 37667 92504
rect 37601 92499 37667 92502
rect 405969 92426 406035 92429
rect 409054 92426 409114 92532
rect 405969 92424 409114 92426
rect 405969 92368 405974 92424
rect 406030 92368 409114 92424
rect 405969 92366 409114 92368
rect 405969 92363 406035 92366
rect 82681 92290 82747 92293
rect 137605 92290 137671 92293
rect 82681 92288 84538 92290
rect 82681 92232 82686 92288
rect 82742 92232 84538 92288
rect 82681 92230 84538 92232
rect 82681 92227 82747 92230
rect 84478 92222 84538 92230
rect 134710 92288 137671 92290
rect 134710 92232 137610 92288
rect 137666 92232 137671 92288
rect 134710 92230 137671 92232
rect 84478 92162 85060 92222
rect 134710 91648 134770 92230
rect 137605 92227 137671 92230
rect 175509 92290 175575 92293
rect 231445 92290 231511 92293
rect 175509 92288 178378 92290
rect 175509 92232 175514 92288
rect 175570 92232 178378 92288
rect 175509 92230 178378 92232
rect 175509 92227 175575 92230
rect 178318 92222 178378 92230
rect 228734 92288 231511 92290
rect 228734 92232 231450 92288
rect 231506 92232 231511 92288
rect 228734 92230 231511 92232
rect 178318 92162 178900 92222
rect 228734 91648 228794 92230
rect 231445 92227 231511 92230
rect 270361 92290 270427 92293
rect 325285 92290 325351 92293
rect 270361 92288 272402 92290
rect 270361 92232 270366 92288
rect 270422 92232 272402 92288
rect 270361 92230 272402 92232
rect 270361 92227 270427 92230
rect 272342 92222 272402 92230
rect 322758 92288 325351 92290
rect 322758 92232 325290 92288
rect 325346 92232 325351 92288
rect 322758 92230 325351 92232
rect 272342 92162 272924 92222
rect 322758 91648 322818 92230
rect 325285 92227 325351 92230
rect 427589 91610 427655 91613
rect 424694 91608 427655 91610
rect 424694 91552 427594 91608
rect 427650 91552 427655 91608
rect 424694 91550 427655 91552
rect 424694 91376 424754 91550
rect 427589 91547 427655 91550
rect 18097 91338 18163 91341
rect 52597 91338 52663 91341
rect 356197 91338 356263 91341
rect 18097 91336 19924 91338
rect 18097 91280 18102 91336
rect 18158 91280 19924 91336
rect 18097 91278 19924 91280
rect 52597 91336 55068 91338
rect 52597 91280 52602 91336
rect 52658 91280 55068 91336
rect 52597 91278 55068 91280
rect 352780 91336 356263 91338
rect 352780 91280 356202 91336
rect 356258 91280 356263 91336
rect 352780 91278 356263 91280
rect 18097 91275 18163 91278
rect 52597 91275 52663 91278
rect 356197 91275 356263 91278
rect 73389 91202 73455 91205
rect 70862 91200 73455 91202
rect 70862 91144 73394 91200
rect 73450 91144 73455 91200
rect 70862 91142 73455 91144
rect 70862 90628 70922 91142
rect 73389 91139 73455 91142
rect 405969 90250 406035 90253
rect 430165 90250 430231 90253
rect 434416 90250 434896 90280
rect 405969 90248 408930 90250
rect 405969 90192 405974 90248
rect 406030 90192 408930 90248
rect 405969 90190 408930 90192
rect 405969 90187 406035 90190
rect 38797 90114 38863 90117
rect 35748 90112 38863 90114
rect 35748 90056 38802 90112
rect 38858 90056 38863 90112
rect 35748 90054 38863 90056
rect 38797 90051 38863 90054
rect 145793 90114 145859 90117
rect 148870 90114 148876 90116
rect 145793 90112 148876 90114
rect 145793 90056 145798 90112
rect 145854 90056 148876 90112
rect 145793 90054 148876 90056
rect 145793 90051 145859 90054
rect 148870 90052 148876 90054
rect 148940 90052 148946 90116
rect 152182 90052 152188 90116
rect 152252 90114 152258 90116
rect 155494 90114 155500 90116
rect 152252 90054 155500 90114
rect 152252 90052 152258 90054
rect 155494 90052 155500 90054
rect 155564 90052 155570 90116
rect 351638 90052 351644 90116
rect 351708 90114 351714 90116
rect 352793 90114 352859 90117
rect 351708 90112 352859 90114
rect 351708 90056 352798 90112
rect 352854 90056 352859 90112
rect 408870 90084 408930 90190
rect 430165 90248 434896 90250
rect 430165 90192 430170 90248
rect 430226 90192 434896 90248
rect 430165 90190 434896 90192
rect 430165 90187 430231 90190
rect 434416 90160 434896 90190
rect 351708 90054 352859 90056
rect 351708 90052 351714 90054
rect 352793 90051 352859 90054
rect 74033 89842 74099 89845
rect 74166 89842 74172 89844
rect 74033 89840 74172 89842
rect 74033 89784 74038 89840
rect 74094 89784 74172 89840
rect 74033 89782 74172 89784
rect 74033 89779 74099 89782
rect 74166 89780 74172 89782
rect 74236 89780 74242 89844
rect 245838 89100 245844 89164
rect 245908 89162 245914 89164
rect 248925 89162 248991 89165
rect 245908 89160 248991 89162
rect 245908 89104 248930 89160
rect 248986 89104 248991 89160
rect 245908 89102 248991 89104
rect 245908 89100 245914 89102
rect 248925 89099 248991 89102
rect 241974 88964 241980 89028
rect 242044 89026 242050 89028
rect 250213 89026 250279 89029
rect 242044 89024 250279 89026
rect 242044 88968 250218 89024
rect 250274 88968 250279 89024
rect 242044 88966 250279 88968
rect 242044 88964 242050 88966
rect 155453 88892 155519 88893
rect 155729 88892 155795 88893
rect 155453 88888 155500 88892
rect 155564 88890 155570 88892
rect 155453 88832 155458 88888
rect 155453 88828 155500 88832
rect 155564 88830 155610 88890
rect 155564 88828 155570 88830
rect 155678 88828 155684 88892
rect 155748 88890 155795 88892
rect 231537 88890 231603 88893
rect 241982 88892 242042 88964
rect 250213 88963 250279 88966
rect 155748 88888 155840 88890
rect 155790 88832 155840 88888
rect 155748 88830 155840 88832
rect 228734 88888 231603 88890
rect 228734 88832 231542 88888
rect 231598 88832 231603 88888
rect 228734 88830 231603 88832
rect 155748 88828 155795 88830
rect 155453 88827 155519 88828
rect 155729 88827 155795 88828
rect 137697 88754 137763 88757
rect 134710 88752 137763 88754
rect 134710 88696 137702 88752
rect 137758 88696 137763 88752
rect 134710 88694 137763 88696
rect 134710 88520 134770 88694
rect 137697 88691 137763 88694
rect 228734 88520 228794 88830
rect 231537 88827 231603 88830
rect 241974 88828 241980 88892
rect 242044 88828 242050 88892
rect 249518 88828 249524 88892
rect 249588 88890 249594 88892
rect 249661 88890 249727 88893
rect 325377 88890 325443 88893
rect 249588 88888 249727 88890
rect 249588 88832 249666 88888
rect 249722 88832 249727 88888
rect 249588 88830 249727 88832
rect 249588 88828 249594 88830
rect 249661 88827 249727 88830
rect 322758 88888 325443 88890
rect 322758 88832 325382 88888
rect 325438 88832 325443 88888
rect 322758 88830 325443 88832
rect 251731 88620 251797 88621
rect 251726 88618 251732 88620
rect 251640 88558 251732 88618
rect 251726 88556 251732 88558
rect 251796 88556 251802 88620
rect 251731 88555 251797 88556
rect 322758 88520 322818 88830
rect 325377 88827 325443 88830
rect 72009 87530 72075 87533
rect 74166 87530 74172 87532
rect 72009 87528 74172 87530
rect 72009 87472 72014 87528
rect 72070 87472 74172 87528
rect 72009 87470 74172 87472
rect 72009 87467 72075 87470
rect 74166 87468 74172 87470
rect 74236 87468 74242 87532
rect 156097 87530 156163 87533
rect 156097 87528 156298 87530
rect 156097 87472 156102 87528
rect 156158 87472 156298 87528
rect 156097 87470 156298 87472
rect 156097 87467 156163 87470
rect 155269 87394 155335 87397
rect 156046 87394 156052 87396
rect 155269 87392 156052 87394
rect 155269 87336 155274 87392
rect 155330 87336 156052 87392
rect 155269 87334 156052 87336
rect 155269 87331 155335 87334
rect 156046 87332 156052 87334
rect 156116 87332 156122 87396
rect 156238 87394 156298 87470
rect 246206 87468 246212 87532
rect 246276 87530 246282 87532
rect 246276 87470 250506 87530
rect 246276 87468 246282 87470
rect 167638 87394 167644 87396
rect 156238 87334 167644 87394
rect 167638 87332 167644 87334
rect 167708 87332 167714 87396
rect 250446 87394 250506 87470
rect 251174 87394 251180 87396
rect 250446 87334 251180 87394
rect 251174 87332 251180 87334
rect 251244 87332 251250 87396
rect 148502 87196 148508 87260
rect 148572 87258 148578 87260
rect 157753 87258 157819 87261
rect 148572 87256 157819 87258
rect 148572 87200 157758 87256
rect 157814 87200 157819 87256
rect 148572 87198 157819 87200
rect 148572 87196 148578 87198
rect 157753 87195 157819 87198
rect 159041 87122 159107 87125
rect 168742 87122 168748 87124
rect 159041 87120 168748 87122
rect 159041 87064 159046 87120
rect 159102 87064 168748 87120
rect 159041 87062 168748 87064
rect 159041 87059 159107 87062
rect 168742 87060 168748 87062
rect 168812 87060 168818 87124
rect 158397 86986 158463 86989
rect 169294 86986 169300 86988
rect 158397 86984 169300 86986
rect 158397 86928 158402 86984
rect 158458 86928 169300 86984
rect 158397 86926 169300 86928
rect 158397 86923 158463 86926
rect 169294 86924 169300 86926
rect 169364 86924 169370 86988
rect 156557 86850 156623 86853
rect 168006 86850 168012 86852
rect 156557 86848 168012 86850
rect 156557 86792 156562 86848
rect 156618 86792 168012 86848
rect 156557 86790 168012 86792
rect 156557 86787 156623 86790
rect 168006 86788 168012 86790
rect 168076 86788 168082 86852
rect 253341 86850 253407 86853
rect 262398 86850 262404 86852
rect 253341 86848 262404 86850
rect 253341 86792 253346 86848
rect 253402 86792 262404 86848
rect 253341 86790 262404 86792
rect 253341 86787 253407 86790
rect 262398 86788 262404 86790
rect 262468 86788 262474 86852
rect 157201 86714 157267 86717
rect 169110 86714 169116 86716
rect 157201 86712 169116 86714
rect 157201 86656 157206 86712
rect 157262 86656 169116 86712
rect 157201 86654 169116 86656
rect 157201 86651 157267 86654
rect 169110 86652 169116 86654
rect 169180 86652 169186 86716
rect 251317 86714 251383 86717
rect 262582 86714 262588 86716
rect 251317 86712 262588 86714
rect 251317 86656 251322 86712
rect 251378 86656 262588 86712
rect 251317 86654 262588 86656
rect 251317 86651 251383 86654
rect 262582 86652 262588 86654
rect 262652 86652 262658 86716
rect 326573 86714 326639 86717
rect 336366 86714 336372 86716
rect 326573 86712 336372 86714
rect 326573 86656 326578 86712
rect 326634 86656 336372 86712
rect 326573 86654 336372 86656
rect 326573 86651 326639 86654
rect 336366 86652 336372 86654
rect 336436 86714 336442 86716
rect 412869 86714 412935 86717
rect 336436 86712 412935 86714
rect 336436 86656 412874 86712
rect 412930 86656 412935 86712
rect 336436 86654 412935 86656
rect 336436 86652 336442 86654
rect 412869 86651 412935 86654
rect 73849 86442 73915 86445
rect 74534 86442 74540 86444
rect 73849 86440 74540 86442
rect 73849 86384 73854 86440
rect 73910 86384 74540 86440
rect 73849 86382 74540 86384
rect 73849 86379 73915 86382
rect 74534 86380 74540 86382
rect 74604 86380 74610 86444
rect 72878 86244 72884 86308
rect 72948 86306 72954 86308
rect 73573 86306 73639 86309
rect 72948 86304 73639 86306
rect 72948 86248 73578 86304
rect 73634 86248 73639 86304
rect 72948 86246 73639 86248
rect 72948 86244 72954 86246
rect 73573 86243 73639 86246
rect 251174 86244 251180 86308
rect 251244 86306 251250 86308
rect 252053 86306 252119 86309
rect 251244 86304 252119 86306
rect 251244 86248 252058 86304
rect 252114 86248 252119 86304
rect 251244 86246 252119 86248
rect 251244 86244 251250 86246
rect 252053 86243 252119 86246
rect 72694 86108 72700 86172
rect 72764 86170 72770 86172
rect 73481 86170 73547 86173
rect 72764 86168 73547 86170
rect 72764 86112 73486 86168
rect 73542 86112 73547 86168
rect 72764 86110 73547 86112
rect 72764 86108 72770 86110
rect 73481 86107 73547 86110
rect 73665 86170 73731 86173
rect 73982 86170 73988 86172
rect 73665 86168 73988 86170
rect 73665 86112 73670 86168
rect 73726 86112 73988 86168
rect 73665 86110 73988 86112
rect 73665 86107 73731 86110
rect 73982 86108 73988 86110
rect 74052 86108 74058 86172
rect 249569 86170 249635 86173
rect 249886 86170 249892 86172
rect 249569 86168 249892 86170
rect 249569 86112 249574 86168
rect 249630 86112 249892 86168
rect 249569 86110 249892 86112
rect 249569 86107 249635 86110
rect 249886 86108 249892 86110
rect 249956 86108 249962 86172
rect 137881 85762 137947 85765
rect 231077 85762 231143 85765
rect 324549 85762 324615 85765
rect 134710 85760 137947 85762
rect 134710 85704 137886 85760
rect 137942 85704 137947 85760
rect 134710 85702 137947 85704
rect 134710 85392 134770 85702
rect 137881 85699 137947 85702
rect 228734 85760 231143 85762
rect 228734 85704 231082 85760
rect 231138 85704 231143 85760
rect 228734 85702 231143 85704
rect 228734 85392 228794 85702
rect 231077 85699 231143 85702
rect 322758 85760 324615 85762
rect 322758 85704 324554 85760
rect 324610 85704 324615 85760
rect 322758 85702 324615 85704
rect 322758 85392 322818 85702
rect 324549 85699 324615 85702
rect 178729 84268 178795 84269
rect 178678 84266 178684 84268
rect 178602 84206 178684 84266
rect 178748 84266 178795 84268
rect 182317 84266 182383 84269
rect 178748 84264 182383 84266
rect 178790 84208 182322 84264
rect 182378 84208 182383 84264
rect 178678 84204 178684 84206
rect 178748 84206 182383 84208
rect 178748 84204 178795 84206
rect 178729 84203 178795 84204
rect 182317 84203 182383 84206
rect 242158 83388 242164 83452
rect 242228 83450 242234 83452
rect 242894 83450 242900 83452
rect 242228 83390 242900 83450
rect 242228 83388 242234 83390
rect 242894 83388 242900 83390
rect 242964 83388 242970 83452
rect 9896 82362 10376 82392
rect 13497 82362 13563 82365
rect 9896 82360 13563 82362
rect 9896 82304 13502 82360
rect 13558 82304 13563 82360
rect 9896 82302 13563 82304
rect 9896 82272 10376 82302
rect 13497 82299 13563 82302
rect 54069 78010 54135 78013
rect 54846 78010 54852 78012
rect 54069 78008 54852 78010
rect 54069 77952 54074 78008
rect 54130 77952 54852 78008
rect 54069 77950 54852 77952
rect 54069 77947 54135 77950
rect 54846 77948 54852 77950
rect 54916 77948 54922 78012
rect 52638 77812 52644 77876
rect 52708 77874 52714 77876
rect 53057 77874 53123 77877
rect 52708 77872 53123 77874
rect 52708 77816 53062 77872
rect 53118 77816 53123 77872
rect 52708 77814 53123 77816
rect 52708 77812 52714 77814
rect 53057 77811 53123 77814
rect 54662 77812 54668 77876
rect 54732 77874 54738 77876
rect 55081 77874 55147 77877
rect 54732 77872 55147 77874
rect 54732 77816 55086 77872
rect 55142 77816 55147 77872
rect 54732 77814 55147 77816
rect 54732 77812 54738 77814
rect 55081 77811 55147 77814
rect 55398 77812 55404 77876
rect 55468 77874 55474 77876
rect 56093 77874 56159 77877
rect 55468 77872 56159 77874
rect 55468 77816 56098 77872
rect 56154 77816 56159 77872
rect 55468 77814 56159 77816
rect 55468 77812 55474 77814
rect 56093 77811 56159 77814
rect 350953 77874 351019 77877
rect 351638 77874 351644 77876
rect 350953 77872 351644 77874
rect 350953 77816 350958 77872
rect 351014 77816 351644 77872
rect 350953 77814 351644 77816
rect 350953 77811 351019 77814
rect 351638 77812 351644 77814
rect 351708 77812 351714 77876
rect 351822 77812 351828 77876
rect 351892 77874 351898 77876
rect 352057 77874 352123 77877
rect 351892 77872 352123 77874
rect 351892 77816 352062 77872
rect 352118 77816 352123 77872
rect 351892 77814 352123 77816
rect 351892 77812 351898 77814
rect 352057 77811 352123 77814
rect 429521 77738 429587 77741
rect 434416 77738 434896 77768
rect 429521 77736 434896 77738
rect 429521 77680 429526 77736
rect 429582 77680 434896 77736
rect 429521 77678 434896 77680
rect 429521 77675 429587 77678
rect 434416 77648 434896 77678
rect 79461 75834 79527 75837
rect 76198 75832 79527 75834
rect 76198 75776 79466 75832
rect 79522 75776 79527 75832
rect 76198 75774 79527 75776
rect 76198 75260 76258 75774
rect 79461 75771 79527 75774
rect 238662 75364 238668 75428
rect 238732 75426 238738 75428
rect 242894 75426 242900 75428
rect 238732 75366 242900 75426
rect 238732 75364 238738 75366
rect 242894 75364 242900 75366
rect 242964 75364 242970 75428
rect 251174 75364 251180 75428
rect 251244 75426 251250 75428
rect 261846 75426 261852 75428
rect 251244 75366 261852 75426
rect 251244 75364 251250 75366
rect 261846 75364 261852 75366
rect 261916 75364 261922 75428
rect 139629 75290 139695 75293
rect 173853 75290 173919 75293
rect 139629 75288 143020 75290
rect 139629 75232 139634 75288
rect 139690 75232 143020 75288
rect 139629 75230 143020 75232
rect 170804 75288 173919 75290
rect 170804 75232 173858 75288
rect 173914 75232 173919 75288
rect 170804 75230 173919 75232
rect 139629 75227 139695 75230
rect 173853 75227 173919 75230
rect 233469 75290 233535 75293
rect 266589 75290 266655 75293
rect 233469 75288 237044 75290
rect 233469 75232 233474 75288
rect 233530 75232 237044 75288
rect 233469 75230 237044 75232
rect 264828 75288 266655 75290
rect 264828 75232 266594 75288
rect 266650 75232 266655 75288
rect 264828 75230 266655 75232
rect 233469 75227 233535 75230
rect 266589 75227 266655 75230
rect 328413 75290 328479 75293
rect 328413 75288 331068 75290
rect 328413 75232 328418 75288
rect 328474 75232 331068 75288
rect 328413 75230 331068 75232
rect 328413 75227 328479 75230
rect 174037 74202 174103 74205
rect 266589 74202 266655 74205
rect 170804 74200 174103 74202
rect 76382 73930 76442 74172
rect 170804 74144 174042 74200
rect 174098 74144 174103 74200
rect 170804 74142 174103 74144
rect 264828 74200 266655 74202
rect 264828 74144 266594 74200
rect 266650 74144 266655 74200
rect 264828 74142 266655 74144
rect 174037 74139 174103 74142
rect 266589 74139 266655 74142
rect 328321 74202 328387 74205
rect 328321 74200 331068 74202
rect 328321 74144 328326 74200
rect 328382 74144 331068 74200
rect 328321 74142 331068 74144
rect 328321 74139 328387 74142
rect 80197 73930 80263 73933
rect 76382 73928 80263 73930
rect 76382 73872 80202 73928
rect 80258 73872 80263 73928
rect 76382 73870 80263 73872
rect 80197 73867 80263 73870
rect 139721 73794 139787 73797
rect 142990 73794 143050 74104
rect 139721 73792 143050 73794
rect 139721 73736 139726 73792
rect 139782 73736 143050 73792
rect 139721 73734 143050 73736
rect 233469 73794 233535 73797
rect 237014 73794 237074 74104
rect 233469 73792 237074 73794
rect 233469 73736 233474 73792
rect 233530 73736 237074 73792
rect 233469 73734 237074 73736
rect 139721 73731 139787 73734
rect 233469 73731 233535 73734
rect 172933 73250 172999 73253
rect 266589 73250 266655 73253
rect 170804 73248 172999 73250
rect 76382 72842 76442 73220
rect 170804 73192 172938 73248
rect 172994 73192 172999 73248
rect 170804 73190 172999 73192
rect 264828 73248 266655 73250
rect 264828 73192 266594 73248
rect 266650 73192 266655 73248
rect 264828 73190 266655 73192
rect 172933 73187 172999 73190
rect 266589 73187 266655 73190
rect 79829 72842 79895 72845
rect 76382 72840 79895 72842
rect 76382 72784 79834 72840
rect 79890 72784 79895 72840
rect 76382 72782 79895 72784
rect 79829 72779 79895 72782
rect 139537 72570 139603 72573
rect 142990 72570 143050 73152
rect 139537 72568 143050 72570
rect 139537 72512 139542 72568
rect 139598 72512 143050 72568
rect 139537 72510 143050 72512
rect 233469 72570 233535 72573
rect 237014 72570 237074 73152
rect 233469 72568 237074 72570
rect 233469 72512 233474 72568
rect 233530 72512 237074 72568
rect 233469 72510 237074 72512
rect 327217 72570 327283 72573
rect 331038 72570 331098 73152
rect 327217 72568 331098 72570
rect 327217 72512 327222 72568
rect 327278 72512 331098 72568
rect 327217 72510 331098 72512
rect 139537 72507 139603 72510
rect 233469 72507 233535 72510
rect 327217 72507 327283 72510
rect 173301 72162 173367 72165
rect 266681 72162 266747 72165
rect 170804 72160 173367 72162
rect 76382 71618 76442 72132
rect 170804 72104 173306 72160
rect 173362 72104 173367 72160
rect 170804 72102 173367 72104
rect 264828 72160 266747 72162
rect 264828 72104 266686 72160
rect 266742 72104 266747 72160
rect 264828 72102 266747 72104
rect 173301 72099 173367 72102
rect 266681 72099 266747 72102
rect 78909 71618 78975 71621
rect 76382 71616 78975 71618
rect 76382 71560 78914 71616
rect 78970 71560 78975 71616
rect 76382 71558 78975 71560
rect 78909 71555 78975 71558
rect 139905 71482 139971 71485
rect 142990 71482 143050 72064
rect 139905 71480 143050 71482
rect 139905 71424 139910 71480
rect 139966 71424 143050 71480
rect 139905 71422 143050 71424
rect 233469 71482 233535 71485
rect 237014 71482 237074 72064
rect 233469 71480 237074 71482
rect 233469 71424 233474 71480
rect 233530 71424 237074 71480
rect 233469 71422 237074 71424
rect 327033 71482 327099 71485
rect 331038 71482 331098 72064
rect 327033 71480 331098 71482
rect 327033 71424 327038 71480
rect 327094 71424 331098 71480
rect 327033 71422 331098 71424
rect 139905 71419 139971 71422
rect 233469 71419 233535 71422
rect 327033 71419 327099 71422
rect 80197 71210 80263 71213
rect 76198 71208 80263 71210
rect 76198 71152 80202 71208
rect 80258 71152 80263 71208
rect 76198 71150 80263 71152
rect 76198 71044 76258 71150
rect 80197 71147 80263 71150
rect 139629 71074 139695 71077
rect 174037 71074 174103 71077
rect 139629 71072 143020 71074
rect 139629 71016 139634 71072
rect 139690 71016 143020 71072
rect 139629 71014 143020 71016
rect 170804 71072 174103 71074
rect 170804 71016 174042 71072
rect 174098 71016 174103 71072
rect 170804 71014 174103 71016
rect 139629 71011 139695 71014
rect 174037 71011 174103 71014
rect 233561 71074 233627 71077
rect 266589 71074 266655 71077
rect 233561 71072 237044 71074
rect 233561 71016 233566 71072
rect 233622 71016 237044 71072
rect 233561 71014 237044 71016
rect 264828 71072 266655 71074
rect 264828 71016 266594 71072
rect 266650 71016 266655 71072
rect 264828 71014 266655 71016
rect 233561 71011 233627 71014
rect 266589 71011 266655 71014
rect 328505 71074 328571 71077
rect 328505 71072 331068 71074
rect 328505 71016 328510 71072
rect 328566 71016 331068 71072
rect 328505 71014 331068 71016
rect 328505 71011 328571 71014
rect 174037 70122 174103 70125
rect 266589 70122 266655 70125
rect 170804 70120 174103 70122
rect 76382 69850 76442 70092
rect 170804 70064 174042 70120
rect 174098 70064 174103 70120
rect 170804 70062 174103 70064
rect 264828 70120 266655 70122
rect 264828 70064 266594 70120
rect 266650 70064 266655 70120
rect 264828 70062 266655 70064
rect 174037 70059 174103 70062
rect 266589 70059 266655 70062
rect 80197 69850 80263 69853
rect 76382 69848 80263 69850
rect 76382 69792 80202 69848
rect 80258 69792 80263 69848
rect 76382 69790 80263 69792
rect 80197 69787 80263 69790
rect 139813 69578 139879 69581
rect 142990 69578 143050 70024
rect 139813 69576 143050 69578
rect 139813 69520 139818 69576
rect 139874 69520 143050 69576
rect 139813 69518 143050 69520
rect 233561 69578 233627 69581
rect 237014 69578 237074 70024
rect 233561 69576 237074 69578
rect 233561 69520 233566 69576
rect 233622 69520 237074 69576
rect 233561 69518 237074 69520
rect 327125 69578 327191 69581
rect 331038 69578 331098 70024
rect 327125 69576 331098 69578
rect 327125 69520 327130 69576
rect 327186 69520 331098 69576
rect 327125 69518 331098 69520
rect 139813 69515 139879 69518
rect 233561 69515 233627 69518
rect 327125 69515 327191 69518
rect 87925 69442 87991 69445
rect 131349 69442 131415 69445
rect 87925 69440 90028 69442
rect 87925 69384 87930 69440
rect 87986 69384 90028 69440
rect 87925 69382 90028 69384
rect 129772 69440 131415 69442
rect 129772 69384 131354 69440
rect 131410 69384 131415 69440
rect 129772 69382 131415 69384
rect 87925 69379 87991 69382
rect 131349 69379 131415 69382
rect 181029 69442 181095 69445
rect 226477 69442 226543 69445
rect 181029 69440 184052 69442
rect 181029 69384 181034 69440
rect 181090 69384 184052 69440
rect 181029 69382 184052 69384
rect 223796 69440 226543 69442
rect 223796 69384 226482 69440
rect 226538 69384 226543 69440
rect 223796 69382 226543 69384
rect 181029 69379 181095 69382
rect 226477 69379 226543 69382
rect 274869 69442 274935 69445
rect 321697 69442 321763 69445
rect 274869 69440 278076 69442
rect 274869 69384 274874 69440
rect 274930 69384 278076 69440
rect 274869 69382 278076 69384
rect 317820 69440 321763 69442
rect 317820 69384 321702 69440
rect 321758 69384 321763 69440
rect 317820 69382 321763 69384
rect 274869 69379 274935 69382
rect 321697 69379 321763 69382
rect 9896 69034 10376 69064
rect 13313 69034 13379 69037
rect 172933 69034 172999 69037
rect 266589 69034 266655 69037
rect 9896 69032 13379 69034
rect 9896 68976 13318 69032
rect 13374 68976 13379 69032
rect 170804 69032 172999 69034
rect 9896 68974 13379 68976
rect 9896 68944 10376 68974
rect 13313 68971 13379 68974
rect 76382 68626 76442 69004
rect 170804 68976 172938 69032
rect 172994 68976 172999 69032
rect 170804 68974 172999 68976
rect 264828 69032 266655 69034
rect 264828 68976 266594 69032
rect 266650 68976 266655 69032
rect 264828 68974 266655 68976
rect 172933 68971 172999 68974
rect 266589 68971 266655 68974
rect 79277 68626 79343 68629
rect 76382 68624 79343 68626
rect 76382 68568 79282 68624
rect 79338 68568 79343 68624
rect 76382 68566 79343 68568
rect 79277 68563 79343 68566
rect 87649 68490 87715 68493
rect 131809 68490 131875 68493
rect 87649 68488 90028 68490
rect 87649 68432 87654 68488
rect 87710 68432 90028 68488
rect 87649 68430 90028 68432
rect 129772 68488 131875 68490
rect 129772 68432 131814 68488
rect 131870 68432 131875 68488
rect 129772 68430 131875 68432
rect 87649 68427 87715 68430
rect 131809 68427 131875 68430
rect 139629 68354 139695 68357
rect 142990 68354 143050 68936
rect 180937 68490 181003 68493
rect 225925 68490 225991 68493
rect 180937 68488 184052 68490
rect 180937 68432 180942 68488
rect 180998 68432 184052 68488
rect 180937 68430 184052 68432
rect 223796 68488 225991 68490
rect 223796 68432 225930 68488
rect 225986 68432 225991 68488
rect 223796 68430 225991 68432
rect 180937 68427 181003 68430
rect 225925 68427 225991 68430
rect 139629 68352 143050 68354
rect 139629 68296 139634 68352
rect 139690 68296 143050 68352
rect 139629 68294 143050 68296
rect 233653 68354 233719 68357
rect 237014 68354 237074 68936
rect 274685 68490 274751 68493
rect 321605 68490 321671 68493
rect 274685 68488 278076 68490
rect 274685 68432 274690 68488
rect 274746 68432 278076 68488
rect 274685 68430 278076 68432
rect 317820 68488 321671 68490
rect 317820 68432 321610 68488
rect 321666 68432 321671 68488
rect 317820 68430 321671 68432
rect 274685 68427 274751 68430
rect 321605 68427 321671 68430
rect 233653 68352 237074 68354
rect 233653 68296 233658 68352
rect 233714 68296 237074 68352
rect 233653 68294 237074 68296
rect 327217 68354 327283 68357
rect 331038 68354 331098 68936
rect 327217 68352 331098 68354
rect 327217 68296 327222 68352
rect 327278 68296 331098 68352
rect 327217 68294 331098 68296
rect 139629 68291 139695 68294
rect 233653 68291 233719 68294
rect 327217 68291 327283 68294
rect 173853 67946 173919 67949
rect 266681 67946 266747 67949
rect 170804 67944 173919 67946
rect 76382 67402 76442 67916
rect 170804 67888 173858 67944
rect 173914 67888 173919 67944
rect 170804 67886 173919 67888
rect 264828 67944 266747 67946
rect 264828 67888 266686 67944
rect 266742 67888 266747 67944
rect 264828 67886 266747 67888
rect 173853 67883 173919 67886
rect 266681 67883 266747 67886
rect 87833 67674 87899 67677
rect 132361 67674 132427 67677
rect 87833 67672 90028 67674
rect 87833 67616 87838 67672
rect 87894 67616 90028 67672
rect 87833 67614 90028 67616
rect 129772 67672 132427 67674
rect 129772 67616 132366 67672
rect 132422 67616 132427 67672
rect 129772 67614 132427 67616
rect 87833 67611 87899 67614
rect 132361 67611 132427 67614
rect 80197 67402 80263 67405
rect 76382 67400 80263 67402
rect 76382 67344 80202 67400
rect 80258 67344 80263 67400
rect 76382 67342 80263 67344
rect 80197 67339 80263 67342
rect 139721 67402 139787 67405
rect 142990 67402 143050 67848
rect 181397 67674 181463 67677
rect 226293 67674 226359 67677
rect 181397 67672 184052 67674
rect 181397 67616 181402 67672
rect 181458 67616 184052 67672
rect 181397 67614 184052 67616
rect 223796 67672 226359 67674
rect 223796 67616 226298 67672
rect 226354 67616 226359 67672
rect 223796 67614 226359 67616
rect 181397 67611 181463 67614
rect 226293 67611 226359 67614
rect 139721 67400 143050 67402
rect 139721 67344 139726 67400
rect 139782 67344 143050 67400
rect 139721 67342 143050 67344
rect 139721 67339 139787 67342
rect 233469 67266 233535 67269
rect 237014 67266 237074 67848
rect 274777 67674 274843 67677
rect 321605 67674 321671 67677
rect 274777 67672 278076 67674
rect 274777 67616 274782 67672
rect 274838 67616 278076 67672
rect 274777 67614 278076 67616
rect 317820 67672 321671 67674
rect 317820 67616 321610 67672
rect 321666 67616 321671 67672
rect 317820 67614 321671 67616
rect 274777 67611 274843 67614
rect 321605 67611 321671 67614
rect 233469 67264 237074 67266
rect 233469 67208 233474 67264
rect 233530 67208 237074 67264
rect 233469 67206 237074 67208
rect 328229 67266 328295 67269
rect 331038 67266 331098 67848
rect 328229 67264 331098 67266
rect 328229 67208 328234 67264
rect 328290 67208 331098 67264
rect 328229 67206 331098 67208
rect 233469 67203 233535 67206
rect 328229 67203 328295 67206
rect 139629 67130 139695 67133
rect 139629 67128 142314 67130
rect 139629 67072 139634 67128
rect 139690 67072 142314 67128
rect 139629 67070 142314 67072
rect 139629 67067 139695 67070
rect 76382 66858 76442 66964
rect 142254 66926 142314 67070
rect 174037 66994 174103 66997
rect 170804 66992 174103 66994
rect 170804 66936 174042 66992
rect 174098 66936 174103 66992
rect 170804 66934 174103 66936
rect 174037 66931 174103 66934
rect 234205 66994 234271 66997
rect 266589 66994 266655 66997
rect 234205 66992 237044 66994
rect 234205 66936 234210 66992
rect 234266 66936 237044 66992
rect 234205 66934 237044 66936
rect 264828 66992 266655 66994
rect 264828 66936 266594 66992
rect 266650 66936 266655 66992
rect 264828 66934 266655 66936
rect 234205 66931 234271 66934
rect 266589 66931 266655 66934
rect 326941 66994 327007 66997
rect 326941 66992 331068 66994
rect 326941 66936 326946 66992
rect 327002 66936 331068 66992
rect 326941 66934 331068 66936
rect 326941 66931 327007 66934
rect 142254 66866 143020 66926
rect 80197 66858 80263 66861
rect 76382 66856 80263 66858
rect 76382 66800 80202 66856
rect 80258 66800 80263 66856
rect 76382 66798 80263 66800
rect 80197 66795 80263 66798
rect 87189 66722 87255 66725
rect 132545 66722 132611 66725
rect 226293 66722 226359 66725
rect 87189 66720 90028 66722
rect 87189 66664 87194 66720
rect 87250 66664 90028 66720
rect 87189 66662 90028 66664
rect 129772 66720 132611 66722
rect 129772 66664 132550 66720
rect 132606 66664 132611 66720
rect 129772 66662 132611 66664
rect 223796 66720 226359 66722
rect 223796 66664 226298 66720
rect 226354 66664 226359 66720
rect 223796 66662 226359 66664
rect 87189 66659 87255 66662
rect 132545 66659 132611 66662
rect 226293 66659 226359 66662
rect 274869 66722 274935 66725
rect 321237 66722 321303 66725
rect 274869 66720 278076 66722
rect 274869 66664 274874 66720
rect 274930 66664 278076 66720
rect 274869 66662 278076 66664
rect 317820 66720 321303 66722
rect 317820 66664 321242 66720
rect 321298 66664 321303 66720
rect 317820 66662 321303 66664
rect 274869 66659 274935 66662
rect 321237 66659 321303 66662
rect 181949 66450 182015 66453
rect 184022 66450 184082 66624
rect 181949 66448 184082 66450
rect 181949 66392 181954 66448
rect 182010 66392 184082 66448
rect 181949 66390 184082 66392
rect 181949 66387 182015 66390
rect 87281 65906 87347 65909
rect 132361 65906 132427 65909
rect 173853 65906 173919 65909
rect 87281 65904 90028 65906
rect 76382 65634 76442 65876
rect 87281 65848 87286 65904
rect 87342 65848 90028 65904
rect 87281 65846 90028 65848
rect 129772 65904 132427 65906
rect 129772 65848 132366 65904
rect 132422 65848 132427 65904
rect 129772 65846 132427 65848
rect 170804 65904 173919 65906
rect 170804 65848 173858 65904
rect 173914 65848 173919 65904
rect 170804 65846 173919 65848
rect 87281 65843 87347 65846
rect 132361 65843 132427 65846
rect 173853 65843 173919 65846
rect 182133 65906 182199 65909
rect 226385 65906 226451 65909
rect 266589 65906 266655 65909
rect 182133 65904 184052 65906
rect 182133 65848 182138 65904
rect 182194 65848 184052 65904
rect 182133 65846 184052 65848
rect 223796 65904 226451 65906
rect 223796 65848 226390 65904
rect 226446 65848 226451 65904
rect 223796 65846 226451 65848
rect 264828 65904 266655 65906
rect 264828 65848 266594 65904
rect 266650 65848 266655 65904
rect 264828 65846 266655 65848
rect 182133 65843 182199 65846
rect 226385 65843 226451 65846
rect 266589 65843 266655 65846
rect 274961 65906 275027 65909
rect 321605 65906 321671 65909
rect 274961 65904 278076 65906
rect 274961 65848 274966 65904
rect 275022 65848 278076 65904
rect 274961 65846 278076 65848
rect 317820 65904 321671 65906
rect 317820 65848 321610 65904
rect 321666 65848 321671 65904
rect 317820 65846 321671 65848
rect 274961 65843 275027 65846
rect 321605 65843 321671 65846
rect 80197 65634 80263 65637
rect 76382 65632 80263 65634
rect 76382 65576 80202 65632
rect 80258 65576 80263 65632
rect 76382 65574 80263 65576
rect 80197 65571 80263 65574
rect 139905 65498 139971 65501
rect 142990 65498 143050 65808
rect 139905 65496 143050 65498
rect 139905 65440 139910 65496
rect 139966 65440 143050 65496
rect 139905 65438 143050 65440
rect 234389 65498 234455 65501
rect 237014 65498 237074 65808
rect 234389 65496 237074 65498
rect 234389 65440 234394 65496
rect 234450 65440 237074 65496
rect 234389 65438 237074 65440
rect 327125 65498 327191 65501
rect 331038 65498 331098 65808
rect 327125 65496 331098 65498
rect 327125 65440 327130 65496
rect 327186 65440 331098 65496
rect 327125 65438 331098 65440
rect 139905 65435 139971 65438
rect 234389 65435 234455 65438
rect 327125 65435 327191 65438
rect 430073 65226 430139 65229
rect 434416 65226 434896 65256
rect 430073 65224 434896 65226
rect 430073 65168 430078 65224
rect 430134 65168 434896 65224
rect 430073 65166 434896 65168
rect 430073 65163 430139 65166
rect 434416 65136 434896 65166
rect 87465 64954 87531 64957
rect 131349 64954 131415 64957
rect 173485 64954 173551 64957
rect 226201 64954 226267 64957
rect 266589 64954 266655 64957
rect 87465 64952 90028 64954
rect 76382 64546 76442 64924
rect 87465 64896 87470 64952
rect 87526 64896 90028 64952
rect 87465 64894 90028 64896
rect 129772 64952 131415 64954
rect 129772 64896 131354 64952
rect 131410 64896 131415 64952
rect 129772 64894 131415 64896
rect 170804 64952 173551 64954
rect 170804 64896 173490 64952
rect 173546 64896 173551 64952
rect 170804 64894 173551 64896
rect 223796 64952 226267 64954
rect 223796 64896 226206 64952
rect 226262 64896 226267 64952
rect 223796 64894 226267 64896
rect 264828 64952 266655 64954
rect 264828 64896 266594 64952
rect 266650 64896 266655 64952
rect 264828 64894 266655 64896
rect 87465 64891 87531 64894
rect 131349 64891 131415 64894
rect 173485 64891 173551 64894
rect 226201 64891 226267 64894
rect 266589 64891 266655 64894
rect 274685 64954 274751 64957
rect 321605 64954 321671 64957
rect 274685 64952 278076 64954
rect 274685 64896 274690 64952
rect 274746 64896 278076 64952
rect 274685 64894 278076 64896
rect 317820 64952 321671 64954
rect 317820 64896 321610 64952
rect 321666 64896 321671 64952
rect 317820 64894 321671 64896
rect 274685 64891 274751 64894
rect 321605 64891 321671 64894
rect 79461 64546 79527 64549
rect 76382 64544 79527 64546
rect 76382 64488 79466 64544
rect 79522 64488 79527 64544
rect 76382 64486 79527 64488
rect 79461 64483 79527 64486
rect 139629 64274 139695 64277
rect 142990 64274 143050 64856
rect 180937 64410 181003 64413
rect 184022 64410 184082 64856
rect 233469 64546 233535 64549
rect 237014 64546 237074 64856
rect 233469 64544 237074 64546
rect 233469 64488 233474 64544
rect 233530 64488 237074 64544
rect 233469 64486 237074 64488
rect 327309 64546 327375 64549
rect 331038 64546 331098 64856
rect 327309 64544 331098 64546
rect 327309 64488 327314 64544
rect 327370 64488 331098 64544
rect 327309 64486 331098 64488
rect 233469 64483 233535 64486
rect 327309 64483 327375 64486
rect 180937 64408 184082 64410
rect 180937 64352 180942 64408
rect 180998 64352 184082 64408
rect 180937 64350 184082 64352
rect 180937 64347 181003 64350
rect 139629 64272 143050 64274
rect 139629 64216 139634 64272
rect 139690 64216 143050 64272
rect 139629 64214 143050 64216
rect 139629 64211 139695 64214
rect 87189 64138 87255 64141
rect 132177 64138 132243 64141
rect 87189 64136 90028 64138
rect 87189 64080 87194 64136
rect 87250 64080 90028 64136
rect 87189 64078 90028 64080
rect 129772 64136 132243 64138
rect 129772 64080 132182 64136
rect 132238 64080 132243 64136
rect 129772 64078 132243 64080
rect 87189 64075 87255 64078
rect 132177 64075 132243 64078
rect 181765 64138 181831 64141
rect 225925 64138 225991 64141
rect 181765 64136 184052 64138
rect 181765 64080 181770 64136
rect 181826 64080 184052 64136
rect 181765 64078 184052 64080
rect 223796 64136 225991 64138
rect 223796 64080 225930 64136
rect 225986 64080 225991 64136
rect 223796 64078 225991 64080
rect 181765 64075 181831 64078
rect 225925 64075 225991 64078
rect 274869 64138 274935 64141
rect 321605 64138 321671 64141
rect 274869 64136 278076 64138
rect 274869 64080 274874 64136
rect 274930 64080 278076 64136
rect 274869 64078 278076 64080
rect 317820 64136 321671 64138
rect 317820 64080 321610 64136
rect 321666 64080 321671 64136
rect 317820 64078 321671 64080
rect 274869 64075 274935 64078
rect 321605 64075 321671 64078
rect 173485 63866 173551 63869
rect 266681 63866 266747 63869
rect 170804 63864 173551 63866
rect 76382 63322 76442 63836
rect 170804 63808 173490 63864
rect 173546 63808 173551 63864
rect 170804 63806 173551 63808
rect 264828 63864 266747 63866
rect 264828 63808 266686 63864
rect 266742 63808 266747 63864
rect 264828 63806 266747 63808
rect 173485 63803 173551 63806
rect 266681 63803 266747 63806
rect 80197 63322 80263 63325
rect 76382 63320 80263 63322
rect 76382 63264 80202 63320
rect 80258 63264 80263 63320
rect 76382 63262 80263 63264
rect 80197 63259 80263 63262
rect 87373 63186 87439 63189
rect 132361 63186 132427 63189
rect 87373 63184 90028 63186
rect 87373 63128 87378 63184
rect 87434 63128 90028 63184
rect 87373 63126 90028 63128
rect 129772 63184 132427 63186
rect 129772 63128 132366 63184
rect 132422 63128 132427 63184
rect 129772 63126 132427 63128
rect 87373 63123 87439 63126
rect 132361 63123 132427 63126
rect 139721 63186 139787 63189
rect 142990 63186 143050 63768
rect 139721 63184 143050 63186
rect 139721 63128 139726 63184
rect 139782 63128 143050 63184
rect 139721 63126 143050 63128
rect 182317 63186 182383 63189
rect 225741 63186 225807 63189
rect 182317 63184 184052 63186
rect 182317 63128 182322 63184
rect 182378 63128 184052 63184
rect 182317 63126 184052 63128
rect 223796 63184 225807 63186
rect 223796 63128 225746 63184
rect 225802 63128 225807 63184
rect 223796 63126 225807 63128
rect 139721 63123 139787 63126
rect 182317 63123 182383 63126
rect 225741 63123 225807 63126
rect 233469 63186 233535 63189
rect 237014 63186 237074 63768
rect 233469 63184 237074 63186
rect 233469 63128 233474 63184
rect 233530 63128 237074 63184
rect 233469 63126 237074 63128
rect 274225 63186 274291 63189
rect 328413 63186 328479 63189
rect 331038 63186 331098 63768
rect 274225 63184 278076 63186
rect 274225 63128 274230 63184
rect 274286 63128 278076 63184
rect 328413 63184 331098 63186
rect 274225 63126 278076 63128
rect 233469 63123 233535 63126
rect 274225 63123 274291 63126
rect 80197 62914 80263 62917
rect 76198 62912 80263 62914
rect 76198 62856 80202 62912
rect 80258 62856 80263 62912
rect 76198 62854 80263 62856
rect 76198 62748 76258 62854
rect 80197 62851 80263 62854
rect 139813 62778 139879 62781
rect 174037 62778 174103 62781
rect 139813 62776 143020 62778
rect 139813 62720 139818 62776
rect 139874 62720 143020 62776
rect 139813 62718 143020 62720
rect 170804 62776 174103 62778
rect 170804 62720 174042 62776
rect 174098 62720 174103 62776
rect 170804 62718 174103 62720
rect 139813 62715 139879 62718
rect 174037 62715 174103 62718
rect 233561 62778 233627 62781
rect 266589 62778 266655 62781
rect 233561 62776 237044 62778
rect 233561 62720 233566 62776
rect 233622 62720 237044 62776
rect 233561 62718 237044 62720
rect 264828 62776 266655 62778
rect 264828 62720 266594 62776
rect 266650 62720 266655 62776
rect 264828 62718 266655 62720
rect 317790 62778 317850 63156
rect 328413 63128 328418 63184
rect 328474 63128 331098 63184
rect 328413 63126 331098 63128
rect 328413 63123 328479 63126
rect 320501 62778 320567 62781
rect 317790 62776 320567 62778
rect 317790 62720 320506 62776
rect 320562 62720 320567 62776
rect 317790 62718 320567 62720
rect 233561 62715 233627 62718
rect 266589 62715 266655 62718
rect 320501 62715 320567 62718
rect 327217 62778 327283 62781
rect 327217 62776 331068 62778
rect 327217 62720 327222 62776
rect 327278 62720 331068 62776
rect 327217 62718 331068 62720
rect 327217 62715 327283 62718
rect 87281 62370 87347 62373
rect 131349 62370 131415 62373
rect 87281 62368 90028 62370
rect 87281 62312 87286 62368
rect 87342 62312 90028 62368
rect 87281 62310 90028 62312
rect 129772 62368 131415 62370
rect 129772 62312 131354 62368
rect 131410 62312 131415 62368
rect 129772 62310 131415 62312
rect 87281 62307 87347 62310
rect 131349 62307 131415 62310
rect 182317 62370 182383 62373
rect 226293 62370 226359 62373
rect 182317 62368 184052 62370
rect 182317 62312 182322 62368
rect 182378 62312 184052 62368
rect 182317 62310 184052 62312
rect 223796 62368 226359 62370
rect 223796 62312 226298 62368
rect 226354 62312 226359 62368
rect 223796 62310 226359 62312
rect 182317 62307 182383 62310
rect 226293 62307 226359 62310
rect 274777 62370 274843 62373
rect 274777 62368 278076 62370
rect 274777 62312 274782 62368
rect 274838 62312 278076 62368
rect 274777 62310 278076 62312
rect 274777 62307 274843 62310
rect 173117 61826 173183 61829
rect 266589 61826 266655 61829
rect 170804 61824 173183 61826
rect 76382 61418 76442 61796
rect 170804 61768 173122 61824
rect 173178 61768 173183 61824
rect 170804 61766 173183 61768
rect 264828 61824 266655 61826
rect 264828 61768 266594 61824
rect 266650 61768 266655 61824
rect 264828 61766 266655 61768
rect 317790 61826 317850 62340
rect 318385 61826 318451 61829
rect 317790 61824 318451 61826
rect 317790 61768 318390 61824
rect 318446 61768 318451 61824
rect 317790 61766 318451 61768
rect 173117 61763 173183 61766
rect 266589 61763 266655 61766
rect 318385 61763 318451 61766
rect 80197 61418 80263 61421
rect 76382 61416 80263 61418
rect 76382 61360 80202 61416
rect 80258 61360 80263 61416
rect 76382 61358 80263 61360
rect 80197 61355 80263 61358
rect 87189 61418 87255 61421
rect 131717 61418 131783 61421
rect 87189 61416 90028 61418
rect 87189 61360 87194 61416
rect 87250 61360 90028 61416
rect 87189 61358 90028 61360
rect 129772 61416 131783 61418
rect 129772 61360 131722 61416
rect 131778 61360 131783 61416
rect 129772 61358 131783 61360
rect 87189 61355 87255 61358
rect 131717 61355 131783 61358
rect 139629 61418 139695 61421
rect 142990 61418 143050 61728
rect 139629 61416 143050 61418
rect 139629 61360 139634 61416
rect 139690 61360 143050 61416
rect 139629 61358 143050 61360
rect 181581 61418 181647 61421
rect 226293 61418 226359 61421
rect 181581 61416 184052 61418
rect 181581 61360 181586 61416
rect 181642 61360 184052 61416
rect 181581 61358 184052 61360
rect 223796 61416 226359 61418
rect 223796 61360 226298 61416
rect 226354 61360 226359 61416
rect 223796 61358 226359 61360
rect 139629 61355 139695 61358
rect 181581 61355 181647 61358
rect 226293 61355 226359 61358
rect 233469 61418 233535 61421
rect 237014 61418 237074 61728
rect 320685 61554 320751 61557
rect 317790 61552 320751 61554
rect 317790 61496 320690 61552
rect 320746 61496 320751 61552
rect 317790 61494 320751 61496
rect 233469 61416 237074 61418
rect 233469 61360 233474 61416
rect 233530 61360 237074 61416
rect 233469 61358 237074 61360
rect 274961 61418 275027 61421
rect 274961 61416 278076 61418
rect 274961 61360 274966 61416
rect 275022 61360 278076 61416
rect 317790 61388 317850 61494
rect 320685 61491 320751 61494
rect 318385 61418 318451 61421
rect 321053 61418 321119 61421
rect 318385 61416 321119 61418
rect 274961 61358 278076 61360
rect 318385 61360 318390 61416
rect 318446 61360 321058 61416
rect 321114 61360 321119 61416
rect 318385 61358 321119 61360
rect 233469 61355 233535 61358
rect 274961 61355 275027 61358
rect 318385 61355 318451 61358
rect 321053 61355 321119 61358
rect 328321 61418 328387 61421
rect 331038 61418 331098 61728
rect 328321 61416 331098 61418
rect 328321 61360 328326 61416
rect 328382 61360 331098 61416
rect 328321 61358 331098 61360
rect 328321 61355 328387 61358
rect 173117 60738 173183 60741
rect 266589 60738 266655 60741
rect 170804 60736 173183 60738
rect 76382 60194 76442 60708
rect 170804 60680 173122 60736
rect 173178 60680 173183 60736
rect 170804 60678 173183 60680
rect 264828 60736 266655 60738
rect 264828 60680 266594 60736
rect 266650 60680 266655 60736
rect 264828 60678 266655 60680
rect 173117 60675 173183 60678
rect 266589 60675 266655 60678
rect 87189 60466 87255 60469
rect 131349 60466 131415 60469
rect 87189 60464 90028 60466
rect 87189 60408 87194 60464
rect 87250 60408 90028 60464
rect 87189 60406 90028 60408
rect 129772 60464 131415 60466
rect 129772 60408 131354 60464
rect 131410 60408 131415 60464
rect 129772 60406 131415 60408
rect 87189 60403 87255 60406
rect 131349 60403 131415 60406
rect 80197 60194 80263 60197
rect 76382 60192 80263 60194
rect 76382 60136 80202 60192
rect 80258 60136 80263 60192
rect 76382 60134 80263 60136
rect 80197 60131 80263 60134
rect 139721 60058 139787 60061
rect 142990 60058 143050 60640
rect 181213 60466 181279 60469
rect 225741 60466 225807 60469
rect 181213 60464 184052 60466
rect 181213 60408 181218 60464
rect 181274 60408 184052 60464
rect 181213 60406 184052 60408
rect 223796 60464 225807 60466
rect 223796 60408 225746 60464
rect 225802 60408 225807 60464
rect 223796 60406 225807 60408
rect 181213 60403 181279 60406
rect 225741 60403 225807 60406
rect 139721 60056 143050 60058
rect 139721 60000 139726 60056
rect 139782 60000 143050 60056
rect 139721 59998 143050 60000
rect 233469 60058 233535 60061
rect 237014 60058 237074 60640
rect 274869 60466 274935 60469
rect 274869 60464 278076 60466
rect 274869 60408 274874 60464
rect 274930 60408 278076 60464
rect 274869 60406 278076 60408
rect 274869 60403 274935 60406
rect 233469 60056 237074 60058
rect 233469 60000 233474 60056
rect 233530 60000 237074 60056
rect 233469 59998 237074 60000
rect 139721 59995 139787 59998
rect 233469 59995 233535 59998
rect 317790 59922 317850 60436
rect 328413 60058 328479 60061
rect 331038 60058 331098 60640
rect 328413 60056 331098 60058
rect 328413 60000 328418 60056
rect 328474 60000 331098 60056
rect 328413 59998 331098 60000
rect 328413 59995 328479 59998
rect 321053 59922 321119 59925
rect 317790 59920 321119 59922
rect 317790 59864 321058 59920
rect 321114 59864 321119 59920
rect 317790 59862 321119 59864
rect 321053 59859 321119 59862
rect 87833 59650 87899 59653
rect 131349 59650 131415 59653
rect 173025 59650 173091 59653
rect 87833 59648 90028 59650
rect 76382 59106 76442 59620
rect 87833 59592 87838 59648
rect 87894 59592 90028 59648
rect 87833 59590 90028 59592
rect 129772 59648 131415 59650
rect 129772 59592 131354 59648
rect 131410 59592 131415 59648
rect 129772 59590 131415 59592
rect 170804 59648 173091 59650
rect 170804 59592 173030 59648
rect 173086 59592 173091 59648
rect 170804 59590 173091 59592
rect 87833 59587 87899 59590
rect 131349 59587 131415 59590
rect 173025 59587 173091 59590
rect 181029 59650 181095 59653
rect 226293 59650 226359 59653
rect 267325 59650 267391 59653
rect 181029 59648 184052 59650
rect 181029 59592 181034 59648
rect 181090 59592 184052 59648
rect 181029 59590 184052 59592
rect 223796 59648 226359 59650
rect 223796 59592 226298 59648
rect 226354 59592 226359 59648
rect 223796 59590 226359 59592
rect 264828 59648 267391 59650
rect 264828 59592 267330 59648
rect 267386 59592 267391 59648
rect 264828 59590 267391 59592
rect 181029 59587 181095 59590
rect 226293 59587 226359 59590
rect 267325 59587 267391 59590
rect 275697 59650 275763 59653
rect 320501 59650 320567 59653
rect 275697 59648 278076 59650
rect 275697 59592 275702 59648
rect 275758 59592 278076 59648
rect 275697 59590 278076 59592
rect 317820 59648 320567 59650
rect 317820 59592 320506 59648
rect 320562 59592 320567 59648
rect 317820 59590 320567 59592
rect 275697 59587 275763 59590
rect 320501 59587 320567 59590
rect 79645 59106 79711 59109
rect 76382 59104 79711 59106
rect 76382 59048 79650 59104
rect 79706 59048 79711 59104
rect 76382 59046 79711 59048
rect 79645 59043 79711 59046
rect 140457 58970 140523 58973
rect 142990 58970 143050 59552
rect 140457 58968 143050 58970
rect 140457 58912 140462 58968
rect 140518 58912 143050 58968
rect 140457 58910 143050 58912
rect 233653 58970 233719 58973
rect 237014 58970 237074 59552
rect 233653 58968 237074 58970
rect 233653 58912 233658 58968
rect 233714 58912 237074 58968
rect 233653 58910 237074 58912
rect 328597 58970 328663 58973
rect 331038 58970 331098 59552
rect 328597 58968 331098 58970
rect 328597 58912 328602 58968
rect 328658 58912 331098 58968
rect 328597 58910 331098 58912
rect 140457 58907 140523 58910
rect 233653 58907 233719 58910
rect 328597 58907 328663 58910
rect 87189 58698 87255 58701
rect 131441 58698 131507 58701
rect 87189 58696 90028 58698
rect 76382 58562 76442 58668
rect 87189 58640 87194 58696
rect 87250 58640 90028 58696
rect 87189 58638 90028 58640
rect 129772 58696 131507 58698
rect 129772 58640 131446 58696
rect 131502 58640 131507 58696
rect 129772 58638 131507 58640
rect 87189 58635 87255 58638
rect 131441 58635 131507 58638
rect 140365 58698 140431 58701
rect 173577 58698 173643 58701
rect 140365 58696 143020 58698
rect 140365 58640 140370 58696
rect 140426 58640 143020 58696
rect 140365 58638 143020 58640
rect 170804 58696 173643 58698
rect 170804 58640 173582 58696
rect 173638 58640 173643 58696
rect 170804 58638 173643 58640
rect 140365 58635 140431 58638
rect 173577 58635 173643 58638
rect 181121 58698 181187 58701
rect 225741 58698 225807 58701
rect 181121 58696 184052 58698
rect 181121 58640 181126 58696
rect 181182 58640 184052 58696
rect 181121 58638 184052 58640
rect 223796 58696 225807 58698
rect 223796 58640 225746 58696
rect 225802 58640 225807 58696
rect 223796 58638 225807 58640
rect 181121 58635 181187 58638
rect 225741 58635 225807 58638
rect 233469 58698 233535 58701
rect 267877 58698 267943 58701
rect 233469 58696 237044 58698
rect 233469 58640 233474 58696
rect 233530 58640 237044 58696
rect 233469 58638 237044 58640
rect 264828 58696 267943 58698
rect 264828 58640 267882 58696
rect 267938 58640 267943 58696
rect 264828 58638 267943 58640
rect 233469 58635 233535 58638
rect 267877 58635 267943 58638
rect 275421 58698 275487 58701
rect 320409 58698 320475 58701
rect 275421 58696 278076 58698
rect 275421 58640 275426 58696
rect 275482 58640 278076 58696
rect 275421 58638 278076 58640
rect 317820 58696 320475 58698
rect 317820 58640 320414 58696
rect 320470 58640 320475 58696
rect 317820 58638 320475 58640
rect 275421 58635 275487 58638
rect 320409 58635 320475 58638
rect 327493 58698 327559 58701
rect 327493 58696 331068 58698
rect 327493 58640 327498 58696
rect 327554 58640 331068 58696
rect 327493 58638 331068 58640
rect 327493 58635 327559 58638
rect 80197 58562 80263 58565
rect 76382 58560 80263 58562
rect 76382 58504 80202 58560
rect 80258 58504 80263 58560
rect 76382 58502 80263 58504
rect 80197 58499 80263 58502
rect 87189 57882 87255 57885
rect 131349 57882 131415 57885
rect 87189 57880 90028 57882
rect 87189 57824 87194 57880
rect 87250 57824 90028 57880
rect 87189 57822 90028 57824
rect 129772 57880 131415 57882
rect 129772 57824 131354 57880
rect 131410 57824 131415 57880
rect 129772 57822 131415 57824
rect 87189 57819 87255 57822
rect 131349 57819 131415 57822
rect 181029 57882 181095 57885
rect 225557 57882 225623 57885
rect 181029 57880 184052 57882
rect 181029 57824 181034 57880
rect 181090 57824 184052 57880
rect 181029 57822 184052 57824
rect 223796 57880 225623 57882
rect 223796 57824 225562 57880
rect 225618 57824 225623 57880
rect 223796 57822 225623 57824
rect 181029 57819 181095 57822
rect 225557 57819 225623 57822
rect 275697 57882 275763 57885
rect 320409 57882 320475 57885
rect 275697 57880 278076 57882
rect 275697 57824 275702 57880
rect 275758 57824 278076 57880
rect 275697 57822 278076 57824
rect 317820 57880 320475 57882
rect 317820 57824 320414 57880
rect 320470 57824 320475 57880
rect 317820 57822 320475 57824
rect 275697 57819 275763 57822
rect 320409 57819 320475 57822
rect 173301 57610 173367 57613
rect 267693 57610 267759 57613
rect 170804 57608 173367 57610
rect 76382 57202 76442 57580
rect 170804 57552 173306 57608
rect 173362 57552 173367 57608
rect 170804 57550 173367 57552
rect 264828 57608 267759 57610
rect 264828 57552 267698 57608
rect 267754 57552 267759 57608
rect 264828 57550 267759 57552
rect 173301 57547 173367 57550
rect 267693 57547 267759 57550
rect 80197 57202 80263 57205
rect 76382 57200 80263 57202
rect 76382 57144 80202 57200
rect 80258 57144 80263 57200
rect 76382 57142 80263 57144
rect 80197 57139 80263 57142
rect 140273 57202 140339 57205
rect 142990 57202 143050 57512
rect 140273 57200 143050 57202
rect 140273 57144 140278 57200
rect 140334 57144 143050 57200
rect 140273 57142 143050 57144
rect 233561 57202 233627 57205
rect 237014 57202 237074 57512
rect 233561 57200 237074 57202
rect 233561 57144 233566 57200
rect 233622 57144 237074 57200
rect 233561 57142 237074 57144
rect 328413 57202 328479 57205
rect 331038 57202 331098 57512
rect 328413 57200 331098 57202
rect 328413 57144 328418 57200
rect 328474 57144 331098 57200
rect 328413 57142 331098 57144
rect 140273 57139 140339 57142
rect 233561 57139 233627 57142
rect 328413 57139 328479 57142
rect 87189 56930 87255 56933
rect 131349 56930 131415 56933
rect 226293 56930 226359 56933
rect 87189 56928 90028 56930
rect 87189 56872 87194 56928
rect 87250 56872 90028 56928
rect 87189 56870 90028 56872
rect 129772 56928 131415 56930
rect 129772 56872 131354 56928
rect 131410 56872 131415 56928
rect 129772 56870 131415 56872
rect 223796 56928 226359 56930
rect 223796 56872 226298 56928
rect 226354 56872 226359 56928
rect 223796 56870 226359 56872
rect 87189 56867 87255 56870
rect 131349 56867 131415 56870
rect 226293 56867 226359 56870
rect 275697 56930 275763 56933
rect 320501 56930 320567 56933
rect 275697 56928 278076 56930
rect 275697 56872 275702 56928
rect 275758 56872 278076 56928
rect 275697 56870 278076 56872
rect 317820 56928 320567 56930
rect 317820 56872 320506 56928
rect 320562 56872 320567 56928
rect 317820 56870 320567 56872
rect 275697 56867 275763 56870
rect 320501 56867 320567 56870
rect 173485 56658 173551 56661
rect 170804 56656 173551 56658
rect 76382 56114 76442 56628
rect 170804 56600 173490 56656
rect 173546 56600 173551 56656
rect 170804 56598 173551 56600
rect 173485 56595 173551 56598
rect 181029 56658 181095 56661
rect 184022 56658 184082 56832
rect 267325 56658 267391 56661
rect 181029 56656 184082 56658
rect 181029 56600 181034 56656
rect 181090 56600 184082 56656
rect 181029 56598 184082 56600
rect 264828 56656 267391 56658
rect 264828 56600 267330 56656
rect 267386 56600 267391 56656
rect 264828 56598 267391 56600
rect 181029 56595 181095 56598
rect 267325 56595 267391 56598
rect 140457 56250 140523 56253
rect 142990 56250 143050 56560
rect 140457 56248 143050 56250
rect 140457 56192 140462 56248
rect 140518 56192 143050 56248
rect 140457 56190 143050 56192
rect 140457 56187 140523 56190
rect 78909 56114 78975 56117
rect 76382 56112 78975 56114
rect 76382 56056 78914 56112
rect 78970 56056 78975 56112
rect 76382 56054 78975 56056
rect 78909 56051 78975 56054
rect 87281 56114 87347 56117
rect 132177 56114 132243 56117
rect 87281 56112 90028 56114
rect 87281 56056 87286 56112
rect 87342 56056 90028 56112
rect 87281 56054 90028 56056
rect 129772 56112 132243 56114
rect 129772 56056 132182 56112
rect 132238 56056 132243 56112
rect 129772 56054 132243 56056
rect 87281 56051 87347 56054
rect 132177 56051 132243 56054
rect 181121 56114 181187 56117
rect 225649 56114 225715 56117
rect 181121 56112 184052 56114
rect 181121 56056 181126 56112
rect 181182 56056 184052 56112
rect 181121 56054 184052 56056
rect 223796 56112 225715 56114
rect 223796 56056 225654 56112
rect 225710 56056 225715 56112
rect 223796 56054 225715 56056
rect 181121 56051 181187 56054
rect 225649 56051 225715 56054
rect 233469 56114 233535 56117
rect 237014 56114 237074 56560
rect 233469 56112 237074 56114
rect 233469 56056 233474 56112
rect 233530 56056 237074 56112
rect 233469 56054 237074 56056
rect 275237 56114 275303 56117
rect 320409 56114 320475 56117
rect 275237 56112 278076 56114
rect 275237 56056 275242 56112
rect 275298 56056 278076 56112
rect 275237 56054 278076 56056
rect 317820 56112 320475 56114
rect 317820 56056 320414 56112
rect 320470 56056 320475 56112
rect 317820 56054 320475 56056
rect 233469 56051 233535 56054
rect 275237 56051 275303 56054
rect 320409 56051 320475 56054
rect 327493 55978 327559 55981
rect 331038 55978 331098 56560
rect 327493 55976 331098 55978
rect 327493 55920 327498 55976
rect 327554 55920 331098 55976
rect 327493 55918 331098 55920
rect 327493 55915 327559 55918
rect 9896 55706 10376 55736
rect 13129 55706 13195 55709
rect 79553 55706 79619 55709
rect 9896 55704 13195 55706
rect 9896 55648 13134 55704
rect 13190 55648 13195 55704
rect 9896 55646 13195 55648
rect 9896 55616 10376 55646
rect 13129 55643 13195 55646
rect 76198 55704 79619 55706
rect 76198 55648 79558 55704
rect 79614 55648 79619 55704
rect 76198 55646 79619 55648
rect 76198 55540 76258 55646
rect 79553 55643 79619 55646
rect 173393 55570 173459 55573
rect 267233 55570 267299 55573
rect 170804 55568 173459 55570
rect 170804 55512 173398 55568
rect 173454 55512 173459 55568
rect 170804 55510 173459 55512
rect 264828 55568 267299 55570
rect 264828 55512 267238 55568
rect 267294 55512 267299 55568
rect 264828 55510 267299 55512
rect 173393 55507 173459 55510
rect 267233 55507 267299 55510
rect 140641 55298 140707 55301
rect 142990 55298 143050 55472
rect 140641 55296 143050 55298
rect 140641 55240 140646 55296
rect 140702 55240 143050 55296
rect 140641 55238 143050 55240
rect 233469 55298 233535 55301
rect 237014 55298 237074 55472
rect 233469 55296 237074 55298
rect 233469 55240 233474 55296
rect 233530 55240 237074 55296
rect 233469 55238 237074 55240
rect 328505 55298 328571 55301
rect 331038 55298 331098 55472
rect 328505 55296 331098 55298
rect 328505 55240 328510 55296
rect 328566 55240 331098 55296
rect 328505 55238 331098 55240
rect 140641 55235 140707 55238
rect 233469 55235 233535 55238
rect 328505 55235 328571 55238
rect 87189 55162 87255 55165
rect 131349 55162 131415 55165
rect 87189 55160 90028 55162
rect 87189 55104 87194 55160
rect 87250 55104 90028 55160
rect 87189 55102 90028 55104
rect 129772 55160 131415 55162
rect 129772 55104 131354 55160
rect 131410 55104 131415 55160
rect 129772 55102 131415 55104
rect 87189 55099 87255 55102
rect 131349 55099 131415 55102
rect 181029 55162 181095 55165
rect 226385 55162 226451 55165
rect 181029 55160 184052 55162
rect 181029 55104 181034 55160
rect 181090 55104 184052 55160
rect 181029 55102 184052 55104
rect 223796 55160 226451 55162
rect 223796 55104 226390 55160
rect 226446 55104 226451 55160
rect 223796 55102 226451 55104
rect 181029 55099 181095 55102
rect 226385 55099 226451 55102
rect 275421 55162 275487 55165
rect 320409 55162 320475 55165
rect 275421 55160 278076 55162
rect 275421 55104 275426 55160
rect 275482 55104 278076 55160
rect 275421 55102 278076 55104
rect 317820 55160 320475 55162
rect 317820 55104 320414 55160
rect 320470 55104 320475 55160
rect 317820 55102 320475 55104
rect 275421 55099 275487 55102
rect 320409 55099 320475 55102
rect 80197 54618 80263 54621
rect 76198 54616 80263 54618
rect 76198 54560 80202 54616
rect 80258 54560 80263 54616
rect 76198 54558 80263 54560
rect 76198 54452 76258 54558
rect 80197 54555 80263 54558
rect 140365 54482 140431 54485
rect 173577 54482 173643 54485
rect 140365 54480 143020 54482
rect 140365 54424 140370 54480
rect 140426 54424 143020 54480
rect 140365 54422 143020 54424
rect 170804 54480 173643 54482
rect 170804 54424 173582 54480
rect 173638 54424 173643 54480
rect 170804 54422 173643 54424
rect 140365 54419 140431 54422
rect 173577 54419 173643 54422
rect 233469 54482 233535 54485
rect 267877 54482 267943 54485
rect 233469 54480 237044 54482
rect 233469 54424 233474 54480
rect 233530 54424 237044 54480
rect 233469 54422 237044 54424
rect 264828 54480 267943 54482
rect 264828 54424 267882 54480
rect 267938 54424 267943 54480
rect 264828 54422 267943 54424
rect 233469 54419 233535 54422
rect 267877 54419 267943 54422
rect 328413 54482 328479 54485
rect 328413 54480 331068 54482
rect 328413 54424 328418 54480
rect 328474 54424 331068 54480
rect 328413 54422 331068 54424
rect 328413 54419 328479 54422
rect 87189 54346 87255 54349
rect 131349 54346 131415 54349
rect 87189 54344 90028 54346
rect 87189 54288 87194 54344
rect 87250 54288 90028 54344
rect 87189 54286 90028 54288
rect 129772 54344 131415 54346
rect 129772 54288 131354 54344
rect 131410 54288 131415 54344
rect 129772 54286 131415 54288
rect 87189 54283 87255 54286
rect 131349 54283 131415 54286
rect 181029 54346 181095 54349
rect 226477 54346 226543 54349
rect 181029 54344 184052 54346
rect 181029 54288 181034 54344
rect 181090 54288 184052 54344
rect 181029 54286 184052 54288
rect 223796 54344 226543 54346
rect 223796 54288 226482 54344
rect 226538 54288 226543 54344
rect 223796 54286 226543 54288
rect 181029 54283 181095 54286
rect 226477 54283 226543 54286
rect 275697 54346 275763 54349
rect 320409 54346 320475 54349
rect 275697 54344 278076 54346
rect 275697 54288 275702 54344
rect 275758 54288 278076 54344
rect 275697 54286 278076 54288
rect 317820 54344 320475 54346
rect 317820 54288 320414 54344
rect 320470 54288 320475 54344
rect 317820 54286 320475 54288
rect 275697 54283 275763 54286
rect 320409 54283 320475 54286
rect 80197 53666 80263 53669
rect 76198 53664 80263 53666
rect 76198 53608 80202 53664
rect 80258 53608 80263 53664
rect 76198 53606 80263 53608
rect 76198 53500 76258 53606
rect 80197 53603 80263 53606
rect 140549 53530 140615 53533
rect 173577 53530 173643 53533
rect 140549 53528 143020 53530
rect 140549 53472 140554 53528
rect 140610 53472 143020 53528
rect 140549 53470 143020 53472
rect 170804 53528 173643 53530
rect 170804 53472 173582 53528
rect 173638 53472 173643 53528
rect 170804 53470 173643 53472
rect 140549 53467 140615 53470
rect 173577 53467 173643 53470
rect 233469 53530 233535 53533
rect 267877 53530 267943 53533
rect 233469 53528 237044 53530
rect 233469 53472 233474 53528
rect 233530 53472 237044 53528
rect 233469 53470 237044 53472
rect 264828 53528 267943 53530
rect 264828 53472 267882 53528
rect 267938 53472 267943 53528
rect 264828 53470 267943 53472
rect 233469 53467 233535 53470
rect 267877 53467 267943 53470
rect 328413 53530 328479 53533
rect 328413 53528 331068 53530
rect 328413 53472 328418 53528
rect 328474 53472 331068 53528
rect 328413 53470 331068 53472
rect 328413 53467 328479 53470
rect 113961 53124 114027 53125
rect 113910 53122 113916 53124
rect 113870 53062 113916 53122
rect 113980 53120 114027 53124
rect 114022 53064 114027 53120
rect 113910 53060 113916 53062
rect 113980 53060 114027 53064
rect 113961 53059 114027 53060
rect 118653 53124 118719 53125
rect 212493 53124 212559 53125
rect 301641 53124 301707 53125
rect 306609 53124 306675 53125
rect 118653 53120 118700 53124
rect 118764 53122 118770 53124
rect 118653 53064 118658 53120
rect 118653 53060 118700 53064
rect 118764 53062 118810 53122
rect 212493 53120 212540 53124
rect 212604 53122 212610 53124
rect 301590 53122 301596 53124
rect 212493 53064 212498 53120
rect 118764 53060 118770 53062
rect 212493 53060 212540 53064
rect 212604 53062 212650 53122
rect 301550 53062 301596 53122
rect 301660 53120 301707 53124
rect 301702 53064 301707 53120
rect 212604 53060 212610 53062
rect 301590 53060 301596 53062
rect 301660 53060 301707 53064
rect 306558 53060 306564 53124
rect 306628 53122 306675 53124
rect 306628 53120 306720 53122
rect 306670 53064 306720 53120
rect 306628 53062 306720 53064
rect 306628 53060 306675 53062
rect 118653 53059 118719 53060
rect 212493 53059 212559 53060
rect 301641 53059 301707 53060
rect 306609 53059 306675 53060
rect 80197 52714 80263 52717
rect 76198 52712 80263 52714
rect 76198 52656 80202 52712
rect 80258 52656 80263 52712
rect 76198 52654 80263 52656
rect 76198 52412 76258 52654
rect 80197 52651 80263 52654
rect 428785 52714 428851 52717
rect 434416 52714 434896 52744
rect 428785 52712 434896 52714
rect 428785 52656 428790 52712
rect 428846 52656 434896 52712
rect 428785 52654 434896 52656
rect 428785 52651 428851 52654
rect 434416 52624 434896 52654
rect 139997 52442 140063 52445
rect 171829 52442 171895 52445
rect 139997 52440 143020 52442
rect 139997 52384 140002 52440
rect 140058 52384 143020 52440
rect 139997 52382 143020 52384
rect 170804 52440 171895 52442
rect 170804 52384 171834 52440
rect 171890 52384 171895 52440
rect 170804 52382 171895 52384
rect 139997 52379 140063 52382
rect 171829 52379 171895 52382
rect 233469 52442 233535 52445
rect 267877 52442 267943 52445
rect 233469 52440 237044 52442
rect 233469 52384 233474 52440
rect 233530 52384 237044 52440
rect 233469 52382 237044 52384
rect 264828 52440 267943 52442
rect 264828 52384 267882 52440
rect 267938 52384 267943 52440
rect 264828 52382 267943 52384
rect 233469 52379 233535 52382
rect 267877 52379 267943 52382
rect 328505 52442 328571 52445
rect 328505 52440 331068 52442
rect 328505 52384 328510 52440
rect 328566 52384 331068 52440
rect 328505 52382 331068 52384
rect 328505 52379 328571 52382
rect 191374 51564 191380 51628
rect 191444 51626 191450 51628
rect 191977 51626 192043 51629
rect 191444 51624 192043 51626
rect 191444 51568 191982 51624
rect 192038 51568 192043 51624
rect 191444 51566 192043 51568
rect 191444 51564 191450 51566
rect 191977 51563 192043 51566
rect 203753 51626 203819 51629
rect 204254 51626 204260 51628
rect 203753 51624 204260 51626
rect 203753 51568 203758 51624
rect 203814 51568 204260 51624
rect 203753 51566 204260 51568
rect 203753 51563 203819 51566
rect 204254 51564 204260 51566
rect 204324 51564 204330 51628
rect 102369 51354 102435 51357
rect 102502 51354 102508 51356
rect 102369 51352 102508 51354
rect 76382 50810 76442 51324
rect 102369 51296 102374 51352
rect 102430 51296 102508 51352
rect 102369 51294 102508 51296
rect 102369 51291 102435 51294
rect 102502 51292 102508 51294
rect 102572 51292 102578 51356
rect 173301 51354 173367 51357
rect 170804 51352 173367 51354
rect 170804 51296 173306 51352
rect 173362 51296 173367 51352
rect 170804 51294 173367 51296
rect 173301 51291 173367 51294
rect 207750 51292 207756 51356
rect 207820 51354 207826 51356
rect 207893 51354 207959 51357
rect 267509 51354 267575 51357
rect 207820 51352 207959 51354
rect 207820 51296 207898 51352
rect 207954 51296 207959 51352
rect 207820 51294 207959 51296
rect 264828 51352 267575 51354
rect 264828 51296 267514 51352
rect 267570 51296 267575 51352
rect 264828 51294 267575 51296
rect 207820 51292 207826 51294
rect 207893 51291 207959 51294
rect 267509 51291 267575 51294
rect 270678 51292 270684 51356
rect 270748 51354 270754 51356
rect 281309 51354 281375 51357
rect 270748 51352 281375 51354
rect 270748 51296 281314 51352
rect 281370 51296 281375 51352
rect 270748 51294 281375 51296
rect 270748 51292 270754 51294
rect 281309 51291 281375 51294
rect 142430 51020 142436 51084
rect 142500 51082 142506 51084
rect 142849 51082 142915 51085
rect 142500 51080 142915 51082
rect 142500 51024 142854 51080
rect 142910 51024 142915 51080
rect 142500 51022 142915 51024
rect 142500 51020 142506 51022
rect 142849 51019 142915 51022
rect 78909 50810 78975 50813
rect 76382 50808 78975 50810
rect 76382 50752 78914 50808
rect 78970 50752 78975 50808
rect 76382 50750 78975 50752
rect 78909 50747 78975 50750
rect 140641 50810 140707 50813
rect 142990 50810 143050 51256
rect 140641 50808 143050 50810
rect 140641 50752 140646 50808
rect 140702 50752 143050 50808
rect 140641 50750 143050 50752
rect 233561 50810 233627 50813
rect 237014 50810 237074 51256
rect 327677 50946 327743 50949
rect 331038 50946 331098 51256
rect 327677 50944 331098 50946
rect 327677 50888 327682 50944
rect 327738 50888 331098 50944
rect 327677 50886 331098 50888
rect 327677 50883 327743 50886
rect 233561 50808 237074 50810
rect 233561 50752 233566 50808
rect 233622 50752 237074 50808
rect 233561 50750 237074 50752
rect 140641 50747 140707 50750
rect 233561 50747 233627 50750
rect 93629 50676 93695 50677
rect 170541 50676 170607 50677
rect 93629 50674 93676 50676
rect 93584 50672 93676 50674
rect 93584 50616 93634 50672
rect 93584 50614 93676 50616
rect 93629 50612 93676 50614
rect 93740 50612 93746 50676
rect 170541 50674 170588 50676
rect 170496 50672 170588 50674
rect 170496 50616 170546 50672
rect 170496 50614 170588 50616
rect 170541 50612 170588 50614
rect 170652 50612 170658 50676
rect 187142 50612 187148 50676
rect 187212 50674 187218 50676
rect 187285 50674 187351 50677
rect 187212 50672 187351 50674
rect 187212 50616 187290 50672
rect 187346 50616 187351 50672
rect 187212 50614 187351 50616
rect 187212 50612 187218 50614
rect 93629 50611 93695 50612
rect 170541 50611 170607 50612
rect 187285 50611 187351 50614
rect 140365 50402 140431 50405
rect 173577 50402 173643 50405
rect 140365 50400 143020 50402
rect 76382 50266 76442 50372
rect 140365 50344 140370 50400
rect 140426 50344 143020 50400
rect 140365 50342 143020 50344
rect 170804 50400 173643 50402
rect 170804 50344 173582 50400
rect 173638 50344 173643 50400
rect 170804 50342 173643 50344
rect 140365 50339 140431 50342
rect 173577 50339 173643 50342
rect 233469 50402 233535 50405
rect 266773 50402 266839 50405
rect 233469 50400 237044 50402
rect 233469 50344 233474 50400
rect 233530 50344 237044 50400
rect 233469 50342 237044 50344
rect 264828 50400 266839 50402
rect 264828 50344 266778 50400
rect 266834 50344 266839 50400
rect 264828 50342 266839 50344
rect 233469 50339 233535 50342
rect 266773 50339 266839 50342
rect 328413 50402 328479 50405
rect 328413 50400 331068 50402
rect 328413 50344 328418 50400
rect 328474 50344 331068 50400
rect 328413 50342 331068 50344
rect 328413 50339 328479 50342
rect 358446 50340 358452 50404
rect 358516 50402 358522 50404
rect 358589 50402 358655 50405
rect 358516 50400 358655 50402
rect 358516 50344 358594 50400
rect 358650 50344 358655 50400
rect 358516 50342 358655 50344
rect 358516 50340 358522 50342
rect 358589 50339 358655 50342
rect 80197 50266 80263 50269
rect 107521 50268 107587 50269
rect 76382 50264 80263 50266
rect 76382 50208 80202 50264
rect 80258 50208 80263 50264
rect 76382 50206 80263 50208
rect 80197 50203 80263 50206
rect 107470 50204 107476 50268
rect 107540 50266 107587 50268
rect 107540 50264 107632 50266
rect 107582 50208 107632 50264
rect 107540 50206 107632 50208
rect 107540 50204 107587 50206
rect 109310 50204 109316 50268
rect 109380 50266 109386 50268
rect 109453 50266 109519 50269
rect 109380 50264 109519 50266
rect 109380 50208 109458 50264
rect 109514 50208 109519 50264
rect 109380 50206 109519 50208
rect 109380 50204 109386 50206
rect 107521 50203 107587 50204
rect 109453 50203 109519 50206
rect 88385 49316 88451 49317
rect 76382 49178 76442 49284
rect 88334 49252 88340 49316
rect 88404 49314 88451 49316
rect 105129 49314 105195 49317
rect 105262 49314 105268 49316
rect 88404 49312 88496 49314
rect 88446 49256 88496 49312
rect 88404 49254 88496 49256
rect 105129 49312 105268 49314
rect 105129 49256 105134 49312
rect 105190 49256 105268 49312
rect 105129 49254 105268 49256
rect 88404 49252 88451 49254
rect 88385 49251 88451 49252
rect 105129 49251 105195 49254
rect 105262 49252 105268 49254
rect 105332 49252 105338 49316
rect 172933 49314 172999 49317
rect 170804 49312 172999 49314
rect 170804 49256 172938 49312
rect 172994 49256 172999 49312
rect 170804 49254 172999 49256
rect 172933 49251 172999 49254
rect 181990 49252 181996 49316
rect 182060 49314 182066 49316
rect 182133 49314 182199 49317
rect 267877 49314 267943 49317
rect 182060 49312 182199 49314
rect 182060 49256 182138 49312
rect 182194 49256 182199 49312
rect 182060 49254 182199 49256
rect 264828 49312 267943 49314
rect 264828 49256 267882 49312
rect 267938 49256 267943 49312
rect 264828 49254 267943 49256
rect 182060 49252 182066 49254
rect 182133 49251 182199 49254
rect 267877 49251 267943 49254
rect 328413 49314 328479 49317
rect 328413 49312 331068 49314
rect 328413 49256 328418 49312
rect 328474 49256 331068 49312
rect 328413 49254 331068 49256
rect 328413 49251 328479 49254
rect 80197 49178 80263 49181
rect 76382 49176 80263 49178
rect 76382 49120 80202 49176
rect 80258 49120 80263 49176
rect 76382 49118 80263 49120
rect 80197 49115 80263 49118
rect 140549 49042 140615 49045
rect 142990 49042 143050 49216
rect 140549 49040 143050 49042
rect 140549 48984 140554 49040
rect 140610 48984 143050 49040
rect 140549 48982 143050 48984
rect 233469 49042 233535 49045
rect 237014 49042 237074 49216
rect 233469 49040 237074 49042
rect 233469 48984 233474 49040
rect 233530 48984 237074 49040
rect 233469 48982 237074 48984
rect 140549 48979 140615 48982
rect 233469 48979 233535 48982
rect 88150 48572 88156 48636
rect 88220 48634 88226 48636
rect 88293 48634 88359 48637
rect 88220 48632 88359 48634
rect 88220 48576 88298 48632
rect 88354 48576 88359 48632
rect 88220 48574 88359 48576
rect 88220 48572 88226 48574
rect 88293 48571 88359 48574
rect 173301 48362 173367 48365
rect 267877 48362 267943 48365
rect 170804 48360 173367 48362
rect 67869 48092 67935 48093
rect 67869 48088 67916 48092
rect 67980 48090 67986 48092
rect 67869 48032 67874 48088
rect 67869 48028 67916 48032
rect 67980 48030 68026 48090
rect 67980 48028 67986 48030
rect 73982 48028 73988 48092
rect 74052 48090 74058 48092
rect 74309 48090 74375 48093
rect 74052 48088 74375 48090
rect 74052 48032 74314 48088
rect 74370 48032 74375 48088
rect 74052 48030 74375 48032
rect 76382 48090 76442 48332
rect 170804 48304 173306 48360
rect 173362 48304 173367 48360
rect 170804 48302 173367 48304
rect 264828 48360 267943 48362
rect 264828 48304 267882 48360
rect 267938 48304 267943 48360
rect 264828 48302 267943 48304
rect 173301 48299 173367 48302
rect 267877 48299 267943 48302
rect 80197 48090 80263 48093
rect 76382 48088 80263 48090
rect 76382 48032 80202 48088
rect 80258 48032 80263 48088
rect 76382 48030 80263 48032
rect 74052 48028 74058 48030
rect 67869 48027 67935 48028
rect 74309 48027 74375 48030
rect 80197 48027 80263 48030
rect 88293 48090 88359 48093
rect 105129 48090 105195 48093
rect 88293 48088 105195 48090
rect 88293 48032 88298 48088
rect 88354 48032 105134 48088
rect 105190 48032 105195 48088
rect 88293 48030 105195 48032
rect 88293 48027 88359 48030
rect 105129 48027 105195 48030
rect 139997 48090 140063 48093
rect 142990 48090 143050 48264
rect 139997 48088 143050 48090
rect 139997 48032 140002 48088
rect 140058 48032 143050 48088
rect 139997 48030 143050 48032
rect 147725 48090 147791 48093
rect 147950 48090 147956 48092
rect 147725 48088 147956 48090
rect 147725 48032 147730 48088
rect 147786 48032 147956 48088
rect 147725 48030 147956 48032
rect 139997 48027 140063 48030
rect 147725 48027 147791 48030
rect 147950 48028 147956 48030
rect 148020 48028 148026 48092
rect 153981 48090 154047 48093
rect 154758 48090 154764 48092
rect 153981 48088 154764 48090
rect 153981 48032 153986 48088
rect 154042 48032 154764 48088
rect 153981 48030 154764 48032
rect 153981 48027 154047 48030
rect 154758 48028 154764 48030
rect 154828 48028 154834 48092
rect 160053 47956 160119 47957
rect 145558 47892 145564 47956
rect 145628 47954 145634 47956
rect 147950 47954 147956 47956
rect 145628 47894 147956 47954
rect 145628 47892 145634 47894
rect 147950 47892 147956 47894
rect 148020 47892 148026 47956
rect 160053 47952 160100 47956
rect 160164 47954 160170 47956
rect 160053 47896 160058 47952
rect 160053 47892 160100 47896
rect 160164 47894 160210 47954
rect 160164 47892 160170 47894
rect 168742 47892 168748 47956
rect 168812 47954 168818 47956
rect 168885 47954 168951 47957
rect 181857 47956 181923 47957
rect 168812 47952 168951 47954
rect 168812 47896 168890 47952
rect 168946 47896 168951 47952
rect 168812 47894 168951 47896
rect 168812 47892 168818 47894
rect 160053 47891 160119 47892
rect 168885 47891 168951 47894
rect 181806 47892 181812 47956
rect 181876 47954 181923 47956
rect 181876 47952 181968 47954
rect 181918 47896 181968 47952
rect 181876 47894 181968 47896
rect 181876 47892 181923 47894
rect 181857 47891 181923 47892
rect 166401 47818 166467 47821
rect 167229 47818 167295 47821
rect 166401 47816 167295 47818
rect 166401 47760 166406 47816
rect 166462 47760 167234 47816
rect 167290 47760 167295 47816
rect 166401 47758 167295 47760
rect 166401 47755 166467 47758
rect 167229 47755 167295 47758
rect 233469 47818 233535 47821
rect 237014 47818 237074 48264
rect 238621 48092 238687 48093
rect 238621 48088 238668 48092
rect 238732 48090 238738 48092
rect 260425 48090 260491 48093
rect 261846 48090 261852 48092
rect 238621 48032 238626 48088
rect 238621 48028 238668 48032
rect 238732 48030 238778 48090
rect 260425 48088 261852 48090
rect 260425 48032 260430 48088
rect 260486 48032 261852 48088
rect 260425 48030 261852 48032
rect 238732 48028 238738 48030
rect 238621 48027 238687 48028
rect 260425 48027 260491 48030
rect 261846 48028 261852 48030
rect 261916 48028 261922 48092
rect 262398 48028 262404 48092
rect 262468 48090 262474 48092
rect 262817 48090 262883 48093
rect 262468 48088 262883 48090
rect 262468 48032 262822 48088
rect 262878 48032 262883 48088
rect 262468 48030 262883 48032
rect 262468 48028 262474 48030
rect 262817 48027 262883 48030
rect 264238 48028 264244 48092
rect 264308 48090 264314 48092
rect 283701 48090 283767 48093
rect 284345 48090 284411 48093
rect 264308 48088 284411 48090
rect 264308 48032 283706 48088
rect 283762 48032 284350 48088
rect 284406 48032 284411 48088
rect 264308 48030 284411 48032
rect 264308 48028 264314 48030
rect 283701 48027 283767 48030
rect 284345 48027 284411 48030
rect 250489 47956 250555 47957
rect 250438 47892 250444 47956
rect 250508 47954 250555 47956
rect 257297 47954 257363 47957
rect 261110 47954 261116 47956
rect 250508 47952 250600 47954
rect 250550 47896 250600 47952
rect 250508 47894 250600 47896
rect 257297 47952 261116 47954
rect 257297 47896 257302 47952
rect 257358 47896 261116 47952
rect 257297 47894 261116 47896
rect 250508 47892 250555 47894
rect 250489 47891 250555 47892
rect 257297 47891 257363 47894
rect 261110 47892 261116 47894
rect 261180 47954 261186 47956
rect 261662 47954 261668 47956
rect 261180 47894 261668 47954
rect 261180 47892 261186 47894
rect 261662 47892 261668 47894
rect 261732 47892 261738 47956
rect 275789 47954 275855 47957
rect 276065 47956 276131 47957
rect 276014 47954 276020 47956
rect 275789 47952 276020 47954
rect 276084 47952 276131 47956
rect 275789 47896 275794 47952
rect 275850 47896 276020 47952
rect 276126 47896 276131 47952
rect 275789 47894 276020 47896
rect 275789 47891 275855 47894
rect 276014 47892 276020 47894
rect 276084 47892 276131 47896
rect 276065 47891 276131 47892
rect 327861 47954 327927 47957
rect 331038 47954 331098 48264
rect 327861 47952 331098 47954
rect 327861 47896 327866 47952
rect 327922 47896 331098 47952
rect 327861 47894 331098 47896
rect 327861 47891 327927 47894
rect 233469 47816 237074 47818
rect 233469 47760 233474 47816
rect 233530 47760 237074 47816
rect 233469 47758 237074 47760
rect 233469 47755 233535 47758
rect 167689 47546 167755 47549
rect 358497 47548 358563 47549
rect 168006 47546 168012 47548
rect 167689 47544 168012 47546
rect 167689 47488 167694 47544
rect 167750 47488 168012 47544
rect 167689 47486 168012 47488
rect 167689 47483 167755 47486
rect 168006 47484 168012 47486
rect 168076 47484 168082 47548
rect 358446 47484 358452 47548
rect 358516 47546 358563 47548
rect 358516 47544 358608 47546
rect 358558 47488 358608 47544
rect 358516 47486 358608 47488
rect 358516 47484 358563 47486
rect 358497 47483 358563 47484
rect 71457 47410 71523 47413
rect 72878 47410 72884 47412
rect 71457 47408 72884 47410
rect 71457 47352 71462 47408
rect 71518 47352 72884 47408
rect 71457 47350 72884 47352
rect 71457 47347 71523 47350
rect 72878 47348 72884 47350
rect 72948 47410 72954 47412
rect 73113 47410 73179 47413
rect 72948 47408 73179 47410
rect 72948 47352 73118 47408
rect 73174 47352 73179 47408
rect 72948 47350 73179 47352
rect 72948 47348 72954 47350
rect 73113 47347 73179 47350
rect 106601 47410 106667 47413
rect 212585 47412 212651 47413
rect 107470 47410 107476 47412
rect 106601 47408 107476 47410
rect 106601 47352 106606 47408
rect 106662 47352 107476 47408
rect 106601 47350 107476 47352
rect 106601 47347 106667 47350
rect 107470 47348 107476 47350
rect 107540 47348 107546 47412
rect 212534 47348 212540 47412
rect 212604 47410 212651 47412
rect 212604 47408 212696 47410
rect 212646 47352 212696 47408
rect 212604 47350 212696 47352
rect 212604 47348 212651 47350
rect 263870 47348 263876 47412
rect 263940 47410 263946 47412
rect 286001 47410 286067 47413
rect 306609 47412 306675 47413
rect 263940 47408 286067 47410
rect 263940 47352 286006 47408
rect 286062 47352 286067 47408
rect 263940 47350 286067 47352
rect 263940 47348 263946 47350
rect 212585 47347 212651 47348
rect 286001 47347 286067 47350
rect 306558 47348 306564 47412
rect 306628 47410 306675 47412
rect 306628 47408 306720 47410
rect 306670 47352 306720 47408
rect 306628 47350 306720 47352
rect 306628 47348 306675 47350
rect 306609 47347 306675 47348
rect 109310 47212 109316 47276
rect 109380 47274 109386 47276
rect 109453 47274 109519 47277
rect 110414 47274 110420 47276
rect 109380 47272 110420 47274
rect 109380 47216 109458 47272
rect 109514 47216 110420 47272
rect 109380 47214 110420 47216
rect 109380 47212 109386 47214
rect 109453 47211 109519 47214
rect 110414 47212 110420 47214
rect 110484 47212 110490 47276
rect 248005 47274 248071 47277
rect 248598 47274 248604 47276
rect 248005 47272 248604 47274
rect 248005 47216 248010 47272
rect 248066 47216 248604 47272
rect 248005 47214 248604 47216
rect 248005 47211 248071 47214
rect 248598 47212 248604 47214
rect 248668 47212 248674 47276
rect 181806 46668 181812 46732
rect 181876 46730 181882 46732
rect 182133 46730 182199 46733
rect 199061 46730 199127 46733
rect 181876 46728 199127 46730
rect 181876 46672 182138 46728
rect 182194 46672 199066 46728
rect 199122 46672 199127 46728
rect 181876 46670 199127 46672
rect 181876 46668 181882 46670
rect 182133 46667 182199 46670
rect 199061 46667 199127 46670
rect 162854 46532 162860 46596
rect 162924 46594 162930 46596
rect 162997 46594 163063 46597
rect 162924 46592 163063 46594
rect 162924 46536 163002 46592
rect 163058 46536 163063 46592
rect 162924 46534 163063 46536
rect 162924 46532 162930 46534
rect 162997 46531 163063 46534
rect 275830 46532 275836 46596
rect 275900 46594 275906 46596
rect 275973 46594 276039 46597
rect 275900 46592 276039 46594
rect 275900 46536 275978 46592
rect 276034 46536 276039 46592
rect 275900 46534 276039 46536
rect 275900 46532 275906 46534
rect 275973 46531 276039 46534
rect 74217 46188 74283 46189
rect 74166 46124 74172 46188
rect 74236 46186 74283 46188
rect 118653 46188 118719 46189
rect 118653 46186 118700 46188
rect 74236 46184 74328 46186
rect 74278 46128 74328 46184
rect 74236 46126 74328 46128
rect 118608 46184 118700 46186
rect 118608 46128 118658 46184
rect 118608 46126 118700 46128
rect 74236 46124 74283 46126
rect 74217 46123 74283 46124
rect 118653 46124 118700 46126
rect 118764 46124 118770 46188
rect 118653 46123 118719 46124
rect 158990 45988 158996 46052
rect 159060 46050 159066 46052
rect 169529 46050 169595 46053
rect 169713 46052 169779 46053
rect 159060 46048 169595 46050
rect 159060 45992 169534 46048
rect 169590 45992 169595 46048
rect 159060 45990 169595 45992
rect 159060 45988 159066 45990
rect 169529 45987 169595 45990
rect 169662 45988 169668 46052
rect 169732 46050 169779 46052
rect 244877 46050 244943 46053
rect 262541 46052 262607 46053
rect 248966 46050 248972 46052
rect 169732 46048 169824 46050
rect 169774 45992 169824 46048
rect 169732 45990 169824 45992
rect 244877 46048 248972 46050
rect 244877 45992 244882 46048
rect 244938 45992 248972 46048
rect 244877 45990 248972 45992
rect 169732 45988 169779 45990
rect 169713 45987 169779 45988
rect 244877 45987 244943 45990
rect 248966 45988 248972 45990
rect 249036 45988 249042 46052
rect 262541 46048 262588 46052
rect 262652 46050 262658 46052
rect 262541 45992 262546 46048
rect 262541 45988 262588 45992
rect 262652 45990 262698 46050
rect 262652 45988 262658 45990
rect 336366 45988 336372 46052
rect 336436 46050 336442 46052
rect 343133 46050 343199 46053
rect 336436 46048 343199 46050
rect 336436 45992 343138 46048
rect 343194 45992 343199 46048
rect 336436 45990 343199 45992
rect 336436 45988 336442 45990
rect 262541 45987 262607 45988
rect 343133 45987 343199 45990
rect 64189 45914 64255 45917
rect 74534 45914 74540 45916
rect 64189 45912 74540 45914
rect 64189 45856 64194 45912
rect 64250 45856 74540 45912
rect 64189 45854 74540 45856
rect 64189 45851 64255 45854
rect 74534 45852 74540 45854
rect 74604 45852 74610 45916
rect 157518 45852 157524 45916
rect 157588 45914 157594 45916
rect 165941 45914 166007 45917
rect 157588 45912 166007 45914
rect 157588 45856 165946 45912
rect 166002 45856 166007 45912
rect 157588 45854 166007 45856
rect 157588 45852 157594 45854
rect 165941 45851 166007 45854
rect 252830 45852 252836 45916
rect 252900 45914 252906 45916
rect 262817 45914 262883 45917
rect 252900 45912 262883 45914
rect 252900 45856 262822 45912
rect 262878 45856 262883 45912
rect 252900 45854 262883 45856
rect 252900 45852 252906 45854
rect 262817 45851 262883 45854
rect 147950 45716 147956 45780
rect 148020 45778 148026 45780
rect 162997 45778 163063 45781
rect 148020 45776 163063 45778
rect 148020 45720 163002 45776
rect 163058 45720 163063 45776
rect 148020 45718 163063 45720
rect 148020 45716 148026 45718
rect 162997 45715 163063 45718
rect 181949 45370 182015 45373
rect 204254 45370 204260 45372
rect 181949 45368 204260 45370
rect 181949 45312 181954 45368
rect 182010 45312 204260 45368
rect 181949 45310 204260 45312
rect 181949 45307 182015 45310
rect 204254 45308 204260 45310
rect 204324 45308 204330 45372
rect 113593 43330 113659 43333
rect 113910 43330 113916 43332
rect 113593 43328 113916 43330
rect 113593 43272 113598 43328
rect 113654 43272 113916 43328
rect 113593 43270 113916 43272
rect 113593 43267 113659 43270
rect 113910 43268 113916 43270
rect 113980 43268 113986 43332
rect 9896 42242 10376 42272
rect 12853 42242 12919 42245
rect 9896 42240 12919 42242
rect 9896 42184 12858 42240
rect 12914 42184 12919 42240
rect 9896 42182 12919 42184
rect 9896 42152 10376 42182
rect 12853 42179 12919 42182
rect 428693 40202 428759 40205
rect 434416 40202 434896 40232
rect 428693 40200 434896 40202
rect 428693 40144 428698 40200
rect 428754 40144 434896 40200
rect 428693 40142 434896 40144
rect 428693 40139 428759 40142
rect 434416 40112 434896 40142
rect 207525 37754 207591 37757
rect 301549 37756 301615 37757
rect 207750 37754 207756 37756
rect 207525 37752 207756 37754
rect 207525 37696 207530 37752
rect 207586 37696 207756 37752
rect 207525 37694 207756 37696
rect 207525 37691 207591 37694
rect 207750 37692 207756 37694
rect 207820 37692 207826 37756
rect 301549 37754 301596 37756
rect 301504 37752 301596 37754
rect 301504 37696 301554 37752
rect 301504 37694 301596 37696
rect 301549 37692 301596 37694
rect 301660 37692 301666 37756
rect 301549 37691 301615 37692
rect 88109 33674 88175 33677
rect 181949 33674 182015 33677
rect 275881 33674 275947 33677
rect 88109 33672 90058 33674
rect 88109 33616 88114 33672
rect 88170 33616 90058 33672
rect 88109 33614 90058 33616
rect 88109 33611 88175 33614
rect 89998 33444 90058 33614
rect 181949 33672 184082 33674
rect 181949 33616 181954 33672
rect 182010 33616 184082 33672
rect 181949 33614 184082 33616
rect 181949 33611 182015 33614
rect 184022 33444 184082 33614
rect 275881 33672 278106 33674
rect 275881 33616 275886 33672
rect 275942 33616 278106 33672
rect 275881 33614 278106 33616
rect 275881 33611 275947 33614
rect 278046 33444 278106 33614
rect 88201 30818 88267 30821
rect 182041 30818 182107 30821
rect 275973 30818 276039 30821
rect 88201 30816 90058 30818
rect 88201 30760 88206 30816
rect 88262 30760 90058 30816
rect 88201 30758 90058 30760
rect 88201 30755 88267 30758
rect 89998 30724 90058 30758
rect 182041 30816 184082 30818
rect 182041 30760 182046 30816
rect 182102 30760 184082 30816
rect 182041 30758 184082 30760
rect 182041 30755 182107 30758
rect 184022 30724 184082 30758
rect 275973 30816 278106 30818
rect 275973 30760 275978 30816
rect 276034 30760 278106 30816
rect 275973 30758 278106 30760
rect 275973 30755 276039 30758
rect 278046 30724 278106 30758
rect 9896 28914 10376 28944
rect 12669 28914 12735 28917
rect 9896 28912 12735 28914
rect 9896 28856 12674 28912
rect 12730 28856 12735 28912
rect 9896 28854 12735 28856
rect 9896 28824 10376 28854
rect 12669 28851 12735 28854
rect 88293 28098 88359 28101
rect 89998 28098 90058 28136
rect 88293 28096 90058 28098
rect 88293 28040 88298 28096
rect 88354 28040 90058 28096
rect 88293 28038 90058 28040
rect 182133 28098 182199 28101
rect 184022 28098 184082 28136
rect 182133 28096 184082 28098
rect 182133 28040 182138 28096
rect 182194 28040 184082 28096
rect 182133 28038 184082 28040
rect 275789 28098 275855 28101
rect 278046 28098 278106 28136
rect 275789 28096 278106 28098
rect 275789 28040 275794 28096
rect 275850 28040 278106 28096
rect 275789 28038 278106 28040
rect 88293 28035 88359 28038
rect 182133 28035 182199 28038
rect 275789 28035 275855 28038
rect 429797 27690 429863 27693
rect 434416 27690 434896 27720
rect 429797 27688 434896 27690
rect 429797 27632 429802 27688
rect 429858 27632 434896 27688
rect 429797 27630 434896 27632
rect 429797 27627 429863 27630
rect 434416 27600 434896 27630
rect 88385 26058 88451 26061
rect 182225 26058 182291 26061
rect 276065 26058 276131 26061
rect 88385 26056 90058 26058
rect 88385 26000 88390 26056
rect 88446 26000 90058 26056
rect 88385 25998 90058 26000
rect 88385 25995 88451 25998
rect 89998 25420 90058 25998
rect 182225 26056 184082 26058
rect 182225 26000 182230 26056
rect 182286 26000 184082 26056
rect 182225 25998 184082 26000
rect 182225 25995 182291 25998
rect 184022 25420 184082 25998
rect 276065 26056 278106 26058
rect 276065 26000 276070 26056
rect 276126 26000 278106 26056
rect 276065 25998 278106 26000
rect 276065 25995 276131 25998
rect 278046 25420 278106 25998
rect 88017 23338 88083 23341
rect 181857 23338 181923 23341
rect 275513 23338 275579 23341
rect 88017 23336 90058 23338
rect 88017 23280 88022 23336
rect 88078 23280 90058 23336
rect 88017 23278 90058 23280
rect 88017 23275 88083 23278
rect 89998 22700 90058 23278
rect 181857 23336 184082 23338
rect 181857 23280 181862 23336
rect 181918 23280 184082 23336
rect 181857 23278 184082 23280
rect 181857 23275 181923 23278
rect 184022 22700 184082 23278
rect 275513 23336 278106 23338
rect 275513 23280 275518 23336
rect 275574 23280 278106 23336
rect 275513 23278 278106 23280
rect 275513 23275 275579 23278
rect 278046 22700 278106 23278
rect 88477 20754 88543 20757
rect 182317 20754 182383 20757
rect 276157 20754 276223 20757
rect 88477 20752 90058 20754
rect 88477 20696 88482 20752
rect 88538 20696 90058 20752
rect 88477 20694 90058 20696
rect 88477 20691 88543 20694
rect 89998 20116 90058 20694
rect 182317 20752 184082 20754
rect 182317 20696 182322 20752
rect 182378 20696 184082 20752
rect 182317 20694 184082 20696
rect 182317 20691 182383 20694
rect 184022 20116 184082 20694
rect 276157 20752 278106 20754
rect 276157 20696 276162 20752
rect 276218 20696 278106 20752
rect 276157 20694 278106 20696
rect 276157 20691 276223 20694
rect 278046 20116 278106 20694
rect 9896 15586 10376 15616
rect 13037 15586 13103 15589
rect 9896 15584 13103 15586
rect 9896 15528 13042 15584
rect 13098 15528 13103 15584
rect 9896 15526 13103 15528
rect 9896 15496 10376 15526
rect 13037 15523 13103 15526
rect 429429 15178 429495 15181
rect 434416 15178 434896 15208
rect 429429 15176 434896 15178
rect 429429 15120 429434 15176
rect 429490 15120 434896 15176
rect 429429 15118 434896 15120
rect 429429 15115 429495 15118
rect 434416 15088 434896 15118
<< via3 >>
rect 280252 393740 280316 393804
rect 323124 393740 323188 393804
rect 323492 393060 323556 393124
rect 97356 367220 97420 367284
rect 285036 367220 285100 367284
rect 97356 352048 97420 352052
rect 97356 351992 97370 352048
rect 97370 351992 97420 352048
rect 97356 351988 97420 351992
rect 285036 351640 285100 351644
rect 285036 351584 285050 351640
rect 285050 351584 285100 351640
rect 285036 351580 285100 351584
rect 104900 333764 104964 333828
rect 212172 333492 212236 333556
rect 231860 333552 231924 333556
rect 231860 333496 231874 333552
rect 231874 333496 231924 333552
rect 231860 333492 231924 333496
rect 306196 333552 306260 333556
rect 306196 333496 306246 333552
rect 306246 333496 306260 333552
rect 306196 333492 306260 333496
rect 280252 333084 280316 333148
rect 137284 332132 137348 332196
rect 198740 332192 198804 332196
rect 198740 332136 198790 332192
rect 198790 332136 198804 332192
rect 198740 332132 198804 332136
rect 231860 332132 231924 332196
rect 296076 332132 296140 332196
rect 137284 331452 137348 331516
rect 204444 331588 204508 331652
rect 294052 331588 294116 331652
rect 231860 331452 231924 331516
rect 159548 330152 159612 330156
rect 159548 330096 159598 330152
rect 159598 330096 159612 330152
rect 159548 330092 159612 330096
rect 252284 330092 252348 330156
rect 251548 329956 251612 330020
rect 253020 329956 253084 330020
rect 161756 329472 161820 329476
rect 161756 329416 161770 329472
rect 161770 329416 161820 329472
rect 161756 329412 161820 329416
rect 262404 327508 262468 327572
rect 52644 327372 52708 327436
rect 54668 327372 54732 327436
rect 55404 327372 55468 327436
rect 168564 327372 168628 327436
rect 339500 327372 339564 327436
rect 340972 327372 341036 327436
rect 153292 326344 153356 326348
rect 153292 326288 153306 326344
rect 153306 326288 153356 326344
rect 153292 326284 153356 326288
rect 55220 317852 55284 317916
rect 55404 315812 55468 315876
rect 153292 315812 153356 315876
rect 340972 314860 341036 314924
rect 351828 314860 351892 314924
rect 339500 314588 339564 314652
rect 352564 314452 352628 314516
rect 55036 310372 55100 310436
rect 54668 306156 54732 306220
rect 74540 305612 74604 305676
rect 73988 303980 74052 304044
rect 52644 300580 52708 300644
rect 73804 300036 73868 300100
rect 134708 298132 134772 298196
rect 323492 295412 323556 295476
rect 136916 294732 136980 294796
rect 228732 294732 228796 294796
rect 231860 294596 231924 294660
rect 74172 292964 74236 293028
rect 136916 292148 136980 292212
rect 230756 292012 230820 292076
rect 322756 291876 322820 291940
rect 73436 291740 73500 291804
rect 73988 291740 74052 291804
rect 261116 290652 261180 290716
rect 270500 290652 270564 290716
rect 138020 289292 138084 289356
rect 228732 289292 228796 289356
rect 323124 289020 323188 289084
rect 73436 286300 73500 286364
rect 74172 286300 74236 286364
rect 353668 285212 353732 285276
rect 84660 284940 84724 285004
rect 134892 284804 134956 284868
rect 73620 282764 73684 282828
rect 84476 282764 84540 282828
rect 73436 281948 73500 282012
rect 74172 281948 74236 282012
rect 352748 279636 352812 279700
rect 138388 279364 138452 279428
rect 138388 279288 138452 279292
rect 138388 279232 138438 279288
rect 138438 279232 138452 279288
rect 138388 279228 138452 279232
rect 73436 277324 73500 277388
rect 73436 277188 73500 277252
rect 73988 277188 74052 277252
rect 73988 277052 74052 277116
rect 149060 274876 149124 274940
rect 168932 274740 168996 274804
rect 262036 274740 262100 274804
rect 168564 274604 168628 274668
rect 262404 274604 262468 274668
rect 167828 274468 167892 274532
rect 262588 274468 262652 274532
rect 168196 274332 168260 274396
rect 261668 274332 261732 274396
rect 247868 273984 247932 273988
rect 247868 273928 247882 273984
rect 247882 273928 247932 273984
rect 247868 273924 247932 273928
rect 136916 273788 136980 273852
rect 154580 273788 154644 273852
rect 242348 273788 242412 273852
rect 74172 271128 74236 271132
rect 74172 271072 74222 271128
rect 74222 271072 74236 271128
rect 74172 271068 74236 271072
rect 73988 270388 74052 270452
rect 73436 270252 73500 270316
rect 73988 270252 74052 270316
rect 73436 270116 73500 270180
rect 138572 269844 138636 269908
rect 138572 269572 138636 269636
rect 138756 269572 138820 269636
rect 182916 269496 182980 269500
rect 182916 269440 182966 269496
rect 182966 269440 182980 269496
rect 182916 269436 182980 269440
rect 219716 268348 219780 268412
rect 351828 266716 351892 266780
rect 55220 266580 55284 266644
rect 352012 266580 352076 266644
rect 52644 265492 52708 265556
rect 54668 265492 54732 265556
rect 55404 265492 55468 265556
rect 241428 263860 241492 263924
rect 242716 263860 242780 263924
rect 73804 263588 73868 263652
rect 75460 263588 75524 263652
rect 74540 263452 74604 263516
rect 73436 263316 73500 263380
rect 74724 263316 74788 263380
rect 245108 263452 245172 263516
rect 251180 263452 251244 263516
rect 183836 262092 183900 262156
rect 193220 262092 193284 262156
rect 278964 261412 279028 261476
rect 288532 261412 288596 261476
rect 298284 261412 298348 261476
rect 307852 261412 307916 261476
rect 317604 261412 317668 261476
rect 327172 261412 327236 261476
rect 203156 260732 203220 260796
rect 212540 260732 212604 260796
rect 138756 259976 138820 259980
rect 138756 259920 138806 259976
rect 138806 259920 138820 259976
rect 138756 259916 138820 259920
rect 48964 259372 49028 259436
rect 48964 255836 49028 255900
rect 138756 250396 138820 250460
rect 48964 249172 49028 249236
rect 49148 246044 49212 246108
rect 138756 245500 138820 245564
rect 46940 243460 47004 243524
rect 96068 241692 96132 241756
rect 104900 241692 104964 241756
rect 84476 241012 84540 241076
rect 93860 241012 93924 241076
rect 138388 240740 138452 240804
rect 196164 240332 196228 240396
rect 305092 240392 305156 240396
rect 305092 240336 305142 240392
rect 305142 240336 305156 240392
rect 305092 240332 305156 240336
rect 49148 239788 49212 239852
rect 295524 239788 295588 239852
rect 95148 239712 95212 239716
rect 95148 239656 95198 239712
rect 95198 239656 95212 239712
rect 95148 239652 95212 239656
rect 187884 239652 187948 239716
rect 324596 239652 324660 239716
rect 92572 239380 92636 239444
rect 192116 239380 192180 239444
rect 283196 239440 283260 239444
rect 283196 239384 283246 239440
rect 283246 239384 283260 239440
rect 283196 239380 283260 239384
rect 198924 238428 198988 238492
rect 290004 238488 290068 238492
rect 290004 238432 290054 238488
rect 290054 238432 290068 238488
rect 290004 238428 290068 238432
rect 100116 237884 100180 237948
rect 231860 237884 231924 237948
rect 219716 237808 219780 237812
rect 219716 237752 219766 237808
rect 219766 237752 219780 237808
rect 219716 237748 219780 237752
rect 141148 237612 141212 237676
rect 143172 237612 143236 237676
rect 89996 236932 90060 236996
rect 100116 236932 100180 236996
rect 186596 236932 186660 236996
rect 198924 236932 198988 236996
rect 264796 236932 264860 236996
rect 273812 236932 273876 236996
rect 74540 236388 74604 236452
rect 75460 236388 75524 236452
rect 81348 236388 81412 236452
rect 73436 236252 73500 236316
rect 74724 236252 74788 236316
rect 76380 236252 76444 236316
rect 203156 236312 203220 236316
rect 203156 236256 203170 236312
rect 203170 236256 203220 236312
rect 203156 236252 203220 236256
rect 286876 236312 286940 236316
rect 286876 236256 286926 236312
rect 286926 236256 286940 236312
rect 286876 236252 286940 236256
rect 73988 236116 74052 236180
rect 76564 236116 76628 236180
rect 167828 236116 167892 236180
rect 177028 236116 177092 236180
rect 244188 236176 244252 236180
rect 244188 236120 244238 236176
rect 244238 236120 244252 236176
rect 244188 236116 244252 236120
rect 73620 235980 73684 236044
rect 76012 235980 76076 236044
rect 147772 235980 147836 236044
rect 168196 235980 168260 236044
rect 75644 235844 75708 235908
rect 76932 235844 76996 235908
rect 116124 235844 116188 235908
rect 148692 235844 148756 235908
rect 247132 235844 247196 235908
rect 105084 235708 105148 235772
rect 167828 235708 167892 235772
rect 262588 235768 262652 235772
rect 262588 235712 262602 235768
rect 262602 235712 262652 235768
rect 262588 235708 262652 235712
rect 74356 235572 74420 235636
rect 74908 235572 74972 235636
rect 124404 235572 124468 235636
rect 133972 235572 134036 235636
rect 152004 235632 152068 235636
rect 152004 235576 152008 235632
rect 152008 235576 152064 235632
rect 152064 235576 152068 235632
rect 152004 235572 152068 235576
rect 158812 235572 158876 235636
rect 246212 235572 246276 235636
rect 74540 235436 74604 235500
rect 75460 235436 75524 235500
rect 145196 235360 145260 235364
rect 145196 235304 145210 235360
rect 145210 235304 145260 235360
rect 145196 235300 145260 235304
rect 75276 235028 75340 235092
rect 136364 235028 136428 235092
rect 137284 234892 137348 234956
rect 148140 234952 148204 234956
rect 148140 234896 148190 234952
rect 148190 234896 148204 234952
rect 148140 234892 148204 234896
rect 231308 234892 231372 234956
rect 245476 234892 245540 234956
rect 301044 234952 301108 234956
rect 301044 234896 301094 234952
rect 301094 234896 301108 234952
rect 301044 234892 301108 234896
rect 207204 234408 207268 234412
rect 207204 234352 207254 234408
rect 207254 234352 207268 234408
rect 207204 234348 207268 234352
rect 283196 234348 283260 234412
rect 137652 234212 137716 234276
rect 73804 234076 73868 234140
rect 75644 234076 75708 234140
rect 230756 234136 230820 234140
rect 230756 234080 230770 234136
rect 230770 234080 230820 234136
rect 230756 234076 230820 234080
rect 74172 233804 74236 233868
rect 74908 233804 74972 233868
rect 74908 233668 74972 233732
rect 156788 233668 156852 233732
rect 261668 233668 261732 233732
rect 249892 233396 249956 233460
rect 262036 233260 262100 233324
rect 52644 232444 52708 232508
rect 54668 232444 54732 232508
rect 55588 232504 55652 232508
rect 55588 232448 55602 232504
rect 55602 232448 55652 232504
rect 55588 232444 55652 232448
rect 239588 232444 239652 232508
rect 351644 232444 351708 232508
rect 351828 232444 351892 232508
rect 185860 227004 185924 227068
rect 193036 227004 193100 227068
rect 55404 226868 55468 226932
rect 174084 226868 174148 226932
rect 116124 226732 116188 226796
rect 135444 226732 135508 226796
rect 154764 226596 154828 226660
rect 185860 226596 185924 226660
rect 92572 226460 92636 226524
rect 109132 226460 109196 226524
rect 109500 226460 109564 226524
rect 116124 226460 116188 226524
rect 135444 226460 135508 226524
rect 154764 226324 154828 226388
rect 174084 226460 174148 226524
rect 178684 226460 178748 226524
rect 182916 226460 182980 226524
rect 193220 226460 193284 226524
rect 73804 224284 73868 224348
rect 73804 224148 73868 224212
rect 74540 224148 74604 224212
rect 73804 224012 73868 224076
rect 74540 224012 74604 224076
rect 73804 223876 73868 223940
rect 55404 221972 55468 222036
rect 55588 221292 55652 221356
rect 56324 221292 56388 221356
rect 242716 216532 242780 216596
rect 258908 216532 258972 216596
rect 272708 216532 272772 216596
rect 322756 216532 322820 216596
rect 336740 216532 336804 216596
rect 352748 216532 352812 216596
rect 358268 216396 358332 216460
rect 357532 215852 357596 215916
rect 405924 215852 405988 215916
rect 73436 213676 73500 213740
rect 54668 210956 54732 211020
rect 147036 208236 147100 208300
rect 52644 206740 52708 206804
rect 73804 205032 73868 205036
rect 73804 204976 73854 205032
rect 73854 204976 73868 205032
rect 73804 204972 73868 204976
rect 73804 204836 73868 204900
rect 74540 204836 74604 204900
rect 134708 204836 134772 204900
rect 72148 204700 72212 204764
rect 73988 204700 74052 204764
rect 74540 204700 74604 204764
rect 73620 204428 73684 204492
rect 84660 204428 84724 204492
rect 242716 204564 242780 204628
rect 237380 204292 237444 204356
rect 239588 204292 239652 204356
rect 322756 204156 322820 204220
rect 73620 203476 73684 203540
rect 73620 202116 73684 202180
rect 74356 202116 74420 202180
rect 242716 201980 242780 202044
rect 136916 200892 136980 200956
rect 228732 200892 228796 200956
rect 322756 200892 322820 200956
rect 74540 199124 74604 199188
rect 164884 198852 164948 198916
rect 176660 198852 176724 198916
rect 322756 198716 322820 198780
rect 136916 198172 136980 198236
rect 230756 197552 230820 197556
rect 230756 197496 230770 197552
rect 230770 197496 230820 197552
rect 230756 197492 230820 197496
rect 261116 197492 261180 197556
rect 270500 197492 270564 197556
rect 74172 195240 74236 195244
rect 74172 195184 74222 195240
rect 74222 195184 74236 195240
rect 74172 195180 74236 195184
rect 74540 195240 74604 195244
rect 74540 195184 74554 195240
rect 74554 195184 74604 195240
rect 74540 195180 74604 195184
rect 74356 195044 74420 195108
rect 74540 195104 74604 195108
rect 74540 195048 74554 195104
rect 74554 195048 74604 195104
rect 74540 195044 74604 195048
rect 230756 194908 230820 194972
rect 138020 194636 138084 194700
rect 322756 194500 322820 194564
rect 72332 192596 72396 192660
rect 72700 192460 72764 192524
rect 242532 192520 242596 192524
rect 242532 192464 242582 192520
rect 242582 192464 242596 192520
rect 242532 192460 242596 192464
rect 352748 191432 352812 191436
rect 352748 191376 352798 191432
rect 352798 191376 352812 191432
rect 352748 191372 352812 191376
rect 73988 191236 74052 191300
rect 74540 185660 74604 185724
rect 73988 185584 74052 185588
rect 73988 185528 74002 185584
rect 74002 185528 74052 185584
rect 73988 185524 74052 185528
rect 74540 185524 74604 185588
rect 73988 185448 74052 185452
rect 73988 185392 74002 185448
rect 74002 185392 74052 185448
rect 73988 185388 74052 185392
rect 71964 185252 72028 185316
rect 72700 185252 72764 185316
rect 351644 184028 351708 184092
rect 242716 183076 242780 183140
rect 271420 182124 271484 182188
rect 322940 182124 323004 182188
rect 174820 181988 174884 182052
rect 228916 181988 228980 182052
rect 271420 181988 271484 182052
rect 322940 181988 323004 182052
rect 147036 181172 147100 181236
rect 169116 181036 169180 181100
rect 168564 180900 168628 180964
rect 167644 180764 167708 180828
rect 261668 180764 261732 180828
rect 169484 180628 169548 180692
rect 242348 180628 242412 180692
rect 262404 180628 262468 180692
rect 147956 180492 148020 180556
rect 167828 180492 167892 180556
rect 262956 180492 263020 180556
rect 241796 180084 241860 180148
rect 242900 179948 242964 180012
rect 287428 179268 287492 179332
rect 289452 179268 289516 179332
rect 310980 179268 311044 179332
rect 317052 179268 317116 179332
rect 286140 179132 286204 179196
rect 288532 179132 288596 179196
rect 309876 179132 309940 179196
rect 311900 179132 311964 179196
rect 178316 178240 178380 178244
rect 178316 178184 178330 178240
rect 178330 178184 178380 178240
rect 178316 178180 178380 178184
rect 73620 177908 73684 177972
rect 75460 177908 75524 177972
rect 71964 176412 72028 176476
rect 71964 175868 72028 175932
rect 72332 175868 72396 175932
rect 182916 175792 182980 175796
rect 182916 175736 182930 175792
rect 182930 175736 182980 175792
rect 182916 175732 182980 175736
rect 219716 175460 219780 175524
rect 74172 173692 74236 173756
rect 52644 172876 52708 172940
rect 54668 172876 54732 172940
rect 55588 172936 55652 172940
rect 55588 172880 55602 172936
rect 55602 172880 55652 172936
rect 55588 172876 55652 172880
rect 55404 172740 55468 172804
rect 351644 172604 351708 172668
rect 351828 172604 351892 172668
rect 75460 169748 75524 169812
rect 76748 169748 76812 169812
rect 74172 169612 74236 169676
rect 76380 169612 76444 169676
rect 73436 169476 73500 169540
rect 73804 169476 73868 169540
rect 75460 169476 75524 169540
rect 74724 169340 74788 169404
rect 75644 169340 75708 169404
rect 72332 169204 72396 169268
rect 75828 169204 75892 169268
rect 144092 169204 144156 169268
rect 147956 169204 148020 169268
rect 237012 167028 237076 167092
rect 48964 162540 49028 162604
rect 49148 158324 49212 158388
rect 76564 157508 76628 157572
rect 76748 157100 76812 157164
rect 49148 155332 49212 155396
rect 49148 152884 49212 152948
rect 49148 148940 49212 149004
rect 76564 148532 76628 148596
rect 236828 147852 236892 147916
rect 237196 147852 237260 147916
rect 49148 145812 49212 145876
rect 76564 145812 76628 145876
rect 176292 145132 176356 145196
rect 187148 145132 187212 145196
rect 197636 144588 197700 144652
rect 196164 144452 196228 144516
rect 290004 144452 290068 144516
rect 98276 144180 98340 144244
rect 142252 144180 142316 144244
rect 76932 144104 76996 144108
rect 76932 144048 76982 144104
rect 76982 144048 76996 144104
rect 76932 144044 76996 144048
rect 142068 144044 142132 144108
rect 236092 144044 236156 144108
rect 197636 143968 197700 143972
rect 197636 143912 197686 143968
rect 197686 143912 197700 143968
rect 197636 143908 197700 143912
rect 110420 143228 110484 143292
rect 136916 143228 136980 143292
rect 210148 143092 210212 143156
rect 294236 143152 294300 143156
rect 294236 143096 294286 143152
rect 294286 143096 294300 143152
rect 294236 143092 294300 143096
rect 89628 142820 89692 142884
rect 73804 142412 73868 142476
rect 74356 142412 74420 142476
rect 74908 142412 74972 142476
rect 74540 142140 74604 142204
rect 75644 142140 75708 142204
rect 73988 142004 74052 142068
rect 74540 142004 74604 142068
rect 75276 142004 75340 142068
rect 76012 141868 76076 141932
rect 142436 142276 142500 142340
rect 151820 142276 151884 142340
rect 142252 142140 142316 142204
rect 144092 142140 144156 142204
rect 167644 142140 167708 142204
rect 142068 142004 142132 142068
rect 219716 142064 219780 142068
rect 238300 142412 238364 142476
rect 242532 142412 242596 142476
rect 238116 142140 238180 142204
rect 261668 142140 261732 142204
rect 219716 142008 219730 142064
rect 219730 142008 219780 142064
rect 219716 142004 219780 142008
rect 105084 141868 105148 141932
rect 230756 141868 230820 141932
rect 74356 141732 74420 141796
rect 76932 141732 76996 141796
rect 78220 141732 78284 141796
rect 167828 141732 167892 141796
rect 168380 141732 168444 141796
rect 237748 141732 237812 141796
rect 241980 141732 242044 141796
rect 256700 141732 256764 141796
rect 137468 141052 137532 141116
rect 149060 141112 149124 141116
rect 149060 141056 149110 141112
rect 149110 141056 149124 141112
rect 149060 141052 149124 141056
rect 207204 141112 207268 141116
rect 207204 141056 207254 141112
rect 207254 141056 207268 141112
rect 207204 141052 207268 141056
rect 296996 141052 297060 141116
rect 152004 140432 152068 140436
rect 152004 140376 152054 140432
rect 152054 140376 152068 140432
rect 152004 140372 152068 140376
rect 137284 140296 137348 140300
rect 137284 140240 137298 140296
rect 137298 140240 137348 140296
rect 137284 140236 137348 140240
rect 230756 139964 230820 140028
rect 147772 139828 147836 139892
rect 148508 139828 148572 139892
rect 169116 139828 169180 139892
rect 243084 139828 243148 139892
rect 262956 139828 263020 139892
rect 242532 139692 242596 139756
rect 251364 139692 251428 139756
rect 52644 139556 52708 139620
rect 54852 139556 54916 139620
rect 351644 139556 351708 139620
rect 351828 139556 351892 139620
rect 73436 139420 73500 139484
rect 252652 138468 252716 138532
rect 249708 138392 249772 138396
rect 249708 138336 249722 138392
rect 249722 138336 249772 138392
rect 249708 138332 249772 138336
rect 252652 137788 252716 137852
rect 298100 137788 298164 137852
rect 73620 137108 73684 137172
rect 198556 135068 198620 135132
rect 55220 134388 55284 134452
rect 249156 134448 249220 134452
rect 249156 134392 249170 134448
rect 249170 134392 249220 134448
rect 249156 134388 249220 134392
rect 351828 134252 351892 134316
rect 352564 134116 352628 134180
rect 55404 132348 55468 132412
rect 178684 132484 178748 132548
rect 182916 132484 182980 132548
rect 198556 132484 198620 132548
rect 199292 132484 199356 132548
rect 298100 132484 298164 132548
rect 246212 130172 246276 130236
rect 241980 129552 242044 129556
rect 241980 129496 242030 129552
rect 242030 129496 242044 129552
rect 241980 129492 242044 129496
rect 84660 127512 84724 127516
rect 84660 127456 84710 127512
rect 84710 127456 84724 127512
rect 84660 127452 84724 127456
rect 252652 127452 252716 127516
rect 259644 127452 259708 127516
rect 55404 127180 55468 127244
rect 248604 126772 248668 126836
rect 249708 126772 249772 126836
rect 73252 124732 73316 124796
rect 242164 124732 242228 124796
rect 73252 124596 73316 124660
rect 148692 122284 148756 122348
rect 148876 122148 148940 122212
rect 54668 122012 54732 122076
rect 55036 122012 55100 122076
rect 231860 119292 231924 119356
rect 73804 117660 73868 117724
rect 74356 117660 74420 117724
rect 54852 117116 54916 117180
rect 136916 116572 136980 116636
rect 229284 116572 229348 116636
rect 238852 116572 238916 116636
rect 146668 113232 146732 113236
rect 146668 113176 146682 113232
rect 146682 113176 146732 113232
rect 146668 113172 146732 113176
rect 147772 113172 147836 113236
rect 52644 113036 52708 113100
rect 230756 112900 230820 112964
rect 74540 112764 74604 112828
rect 241980 110180 242044 110244
rect 242532 110180 242596 110244
rect 84660 109832 84724 109836
rect 84660 109776 84710 109832
rect 84710 109776 84724 109832
rect 84660 109772 84724 109776
rect 134708 109772 134772 109836
rect 240140 109832 240204 109836
rect 240140 109776 240154 109832
rect 240154 109776 240204 109832
rect 240140 109772 240204 109776
rect 322756 109772 322820 109836
rect 73804 109500 73868 109564
rect 148692 108820 148756 108884
rect 148876 108820 148940 108884
rect 230756 107928 230820 107932
rect 230756 107872 230806 107928
rect 230806 107872 230820 107928
rect 230756 107868 230820 107872
rect 137468 106780 137532 106844
rect 324596 106780 324660 106844
rect 138020 104332 138084 104396
rect 231860 104332 231924 104396
rect 228732 103924 228796 103988
rect 322756 103924 322820 103988
rect 261116 102972 261180 103036
rect 270500 102972 270564 103036
rect 171324 102292 171388 102356
rect 177028 102292 177092 102356
rect 74172 102020 74236 102084
rect 164884 100660 164948 100724
rect 178684 100660 178748 100724
rect 241980 100720 242044 100724
rect 241980 100664 242030 100720
rect 242030 100664 242044 100720
rect 241980 100660 242044 100664
rect 258724 100660 258788 100724
rect 272708 100660 272772 100724
rect 322756 100388 322820 100452
rect 178684 99980 178748 100044
rect 228732 99980 228796 100044
rect 145748 99844 145812 99908
rect 258724 99980 258788 100044
rect 272708 99980 272772 100044
rect 242716 99844 242780 99908
rect 164884 98680 164948 98684
rect 164884 98624 164934 98680
rect 164934 98624 164948 98680
rect 164884 98620 164948 98624
rect 73620 98212 73684 98276
rect 352748 97864 352812 97868
rect 352748 97808 352798 97864
rect 352798 97808 352812 97864
rect 352748 97804 352812 97808
rect 241980 95824 242044 95828
rect 241980 95768 242030 95824
rect 242030 95768 242044 95824
rect 241980 95764 242044 95768
rect 148876 95492 148940 95556
rect 74540 93860 74604 93924
rect 84660 93452 84724 93516
rect 148876 90052 148940 90116
rect 152188 90052 152252 90116
rect 155500 90052 155564 90116
rect 351644 90052 351708 90116
rect 74172 89780 74236 89844
rect 245844 89100 245908 89164
rect 241980 88964 242044 89028
rect 155500 88888 155564 88892
rect 155500 88832 155514 88888
rect 155514 88832 155564 88888
rect 155500 88828 155564 88832
rect 155684 88888 155748 88892
rect 155684 88832 155734 88888
rect 155734 88832 155748 88888
rect 155684 88828 155748 88832
rect 241980 88828 242044 88892
rect 249524 88828 249588 88892
rect 251732 88616 251796 88620
rect 251732 88560 251736 88616
rect 251736 88560 251792 88616
rect 251792 88560 251796 88616
rect 251732 88556 251796 88560
rect 74172 87468 74236 87532
rect 156052 87332 156116 87396
rect 246212 87468 246276 87532
rect 167644 87332 167708 87396
rect 251180 87332 251244 87396
rect 148508 87196 148572 87260
rect 168748 87060 168812 87124
rect 169300 86924 169364 86988
rect 168012 86788 168076 86852
rect 262404 86788 262468 86852
rect 169116 86652 169180 86716
rect 262588 86652 262652 86716
rect 336372 86652 336436 86716
rect 74540 86380 74604 86444
rect 72884 86244 72948 86308
rect 251180 86244 251244 86308
rect 72700 86108 72764 86172
rect 73988 86108 74052 86172
rect 249892 86108 249956 86172
rect 178684 84264 178748 84268
rect 178684 84208 178734 84264
rect 178734 84208 178748 84264
rect 178684 84204 178748 84208
rect 242164 83388 242228 83452
rect 242900 83388 242964 83452
rect 54852 77948 54916 78012
rect 52644 77812 52708 77876
rect 54668 77812 54732 77876
rect 55404 77812 55468 77876
rect 351644 77812 351708 77876
rect 351828 77812 351892 77876
rect 238668 75364 238732 75428
rect 242900 75364 242964 75428
rect 251180 75364 251244 75428
rect 261852 75364 261916 75428
rect 113916 53120 113980 53124
rect 113916 53064 113966 53120
rect 113966 53064 113980 53120
rect 113916 53060 113980 53064
rect 118700 53120 118764 53124
rect 118700 53064 118714 53120
rect 118714 53064 118764 53120
rect 118700 53060 118764 53064
rect 212540 53120 212604 53124
rect 212540 53064 212554 53120
rect 212554 53064 212604 53120
rect 212540 53060 212604 53064
rect 301596 53120 301660 53124
rect 301596 53064 301646 53120
rect 301646 53064 301660 53120
rect 301596 53060 301660 53064
rect 306564 53120 306628 53124
rect 306564 53064 306614 53120
rect 306614 53064 306628 53120
rect 306564 53060 306628 53064
rect 191380 51564 191444 51628
rect 204260 51564 204324 51628
rect 102508 51292 102572 51356
rect 207756 51292 207820 51356
rect 270684 51292 270748 51356
rect 142436 51020 142500 51084
rect 93676 50672 93740 50676
rect 93676 50616 93690 50672
rect 93690 50616 93740 50672
rect 93676 50612 93740 50616
rect 170588 50672 170652 50676
rect 170588 50616 170602 50672
rect 170602 50616 170652 50672
rect 170588 50612 170652 50616
rect 187148 50612 187212 50676
rect 358452 50340 358516 50404
rect 107476 50264 107540 50268
rect 107476 50208 107526 50264
rect 107526 50208 107540 50264
rect 107476 50204 107540 50208
rect 109316 50204 109380 50268
rect 88340 49312 88404 49316
rect 88340 49256 88390 49312
rect 88390 49256 88404 49312
rect 88340 49252 88404 49256
rect 105268 49252 105332 49316
rect 181996 49252 182060 49316
rect 88156 48572 88220 48636
rect 67916 48088 67980 48092
rect 67916 48032 67930 48088
rect 67930 48032 67980 48088
rect 67916 48028 67980 48032
rect 73988 48028 74052 48092
rect 147956 48028 148020 48092
rect 154764 48028 154828 48092
rect 145564 47892 145628 47956
rect 147956 47892 148020 47956
rect 160100 47952 160164 47956
rect 160100 47896 160114 47952
rect 160114 47896 160164 47952
rect 160100 47892 160164 47896
rect 168748 47892 168812 47956
rect 181812 47952 181876 47956
rect 181812 47896 181862 47952
rect 181862 47896 181876 47952
rect 181812 47892 181876 47896
rect 238668 48088 238732 48092
rect 238668 48032 238682 48088
rect 238682 48032 238732 48088
rect 238668 48028 238732 48032
rect 261852 48028 261916 48092
rect 262404 48028 262468 48092
rect 264244 48028 264308 48092
rect 250444 47952 250508 47956
rect 250444 47896 250494 47952
rect 250494 47896 250508 47952
rect 250444 47892 250508 47896
rect 261116 47892 261180 47956
rect 261668 47892 261732 47956
rect 276020 47952 276084 47956
rect 276020 47896 276070 47952
rect 276070 47896 276084 47952
rect 276020 47892 276084 47896
rect 168012 47484 168076 47548
rect 358452 47544 358516 47548
rect 358452 47488 358502 47544
rect 358502 47488 358516 47544
rect 358452 47484 358516 47488
rect 72884 47348 72948 47412
rect 107476 47348 107540 47412
rect 212540 47408 212604 47412
rect 212540 47352 212590 47408
rect 212590 47352 212604 47408
rect 212540 47348 212604 47352
rect 263876 47348 263940 47412
rect 306564 47408 306628 47412
rect 306564 47352 306614 47408
rect 306614 47352 306628 47408
rect 306564 47348 306628 47352
rect 109316 47212 109380 47276
rect 110420 47212 110484 47276
rect 248604 47212 248668 47276
rect 181812 46668 181876 46732
rect 162860 46532 162924 46596
rect 275836 46532 275900 46596
rect 74172 46184 74236 46188
rect 74172 46128 74222 46184
rect 74222 46128 74236 46184
rect 74172 46124 74236 46128
rect 118700 46184 118764 46188
rect 118700 46128 118714 46184
rect 118714 46128 118764 46184
rect 118700 46124 118764 46128
rect 158996 45988 159060 46052
rect 169668 46048 169732 46052
rect 169668 45992 169718 46048
rect 169718 45992 169732 46048
rect 169668 45988 169732 45992
rect 248972 45988 249036 46052
rect 262588 46048 262652 46052
rect 262588 45992 262602 46048
rect 262602 45992 262652 46048
rect 262588 45988 262652 45992
rect 336372 45988 336436 46052
rect 74540 45852 74604 45916
rect 157524 45852 157588 45916
rect 252836 45852 252900 45916
rect 147956 45716 148020 45780
rect 204260 45308 204324 45372
rect 113916 43268 113980 43332
rect 207756 37692 207820 37756
rect 301596 37752 301660 37756
rect 301596 37696 301610 37752
rect 301610 37696 301660 37752
rect 301596 37692 301660 37696
<< metal4 >>
rect 0 405398 4000 405520
rect 0 405162 122 405398
rect 358 405162 442 405398
rect 678 405162 762 405398
rect 998 405162 1082 405398
rect 1318 405162 1402 405398
rect 1638 405162 1722 405398
rect 1958 405162 2042 405398
rect 2278 405162 2362 405398
rect 2598 405162 2682 405398
rect 2918 405162 3002 405398
rect 3238 405162 3322 405398
rect 3558 405162 3642 405398
rect 3878 405162 4000 405398
rect 0 405078 4000 405162
rect 0 404842 122 405078
rect 358 404842 442 405078
rect 678 404842 762 405078
rect 998 404842 1082 405078
rect 1318 404842 1402 405078
rect 1638 404842 1722 405078
rect 1958 404842 2042 405078
rect 2278 404842 2362 405078
rect 2598 404842 2682 405078
rect 2918 404842 3002 405078
rect 3238 404842 3322 405078
rect 3558 404842 3642 405078
rect 3878 404842 4000 405078
rect 0 404758 4000 404842
rect 0 404522 122 404758
rect 358 404522 442 404758
rect 678 404522 762 404758
rect 998 404522 1082 404758
rect 1318 404522 1402 404758
rect 1638 404522 1722 404758
rect 1958 404522 2042 404758
rect 2278 404522 2362 404758
rect 2598 404522 2682 404758
rect 2918 404522 3002 404758
rect 3238 404522 3322 404758
rect 3558 404522 3642 404758
rect 3878 404522 4000 404758
rect 0 404438 4000 404522
rect 0 404202 122 404438
rect 358 404202 442 404438
rect 678 404202 762 404438
rect 998 404202 1082 404438
rect 1318 404202 1402 404438
rect 1638 404202 1722 404438
rect 1958 404202 2042 404438
rect 2278 404202 2362 404438
rect 2598 404202 2682 404438
rect 2918 404202 3002 404438
rect 3238 404202 3322 404438
rect 3558 404202 3642 404438
rect 3878 404202 4000 404438
rect 0 404118 4000 404202
rect 0 403882 122 404118
rect 358 403882 442 404118
rect 678 403882 762 404118
rect 998 403882 1082 404118
rect 1318 403882 1402 404118
rect 1638 403882 1722 404118
rect 1958 403882 2042 404118
rect 2278 403882 2362 404118
rect 2598 403882 2682 404118
rect 2918 403882 3002 404118
rect 3238 403882 3322 404118
rect 3558 403882 3642 404118
rect 3878 403882 4000 404118
rect 0 403798 4000 403882
rect 0 403562 122 403798
rect 358 403562 442 403798
rect 678 403562 762 403798
rect 998 403562 1082 403798
rect 1318 403562 1402 403798
rect 1638 403562 1722 403798
rect 1958 403562 2042 403798
rect 2278 403562 2362 403798
rect 2598 403562 2682 403798
rect 2918 403562 3002 403798
rect 3238 403562 3322 403798
rect 3558 403562 3642 403798
rect 3878 403562 4000 403798
rect 0 403478 4000 403562
rect 0 403242 122 403478
rect 358 403242 442 403478
rect 678 403242 762 403478
rect 998 403242 1082 403478
rect 1318 403242 1402 403478
rect 1638 403242 1722 403478
rect 1958 403242 2042 403478
rect 2278 403242 2362 403478
rect 2598 403242 2682 403478
rect 2918 403242 3002 403478
rect 3238 403242 3322 403478
rect 3558 403242 3642 403478
rect 3878 403242 4000 403478
rect 0 403158 4000 403242
rect 0 402922 122 403158
rect 358 402922 442 403158
rect 678 402922 762 403158
rect 998 402922 1082 403158
rect 1318 402922 1402 403158
rect 1638 402922 1722 403158
rect 1958 402922 2042 403158
rect 2278 402922 2362 403158
rect 2598 402922 2682 403158
rect 2918 402922 3002 403158
rect 3238 402922 3322 403158
rect 3558 402922 3642 403158
rect 3878 402922 4000 403158
rect 0 402838 4000 402922
rect 0 402602 122 402838
rect 358 402602 442 402838
rect 678 402602 762 402838
rect 998 402602 1082 402838
rect 1318 402602 1402 402838
rect 1638 402602 1722 402838
rect 1958 402602 2042 402838
rect 2278 402602 2362 402838
rect 2598 402602 2682 402838
rect 2918 402602 3002 402838
rect 3238 402602 3322 402838
rect 3558 402602 3642 402838
rect 3878 402602 4000 402838
rect 0 402518 4000 402602
rect 0 402282 122 402518
rect 358 402282 442 402518
rect 678 402282 762 402518
rect 998 402282 1082 402518
rect 1318 402282 1402 402518
rect 1638 402282 1722 402518
rect 1958 402282 2042 402518
rect 2278 402282 2362 402518
rect 2598 402282 2682 402518
rect 2918 402282 3002 402518
rect 3238 402282 3322 402518
rect 3558 402282 3642 402518
rect 3878 402282 4000 402518
rect 0 402198 4000 402282
rect 0 401962 122 402198
rect 358 401962 442 402198
rect 678 401962 762 402198
rect 998 401962 1082 402198
rect 1318 401962 1402 402198
rect 1638 401962 1722 402198
rect 1958 401962 2042 402198
rect 2278 401962 2362 402198
rect 2598 401962 2682 402198
rect 2918 401962 3002 402198
rect 3238 401962 3322 402198
rect 3558 401962 3642 402198
rect 3878 401962 4000 402198
rect 0 401878 4000 401962
rect 0 401642 122 401878
rect 358 401642 442 401878
rect 678 401642 762 401878
rect 998 401642 1082 401878
rect 1318 401642 1402 401878
rect 1638 401642 1722 401878
rect 1958 401642 2042 401878
rect 2278 401642 2362 401878
rect 2598 401642 2682 401878
rect 2918 401642 3002 401878
rect 3238 401642 3322 401878
rect 3558 401642 3642 401878
rect 3878 401642 4000 401878
rect 0 376432 4000 401642
rect 440740 405398 444740 405520
rect 440740 405162 440862 405398
rect 441098 405162 441182 405398
rect 441418 405162 441502 405398
rect 441738 405162 441822 405398
rect 442058 405162 442142 405398
rect 442378 405162 442462 405398
rect 442698 405162 442782 405398
rect 443018 405162 443102 405398
rect 443338 405162 443422 405398
rect 443658 405162 443742 405398
rect 443978 405162 444062 405398
rect 444298 405162 444382 405398
rect 444618 405162 444740 405398
rect 440740 405078 444740 405162
rect 440740 404842 440862 405078
rect 441098 404842 441182 405078
rect 441418 404842 441502 405078
rect 441738 404842 441822 405078
rect 442058 404842 442142 405078
rect 442378 404842 442462 405078
rect 442698 404842 442782 405078
rect 443018 404842 443102 405078
rect 443338 404842 443422 405078
rect 443658 404842 443742 405078
rect 443978 404842 444062 405078
rect 444298 404842 444382 405078
rect 444618 404842 444740 405078
rect 440740 404758 444740 404842
rect 440740 404522 440862 404758
rect 441098 404522 441182 404758
rect 441418 404522 441502 404758
rect 441738 404522 441822 404758
rect 442058 404522 442142 404758
rect 442378 404522 442462 404758
rect 442698 404522 442782 404758
rect 443018 404522 443102 404758
rect 443338 404522 443422 404758
rect 443658 404522 443742 404758
rect 443978 404522 444062 404758
rect 444298 404522 444382 404758
rect 444618 404522 444740 404758
rect 440740 404438 444740 404522
rect 440740 404202 440862 404438
rect 441098 404202 441182 404438
rect 441418 404202 441502 404438
rect 441738 404202 441822 404438
rect 442058 404202 442142 404438
rect 442378 404202 442462 404438
rect 442698 404202 442782 404438
rect 443018 404202 443102 404438
rect 443338 404202 443422 404438
rect 443658 404202 443742 404438
rect 443978 404202 444062 404438
rect 444298 404202 444382 404438
rect 444618 404202 444740 404438
rect 440740 404118 444740 404202
rect 440740 403882 440862 404118
rect 441098 403882 441182 404118
rect 441418 403882 441502 404118
rect 441738 403882 441822 404118
rect 442058 403882 442142 404118
rect 442378 403882 442462 404118
rect 442698 403882 442782 404118
rect 443018 403882 443102 404118
rect 443338 403882 443422 404118
rect 443658 403882 443742 404118
rect 443978 403882 444062 404118
rect 444298 403882 444382 404118
rect 444618 403882 444740 404118
rect 440740 403798 444740 403882
rect 440740 403562 440862 403798
rect 441098 403562 441182 403798
rect 441418 403562 441502 403798
rect 441738 403562 441822 403798
rect 442058 403562 442142 403798
rect 442378 403562 442462 403798
rect 442698 403562 442782 403798
rect 443018 403562 443102 403798
rect 443338 403562 443422 403798
rect 443658 403562 443742 403798
rect 443978 403562 444062 403798
rect 444298 403562 444382 403798
rect 444618 403562 444740 403798
rect 440740 403478 444740 403562
rect 440740 403242 440862 403478
rect 441098 403242 441182 403478
rect 441418 403242 441502 403478
rect 441738 403242 441822 403478
rect 442058 403242 442142 403478
rect 442378 403242 442462 403478
rect 442698 403242 442782 403478
rect 443018 403242 443102 403478
rect 443338 403242 443422 403478
rect 443658 403242 443742 403478
rect 443978 403242 444062 403478
rect 444298 403242 444382 403478
rect 444618 403242 444740 403478
rect 440740 403158 444740 403242
rect 440740 402922 440862 403158
rect 441098 402922 441182 403158
rect 441418 402922 441502 403158
rect 441738 402922 441822 403158
rect 442058 402922 442142 403158
rect 442378 402922 442462 403158
rect 442698 402922 442782 403158
rect 443018 402922 443102 403158
rect 443338 402922 443422 403158
rect 443658 402922 443742 403158
rect 443978 402922 444062 403158
rect 444298 402922 444382 403158
rect 444618 402922 444740 403158
rect 440740 402838 444740 402922
rect 440740 402602 440862 402838
rect 441098 402602 441182 402838
rect 441418 402602 441502 402838
rect 441738 402602 441822 402838
rect 442058 402602 442142 402838
rect 442378 402602 442462 402838
rect 442698 402602 442782 402838
rect 443018 402602 443102 402838
rect 443338 402602 443422 402838
rect 443658 402602 443742 402838
rect 443978 402602 444062 402838
rect 444298 402602 444382 402838
rect 444618 402602 444740 402838
rect 440740 402518 444740 402602
rect 440740 402282 440862 402518
rect 441098 402282 441182 402518
rect 441418 402282 441502 402518
rect 441738 402282 441822 402518
rect 442058 402282 442142 402518
rect 442378 402282 442462 402518
rect 442698 402282 442782 402518
rect 443018 402282 443102 402518
rect 443338 402282 443422 402518
rect 443658 402282 443742 402518
rect 443978 402282 444062 402518
rect 444298 402282 444382 402518
rect 444618 402282 444740 402518
rect 440740 402198 444740 402282
rect 440740 401962 440862 402198
rect 441098 401962 441182 402198
rect 441418 401962 441502 402198
rect 441738 401962 441822 402198
rect 442058 401962 442142 402198
rect 442378 401962 442462 402198
rect 442698 401962 442782 402198
rect 443018 401962 443102 402198
rect 443338 401962 443422 402198
rect 443658 401962 443742 402198
rect 443978 401962 444062 402198
rect 444298 401962 444382 402198
rect 444618 401962 444740 402198
rect 440740 401878 444740 401962
rect 440740 401642 440862 401878
rect 441098 401642 441182 401878
rect 441418 401642 441502 401878
rect 441738 401642 441822 401878
rect 442058 401642 442142 401878
rect 442378 401642 442462 401878
rect 442698 401642 442782 401878
rect 443018 401642 443102 401878
rect 443338 401642 443422 401878
rect 443658 401642 443742 401878
rect 443978 401642 444062 401878
rect 444298 401642 444382 401878
rect 444618 401642 444740 401878
rect 0 376196 122 376432
rect 358 376196 442 376432
rect 678 376196 762 376432
rect 998 376196 1082 376432
rect 1318 376196 1402 376432
rect 1638 376196 1722 376432
rect 1958 376196 2042 376432
rect 2278 376196 2362 376432
rect 2598 376196 2682 376432
rect 2918 376196 3002 376432
rect 3238 376196 3322 376432
rect 3558 376196 3642 376432
rect 3878 376196 4000 376432
rect 0 345796 4000 376196
rect 0 345560 122 345796
rect 358 345560 442 345796
rect 678 345560 762 345796
rect 998 345560 1082 345796
rect 1318 345560 1402 345796
rect 1638 345560 1722 345796
rect 1958 345560 2042 345796
rect 2278 345560 2362 345796
rect 2598 345560 2682 345796
rect 2918 345560 3002 345796
rect 3238 345560 3322 345796
rect 3558 345560 3642 345796
rect 3878 345560 4000 345796
rect 0 315160 4000 345560
rect 0 314924 122 315160
rect 358 314924 442 315160
rect 678 314924 762 315160
rect 998 314924 1082 315160
rect 1318 314924 1402 315160
rect 1638 314924 1722 315160
rect 1958 314924 2042 315160
rect 2278 314924 2362 315160
rect 2598 314924 2682 315160
rect 2918 314924 3002 315160
rect 3238 314924 3322 315160
rect 3558 314924 3642 315160
rect 3878 314924 4000 315160
rect 0 284524 4000 314924
rect 0 284288 122 284524
rect 358 284288 442 284524
rect 678 284288 762 284524
rect 998 284288 1082 284524
rect 1318 284288 1402 284524
rect 1638 284288 1722 284524
rect 1958 284288 2042 284524
rect 2278 284288 2362 284524
rect 2598 284288 2682 284524
rect 2918 284288 3002 284524
rect 3238 284288 3322 284524
rect 3558 284288 3642 284524
rect 3878 284288 4000 284524
rect 0 253888 4000 284288
rect 0 253652 122 253888
rect 358 253652 442 253888
rect 678 253652 762 253888
rect 998 253652 1082 253888
rect 1318 253652 1402 253888
rect 1638 253652 1722 253888
rect 1958 253652 2042 253888
rect 2278 253652 2362 253888
rect 2598 253652 2682 253888
rect 2918 253652 3002 253888
rect 3238 253652 3322 253888
rect 3558 253652 3642 253888
rect 3878 253652 4000 253888
rect 0 223252 4000 253652
rect 0 223016 122 223252
rect 358 223016 442 223252
rect 678 223016 762 223252
rect 998 223016 1082 223252
rect 1318 223016 1402 223252
rect 1638 223016 1722 223252
rect 1958 223016 2042 223252
rect 2278 223016 2362 223252
rect 2598 223016 2682 223252
rect 2918 223016 3002 223252
rect 3238 223016 3322 223252
rect 3558 223016 3642 223252
rect 3878 223016 4000 223252
rect 0 192616 4000 223016
rect 0 192380 122 192616
rect 358 192380 442 192616
rect 678 192380 762 192616
rect 998 192380 1082 192616
rect 1318 192380 1402 192616
rect 1638 192380 1722 192616
rect 1958 192380 2042 192616
rect 2278 192380 2362 192616
rect 2598 192380 2682 192616
rect 2918 192380 3002 192616
rect 3238 192380 3322 192616
rect 3558 192380 3642 192616
rect 3878 192380 4000 192616
rect 0 161980 4000 192380
rect 0 161744 122 161980
rect 358 161744 442 161980
rect 678 161744 762 161980
rect 998 161744 1082 161980
rect 1318 161744 1402 161980
rect 1638 161744 1722 161980
rect 1958 161744 2042 161980
rect 2278 161744 2362 161980
rect 2598 161744 2682 161980
rect 2918 161744 3002 161980
rect 3238 161744 3322 161980
rect 3558 161744 3642 161980
rect 3878 161744 4000 161980
rect 0 131344 4000 161744
rect 0 131108 122 131344
rect 358 131108 442 131344
rect 678 131108 762 131344
rect 998 131108 1082 131344
rect 1318 131108 1402 131344
rect 1638 131108 1722 131344
rect 1958 131108 2042 131344
rect 2278 131108 2362 131344
rect 2598 131108 2682 131344
rect 2918 131108 3002 131344
rect 3238 131108 3322 131344
rect 3558 131108 3642 131344
rect 3878 131108 4000 131344
rect 0 100708 4000 131108
rect 0 100472 122 100708
rect 358 100472 442 100708
rect 678 100472 762 100708
rect 998 100472 1082 100708
rect 1318 100472 1402 100708
rect 1638 100472 1722 100708
rect 1958 100472 2042 100708
rect 2278 100472 2362 100708
rect 2598 100472 2682 100708
rect 2918 100472 3002 100708
rect 3238 100472 3322 100708
rect 3558 100472 3642 100708
rect 3878 100472 4000 100708
rect 0 70072 4000 100472
rect 0 69836 122 70072
rect 358 69836 442 70072
rect 678 69836 762 70072
rect 998 69836 1082 70072
rect 1318 69836 1402 70072
rect 1638 69836 1722 70072
rect 1958 69836 2042 70072
rect 2278 69836 2362 70072
rect 2598 69836 2682 70072
rect 2918 69836 3002 70072
rect 3238 69836 3322 70072
rect 3558 69836 3642 70072
rect 3878 69836 4000 70072
rect 0 39436 4000 69836
rect 0 39200 122 39436
rect 358 39200 442 39436
rect 678 39200 762 39436
rect 998 39200 1082 39436
rect 1318 39200 1402 39436
rect 1638 39200 1722 39436
rect 1958 39200 2042 39436
rect 2278 39200 2362 39436
rect 2598 39200 2682 39436
rect 2918 39200 3002 39436
rect 3238 39200 3322 39436
rect 3558 39200 3642 39436
rect 3878 39200 4000 39436
rect 0 3878 4000 39200
rect 5000 400398 9000 400520
rect 5000 400162 5122 400398
rect 5358 400162 5442 400398
rect 5678 400162 5762 400398
rect 5998 400162 6082 400398
rect 6318 400162 6402 400398
rect 6638 400162 6722 400398
rect 6958 400162 7042 400398
rect 7278 400162 7362 400398
rect 7598 400162 7682 400398
rect 7918 400162 8002 400398
rect 8238 400162 8322 400398
rect 8558 400162 8642 400398
rect 8878 400162 9000 400398
rect 5000 400078 9000 400162
rect 5000 399842 5122 400078
rect 5358 399842 5442 400078
rect 5678 399842 5762 400078
rect 5998 399842 6082 400078
rect 6318 399842 6402 400078
rect 6638 399842 6722 400078
rect 6958 399842 7042 400078
rect 7278 399842 7362 400078
rect 7598 399842 7682 400078
rect 7918 399842 8002 400078
rect 8238 399842 8322 400078
rect 8558 399842 8642 400078
rect 8878 399842 9000 400078
rect 5000 399758 9000 399842
rect 5000 399522 5122 399758
rect 5358 399522 5442 399758
rect 5678 399522 5762 399758
rect 5998 399522 6082 399758
rect 6318 399522 6402 399758
rect 6638 399522 6722 399758
rect 6958 399522 7042 399758
rect 7278 399522 7362 399758
rect 7598 399522 7682 399758
rect 7918 399522 8002 399758
rect 8238 399522 8322 399758
rect 8558 399522 8642 399758
rect 8878 399522 9000 399758
rect 5000 399438 9000 399522
rect 5000 399202 5122 399438
rect 5358 399202 5442 399438
rect 5678 399202 5762 399438
rect 5998 399202 6082 399438
rect 6318 399202 6402 399438
rect 6638 399202 6722 399438
rect 6958 399202 7042 399438
rect 7278 399202 7362 399438
rect 7598 399202 7682 399438
rect 7918 399202 8002 399438
rect 8238 399202 8322 399438
rect 8558 399202 8642 399438
rect 8878 399202 9000 399438
rect 5000 399118 9000 399202
rect 5000 398882 5122 399118
rect 5358 398882 5442 399118
rect 5678 398882 5762 399118
rect 5998 398882 6082 399118
rect 6318 398882 6402 399118
rect 6638 398882 6722 399118
rect 6958 398882 7042 399118
rect 7278 398882 7362 399118
rect 7598 398882 7682 399118
rect 7918 398882 8002 399118
rect 8238 398882 8322 399118
rect 8558 398882 8642 399118
rect 8878 398882 9000 399118
rect 5000 398798 9000 398882
rect 5000 398562 5122 398798
rect 5358 398562 5442 398798
rect 5678 398562 5762 398798
rect 5998 398562 6082 398798
rect 6318 398562 6402 398798
rect 6638 398562 6722 398798
rect 6958 398562 7042 398798
rect 7278 398562 7362 398798
rect 7598 398562 7682 398798
rect 7918 398562 8002 398798
rect 8238 398562 8322 398798
rect 8558 398562 8642 398798
rect 8878 398562 9000 398798
rect 5000 398478 9000 398562
rect 5000 398242 5122 398478
rect 5358 398242 5442 398478
rect 5678 398242 5762 398478
rect 5998 398242 6082 398478
rect 6318 398242 6402 398478
rect 6638 398242 6722 398478
rect 6958 398242 7042 398478
rect 7278 398242 7362 398478
rect 7598 398242 7682 398478
rect 7918 398242 8002 398478
rect 8238 398242 8322 398478
rect 8558 398242 8642 398478
rect 8878 398242 9000 398478
rect 5000 398158 9000 398242
rect 5000 397922 5122 398158
rect 5358 397922 5442 398158
rect 5678 397922 5762 398158
rect 5998 397922 6082 398158
rect 6318 397922 6402 398158
rect 6638 397922 6722 398158
rect 6958 397922 7042 398158
rect 7278 397922 7362 398158
rect 7598 397922 7682 398158
rect 7918 397922 8002 398158
rect 8238 397922 8322 398158
rect 8558 397922 8642 398158
rect 8878 397922 9000 398158
rect 5000 397838 9000 397922
rect 5000 397602 5122 397838
rect 5358 397602 5442 397838
rect 5678 397602 5762 397838
rect 5998 397602 6082 397838
rect 6318 397602 6402 397838
rect 6638 397602 6722 397838
rect 6958 397602 7042 397838
rect 7278 397602 7362 397838
rect 7598 397602 7682 397838
rect 7918 397602 8002 397838
rect 8238 397602 8322 397838
rect 8558 397602 8642 397838
rect 8878 397602 9000 397838
rect 5000 397518 9000 397602
rect 5000 397282 5122 397518
rect 5358 397282 5442 397518
rect 5678 397282 5762 397518
rect 5998 397282 6082 397518
rect 6318 397282 6402 397518
rect 6638 397282 6722 397518
rect 6958 397282 7042 397518
rect 7278 397282 7362 397518
rect 7598 397282 7682 397518
rect 7918 397282 8002 397518
rect 8238 397282 8322 397518
rect 8558 397282 8642 397518
rect 8878 397282 9000 397518
rect 5000 397198 9000 397282
rect 5000 396962 5122 397198
rect 5358 396962 5442 397198
rect 5678 396962 5762 397198
rect 5998 396962 6082 397198
rect 6318 396962 6402 397198
rect 6638 396962 6722 397198
rect 6958 396962 7042 397198
rect 7278 396962 7362 397198
rect 7598 396962 7682 397198
rect 7918 396962 8002 397198
rect 8238 396962 8322 397198
rect 8558 396962 8642 397198
rect 8878 396962 9000 397198
rect 5000 396878 9000 396962
rect 5000 396642 5122 396878
rect 5358 396642 5442 396878
rect 5678 396642 5762 396878
rect 5998 396642 6082 396878
rect 6318 396642 6402 396878
rect 6638 396642 6722 396878
rect 6958 396642 7042 396878
rect 7278 396642 7362 396878
rect 7598 396642 7682 396878
rect 7918 396642 8002 396878
rect 8238 396642 8322 396878
rect 8558 396642 8642 396878
rect 8878 396642 9000 396878
rect 5000 391750 9000 396642
rect 435740 400398 439740 400520
rect 435740 400162 435862 400398
rect 436098 400162 436182 400398
rect 436418 400162 436502 400398
rect 436738 400162 436822 400398
rect 437058 400162 437142 400398
rect 437378 400162 437462 400398
rect 437698 400162 437782 400398
rect 438018 400162 438102 400398
rect 438338 400162 438422 400398
rect 438658 400162 438742 400398
rect 438978 400162 439062 400398
rect 439298 400162 439382 400398
rect 439618 400162 439740 400398
rect 435740 400078 439740 400162
rect 435740 399842 435862 400078
rect 436098 399842 436182 400078
rect 436418 399842 436502 400078
rect 436738 399842 436822 400078
rect 437058 399842 437142 400078
rect 437378 399842 437462 400078
rect 437698 399842 437782 400078
rect 438018 399842 438102 400078
rect 438338 399842 438422 400078
rect 438658 399842 438742 400078
rect 438978 399842 439062 400078
rect 439298 399842 439382 400078
rect 439618 399842 439740 400078
rect 435740 399758 439740 399842
rect 435740 399522 435862 399758
rect 436098 399522 436182 399758
rect 436418 399522 436502 399758
rect 436738 399522 436822 399758
rect 437058 399522 437142 399758
rect 437378 399522 437462 399758
rect 437698 399522 437782 399758
rect 438018 399522 438102 399758
rect 438338 399522 438422 399758
rect 438658 399522 438742 399758
rect 438978 399522 439062 399758
rect 439298 399522 439382 399758
rect 439618 399522 439740 399758
rect 435740 399438 439740 399522
rect 435740 399202 435862 399438
rect 436098 399202 436182 399438
rect 436418 399202 436502 399438
rect 436738 399202 436822 399438
rect 437058 399202 437142 399438
rect 437378 399202 437462 399438
rect 437698 399202 437782 399438
rect 438018 399202 438102 399438
rect 438338 399202 438422 399438
rect 438658 399202 438742 399438
rect 438978 399202 439062 399438
rect 439298 399202 439382 399438
rect 439618 399202 439740 399438
rect 435740 399118 439740 399202
rect 435740 398882 435862 399118
rect 436098 398882 436182 399118
rect 436418 398882 436502 399118
rect 436738 398882 436822 399118
rect 437058 398882 437142 399118
rect 437378 398882 437462 399118
rect 437698 398882 437782 399118
rect 438018 398882 438102 399118
rect 438338 398882 438422 399118
rect 438658 398882 438742 399118
rect 438978 398882 439062 399118
rect 439298 398882 439382 399118
rect 439618 398882 439740 399118
rect 435740 398798 439740 398882
rect 435740 398562 435862 398798
rect 436098 398562 436182 398798
rect 436418 398562 436502 398798
rect 436738 398562 436822 398798
rect 437058 398562 437142 398798
rect 437378 398562 437462 398798
rect 437698 398562 437782 398798
rect 438018 398562 438102 398798
rect 438338 398562 438422 398798
rect 438658 398562 438742 398798
rect 438978 398562 439062 398798
rect 439298 398562 439382 398798
rect 439618 398562 439740 398798
rect 435740 398478 439740 398562
rect 435740 398242 435862 398478
rect 436098 398242 436182 398478
rect 436418 398242 436502 398478
rect 436738 398242 436822 398478
rect 437058 398242 437142 398478
rect 437378 398242 437462 398478
rect 437698 398242 437782 398478
rect 438018 398242 438102 398478
rect 438338 398242 438422 398478
rect 438658 398242 438742 398478
rect 438978 398242 439062 398478
rect 439298 398242 439382 398478
rect 439618 398242 439740 398478
rect 435740 398158 439740 398242
rect 435740 397922 435862 398158
rect 436098 397922 436182 398158
rect 436418 397922 436502 398158
rect 436738 397922 436822 398158
rect 437058 397922 437142 398158
rect 437378 397922 437462 398158
rect 437698 397922 437782 398158
rect 438018 397922 438102 398158
rect 438338 397922 438422 398158
rect 438658 397922 438742 398158
rect 438978 397922 439062 398158
rect 439298 397922 439382 398158
rect 439618 397922 439740 398158
rect 435740 397838 439740 397922
rect 435740 397602 435862 397838
rect 436098 397602 436182 397838
rect 436418 397602 436502 397838
rect 436738 397602 436822 397838
rect 437058 397602 437142 397838
rect 437378 397602 437462 397838
rect 437698 397602 437782 397838
rect 438018 397602 438102 397838
rect 438338 397602 438422 397838
rect 438658 397602 438742 397838
rect 438978 397602 439062 397838
rect 439298 397602 439382 397838
rect 439618 397602 439740 397838
rect 435740 397518 439740 397602
rect 435740 397282 435862 397518
rect 436098 397282 436182 397518
rect 436418 397282 436502 397518
rect 436738 397282 436822 397518
rect 437058 397282 437142 397518
rect 437378 397282 437462 397518
rect 437698 397282 437782 397518
rect 438018 397282 438102 397518
rect 438338 397282 438422 397518
rect 438658 397282 438742 397518
rect 438978 397282 439062 397518
rect 439298 397282 439382 397518
rect 439618 397282 439740 397518
rect 435740 397198 439740 397282
rect 435740 396962 435862 397198
rect 436098 396962 436182 397198
rect 436418 396962 436502 397198
rect 436738 396962 436822 397198
rect 437058 396962 437142 397198
rect 437378 396962 437462 397198
rect 437698 396962 437782 397198
rect 438018 396962 438102 397198
rect 438338 396962 438422 397198
rect 438658 396962 438742 397198
rect 438978 396962 439062 397198
rect 439298 396962 439382 397198
rect 439618 396962 439740 397198
rect 435740 396878 439740 396962
rect 435740 396642 435862 396878
rect 436098 396642 436182 396878
rect 436418 396642 436502 396878
rect 436738 396642 436822 396878
rect 437058 396642 437142 396878
rect 437378 396642 437462 396878
rect 437698 396642 437782 396878
rect 438018 396642 438102 396878
rect 438338 396642 438422 396878
rect 438658 396642 438742 396878
rect 438978 396642 439062 396878
rect 439298 396642 439382 396878
rect 439618 396642 439740 396878
rect 280251 393804 280317 393805
rect 280251 393740 280252 393804
rect 280316 393740 280317 393804
rect 280251 393739 280317 393740
rect 323123 393804 323189 393805
rect 323123 393740 323124 393804
rect 323188 393740 323189 393804
rect 323123 393739 323189 393740
rect 5000 391514 5122 391750
rect 5358 391514 5442 391750
rect 5678 391514 5762 391750
rect 5998 391514 6082 391750
rect 6318 391514 6402 391750
rect 6638 391514 6722 391750
rect 6958 391514 7042 391750
rect 7278 391514 7362 391750
rect 7598 391514 7682 391750
rect 7918 391514 8002 391750
rect 8238 391514 8322 391750
rect 8558 391514 8642 391750
rect 8878 391514 9000 391750
rect 5000 361114 9000 391514
rect 97355 367284 97421 367285
rect 97355 367220 97356 367284
rect 97420 367220 97421 367284
rect 97355 367219 97421 367220
rect 5000 360878 5122 361114
rect 5358 360878 5442 361114
rect 5678 360878 5762 361114
rect 5998 360878 6082 361114
rect 6318 360878 6402 361114
rect 6638 360878 6722 361114
rect 6958 360878 7042 361114
rect 7278 360878 7362 361114
rect 7598 360878 7682 361114
rect 7918 360878 8002 361114
rect 8238 360878 8322 361114
rect 8558 360878 8642 361114
rect 8878 360878 9000 361114
rect 5000 330478 9000 360878
rect 97358 352053 97418 367219
rect 97355 352052 97421 352053
rect 97355 351988 97356 352052
rect 97420 351988 97421 352052
rect 97355 351987 97421 351988
rect 104899 333828 104965 333829
rect 104899 333764 104900 333828
rect 104964 333764 104965 333828
rect 104899 333763 104965 333764
rect 5000 330242 5122 330478
rect 5358 330242 5442 330478
rect 5678 330242 5762 330478
rect 5998 330242 6082 330478
rect 6318 330242 6402 330478
rect 6638 330242 6722 330478
rect 6958 330242 7042 330478
rect 7278 330242 7362 330478
rect 7598 330242 7682 330478
rect 7918 330242 8002 330478
rect 8238 330242 8322 330478
rect 8558 330242 8642 330478
rect 8878 330242 9000 330478
rect 5000 299842 9000 330242
rect 52643 327436 52709 327437
rect 52643 327372 52644 327436
rect 52708 327372 52709 327436
rect 52643 327371 52709 327372
rect 54667 327436 54733 327437
rect 54667 327372 54668 327436
rect 54732 327372 54733 327436
rect 54667 327371 54733 327372
rect 55403 327436 55469 327437
rect 55403 327372 55404 327436
rect 55468 327372 55469 327436
rect 55403 327371 55469 327372
rect 52646 300645 52706 327371
rect 54670 306221 54730 327371
rect 55219 317916 55285 317917
rect 55219 317852 55220 317916
rect 55284 317852 55285 317916
rect 55219 317851 55285 317852
rect 55035 310436 55101 310437
rect 55035 310372 55036 310436
rect 55100 310434 55101 310436
rect 55222 310434 55282 317851
rect 55406 315877 55466 327371
rect 104902 320042 104962 333763
rect 212171 333556 212237 333557
rect 212171 333492 212172 333556
rect 212236 333492 212237 333556
rect 212171 333491 212237 333492
rect 159550 330157 159610 331366
rect 159547 330156 159613 330157
rect 159547 330092 159548 330156
rect 159612 330092 159613 330156
rect 159547 330091 159613 330092
rect 168566 327437 168626 332046
rect 204443 331652 204509 331653
rect 204443 331602 204444 331652
rect 204508 331602 204509 331652
rect 212174 329562 212234 333491
rect 251550 330021 251610 331366
rect 252286 330157 252346 331366
rect 252283 330156 252349 330157
rect 252283 330092 252284 330156
rect 252348 330092 252349 330156
rect 252283 330091 252349 330092
rect 253022 330021 253082 331366
rect 251547 330020 251613 330021
rect 251547 329956 251548 330020
rect 251612 329956 251613 330020
rect 251547 329955 251613 329956
rect 253019 330020 253085 330021
rect 253019 329956 253020 330020
rect 253084 329956 253085 330020
rect 253019 329955 253085 329956
rect 262406 327573 262466 333406
rect 280254 333149 280314 393739
rect 285035 367284 285101 367285
rect 285035 367220 285036 367284
rect 285100 367220 285101 367284
rect 285035 367219 285101 367220
rect 285038 351645 285098 367219
rect 285035 351644 285101 351645
rect 285035 351580 285036 351644
rect 285100 351580 285101 351644
rect 285035 351579 285101 351580
rect 280251 333148 280317 333149
rect 280251 333084 280252 333148
rect 280316 333084 280317 333148
rect 280251 333083 280317 333084
rect 294051 331652 294117 331653
rect 294051 331602 294052 331652
rect 294116 331602 294117 331652
rect 262403 327572 262469 327573
rect 262403 327508 262404 327572
rect 262468 327508 262469 327572
rect 262403 327507 262469 327508
rect 168563 327436 168629 327437
rect 168563 327372 168564 327436
rect 168628 327372 168629 327436
rect 168563 327371 168629 327372
rect 153291 326348 153357 326349
rect 153291 326284 153292 326348
rect 153356 326284 153357 326348
rect 153291 326283 153357 326284
rect 55403 315876 55469 315877
rect 55403 315812 55404 315876
rect 55468 315812 55469 315876
rect 55403 315811 55469 315812
rect 55100 310374 55282 310434
rect 55100 310372 55101 310374
rect 55035 310371 55101 310372
rect 54667 306220 54733 306221
rect 54667 306156 54668 306220
rect 54732 306156 54733 306220
rect 54667 306155 54733 306156
rect 52643 300644 52709 300645
rect 52643 300580 52644 300644
rect 52708 300580 52709 300644
rect 52643 300579 52709 300580
rect 5000 299606 5122 299842
rect 5358 299606 5442 299842
rect 5678 299606 5762 299842
rect 5998 299606 6082 299842
rect 6318 299606 6402 299842
rect 6638 299606 6722 299842
rect 6958 299606 7042 299842
rect 7278 299606 7362 299842
rect 7598 299606 7682 299842
rect 7918 299606 8002 299842
rect 8238 299606 8322 299842
rect 8558 299606 8642 299842
rect 8878 299606 9000 299842
rect 5000 269206 9000 299606
rect 5000 268970 5122 269206
rect 5358 268970 5442 269206
rect 5678 268970 5762 269206
rect 5998 268970 6082 269206
rect 6318 268970 6402 269206
rect 6638 268970 6722 269206
rect 6958 268970 7042 269206
rect 7278 268970 7362 269206
rect 7598 268970 7682 269206
rect 7918 268970 8002 269206
rect 8238 268970 8322 269206
rect 8558 268970 8642 269206
rect 8878 268970 9000 269206
rect 5000 238570 9000 268970
rect 52646 265557 52706 300579
rect 54670 265557 54730 306155
rect 55222 266645 55282 310374
rect 55219 266644 55285 266645
rect 55219 266580 55220 266644
rect 55284 266580 55285 266644
rect 55219 266579 55285 266580
rect 55406 265557 55466 315811
rect 153294 315877 153354 326283
rect 153291 315876 153357 315877
rect 153291 315812 153292 315876
rect 153356 315812 153357 315876
rect 153291 315811 153357 315812
rect 104718 315202 104778 315726
rect 104464 315160 104784 315202
rect 104464 314924 104506 315160
rect 104742 314924 104784 315160
rect 104464 314882 104784 314924
rect 198464 315160 198784 315202
rect 198464 314924 198506 315160
rect 198742 314924 198784 315160
rect 198464 314882 198784 314924
rect 292464 315160 292784 315202
rect 292464 314924 292506 315160
rect 292742 314924 292784 315160
rect 292464 314882 292784 314924
rect 104718 314602 104778 314882
rect 74539 305676 74605 305677
rect 74539 305612 74540 305676
rect 74604 305612 74605 305676
rect 74539 305611 74605 305612
rect 73987 304044 74053 304045
rect 73987 303980 73988 304044
rect 74052 303980 74053 304044
rect 73987 303979 74053 303980
rect 73803 300100 73869 300101
rect 73803 300036 73804 300100
rect 73868 300036 73869 300100
rect 73803 300035 73869 300036
rect 73435 291804 73501 291805
rect 73435 291740 73436 291804
rect 73500 291740 73501 291804
rect 73435 291739 73501 291740
rect 73438 286365 73498 291739
rect 73435 286364 73501 286365
rect 73435 286300 73436 286364
rect 73500 286300 73501 286364
rect 73435 286299 73501 286300
rect 73619 282828 73685 282829
rect 73619 282764 73620 282828
rect 73684 282764 73685 282828
rect 73619 282763 73685 282764
rect 73435 282012 73501 282013
rect 73435 281948 73436 282012
rect 73500 281948 73501 282012
rect 73435 281947 73501 281948
rect 73438 277389 73498 281947
rect 73435 277388 73501 277389
rect 73435 277324 73436 277388
rect 73500 277324 73501 277388
rect 73435 277323 73501 277324
rect 73435 277252 73501 277253
rect 73435 277188 73436 277252
rect 73500 277188 73501 277252
rect 73435 277187 73501 277188
rect 73438 270317 73498 277187
rect 73435 270316 73501 270317
rect 73435 270252 73436 270316
rect 73500 270252 73501 270316
rect 73435 270251 73501 270252
rect 73435 270180 73501 270181
rect 73435 270116 73436 270180
rect 73500 270116 73501 270180
rect 73435 270115 73501 270116
rect 52643 265556 52709 265557
rect 52643 265492 52644 265556
rect 52708 265492 52709 265556
rect 52643 265491 52709 265492
rect 54667 265556 54733 265557
rect 54667 265492 54668 265556
rect 54732 265492 54733 265556
rect 54667 265491 54733 265492
rect 55403 265556 55469 265557
rect 55403 265492 55404 265556
rect 55468 265492 55469 265556
rect 55403 265491 55469 265492
rect 73438 263381 73498 270115
rect 73435 263380 73501 263381
rect 73435 263316 73436 263380
rect 73500 263316 73501 263380
rect 73435 263315 73501 263316
rect 48963 255836 48964 255886
rect 49028 255836 49029 255886
rect 48963 255835 49029 255836
rect 49147 246108 49213 246109
rect 49147 246044 49148 246108
rect 49212 246044 49213 246108
rect 49147 246043 49213 246044
rect 46939 243524 47005 243525
rect 46939 243460 46940 243524
rect 47004 243460 47005 243524
rect 46939 243459 47005 243460
rect 46942 242522 47002 243459
rect 49150 241162 49210 246043
rect 49147 239852 49213 239853
rect 49147 239802 49148 239852
rect 49212 239802 49213 239852
rect 5000 238334 5122 238570
rect 5358 238334 5442 238570
rect 5678 238334 5762 238570
rect 5998 238334 6082 238570
rect 6318 238334 6402 238570
rect 6638 238334 6722 238570
rect 6958 238334 7042 238570
rect 7278 238334 7362 238570
rect 7598 238334 7682 238570
rect 7918 238334 8002 238570
rect 8238 238334 8322 238570
rect 8558 238334 8642 238570
rect 8878 238334 9000 238570
rect 5000 207934 9000 238334
rect 73435 236316 73501 236317
rect 73435 236252 73436 236316
rect 73500 236252 73501 236316
rect 73435 236251 73501 236252
rect 52643 232508 52709 232509
rect 52643 232444 52644 232508
rect 52708 232444 52709 232508
rect 52643 232443 52709 232444
rect 54667 232508 54733 232509
rect 54667 232444 54668 232508
rect 54732 232444 54733 232508
rect 54667 232443 54733 232444
rect 55587 232508 55653 232509
rect 55587 232444 55588 232508
rect 55652 232444 55653 232508
rect 55587 232443 55653 232444
rect 5000 207698 5122 207934
rect 5358 207698 5442 207934
rect 5678 207698 5762 207934
rect 5998 207698 6082 207934
rect 6318 207698 6402 207934
rect 6638 207698 6722 207934
rect 6958 207698 7042 207934
rect 7278 207698 7362 207934
rect 7598 207698 7682 207934
rect 7918 207698 8002 207934
rect 8238 207698 8322 207934
rect 8558 207698 8642 207934
rect 8878 207698 9000 207934
rect 5000 177298 9000 207698
rect 52646 206805 52706 232443
rect 54670 211021 54730 232443
rect 55403 226932 55469 226933
rect 55403 226868 55404 226932
rect 55468 226868 55469 226932
rect 55403 226867 55469 226868
rect 55406 222037 55466 226867
rect 55403 222036 55469 222037
rect 55403 221972 55404 222036
rect 55468 221972 55469 222036
rect 55403 221971 55469 221972
rect 55406 217954 55466 221971
rect 55590 221357 55650 232443
rect 55587 221356 55653 221357
rect 55587 221292 55588 221356
rect 55652 221292 55653 221356
rect 55587 221291 55653 221292
rect 56323 221356 56389 221357
rect 56323 221292 56324 221356
rect 56388 221292 56389 221356
rect 56323 221291 56389 221292
rect 55406 217894 55834 217954
rect 55774 215234 55834 217894
rect 55406 215174 55834 215234
rect 54667 211020 54733 211021
rect 54667 210956 54668 211020
rect 54732 210956 54733 211020
rect 54667 210955 54733 210956
rect 52643 206804 52709 206805
rect 52643 206740 52644 206804
rect 52708 206740 52709 206804
rect 52643 206739 52709 206740
rect 5000 177062 5122 177298
rect 5358 177062 5442 177298
rect 5678 177062 5762 177298
rect 5998 177062 6082 177298
rect 6318 177062 6402 177298
rect 6638 177062 6722 177298
rect 6958 177062 7042 177298
rect 7278 177062 7362 177298
rect 7598 177062 7682 177298
rect 7918 177062 8002 177298
rect 8238 177062 8322 177298
rect 8558 177062 8642 177298
rect 8878 177062 9000 177298
rect 5000 146662 9000 177062
rect 52646 172941 52706 206739
rect 54670 172941 54730 210955
rect 52643 172940 52709 172941
rect 52643 172876 52644 172940
rect 52708 172876 52709 172940
rect 52643 172875 52709 172876
rect 54667 172940 54733 172941
rect 54667 172876 54668 172940
rect 54732 172876 54733 172940
rect 54667 172875 54733 172876
rect 55406 172805 55466 215174
rect 56326 213874 56386 221291
rect 55590 213814 56386 213874
rect 55590 172941 55650 213814
rect 73438 213741 73498 236251
rect 73622 236045 73682 282763
rect 73806 263653 73866 300035
rect 73990 291805 74050 303979
rect 74171 293028 74237 293029
rect 74171 292964 74172 293028
rect 74236 292964 74237 293028
rect 74171 292963 74237 292964
rect 73987 291804 74053 291805
rect 73987 291740 73988 291804
rect 74052 291740 74053 291804
rect 73987 291739 74053 291740
rect 74174 286634 74234 292963
rect 73990 286574 74234 286634
rect 73990 277253 74050 286574
rect 74171 286364 74237 286365
rect 74171 286300 74172 286364
rect 74236 286300 74237 286364
rect 74171 286299 74237 286300
rect 74174 282013 74234 286299
rect 74171 282012 74237 282013
rect 74171 281948 74172 282012
rect 74236 281948 74237 282012
rect 74171 281947 74237 281948
rect 73987 277252 74053 277253
rect 73987 277188 73988 277252
rect 74052 277188 74053 277252
rect 73987 277187 74053 277188
rect 73987 277116 74053 277117
rect 73987 277052 73988 277116
rect 74052 277052 74053 277116
rect 73987 277051 74053 277052
rect 73990 270453 74050 277051
rect 74171 271132 74237 271133
rect 74171 271068 74172 271132
rect 74236 271068 74237 271132
rect 74171 271067 74237 271068
rect 73987 270452 74053 270453
rect 73987 270388 73988 270452
rect 74052 270388 74053 270452
rect 73987 270387 74053 270388
rect 73987 270316 74053 270317
rect 73987 270252 73988 270316
rect 74052 270252 74053 270316
rect 73987 270251 74053 270252
rect 73803 263652 73869 263653
rect 73803 263588 73804 263652
rect 73868 263588 73869 263652
rect 73803 263587 73869 263588
rect 73806 240394 73866 263587
rect 73990 256034 74050 270251
rect 74174 256714 74234 271067
rect 74542 263517 74602 305611
rect 89104 299842 89424 299884
rect 89104 299606 89146 299842
rect 89382 299606 89424 299842
rect 89104 299564 89424 299606
rect 104718 299554 104778 300766
rect 183104 299842 183424 299884
rect 183104 299606 183146 299842
rect 183382 299606 183424 299842
rect 183104 299564 183424 299606
rect 277104 299842 277424 299884
rect 277104 299606 277146 299842
rect 277382 299606 277424 299842
rect 277104 299564 277424 299606
rect 104682 299494 104778 299554
rect 231862 294661 231922 295326
rect 231859 294660 231925 294661
rect 231859 294596 231860 294660
rect 231924 294596 231925 294660
rect 231859 294595 231925 294596
rect 136915 292212 136981 292213
rect 136915 292162 136916 292212
rect 136980 292162 136981 292212
rect 322755 291876 322756 291926
rect 322820 291876 322821 291926
rect 322755 291875 322821 291876
rect 270499 290716 270565 290717
rect 270499 290652 270500 290716
rect 270564 290652 270565 290716
rect 270499 290651 270565 290652
rect 270502 289442 270562 290651
rect 323126 289442 323186 393739
rect 323491 393124 323557 393125
rect 323491 393060 323492 393124
rect 323556 393060 323557 393124
rect 323491 393059 323557 393060
rect 323494 295562 323554 393059
rect 435740 391750 439740 396642
rect 435740 391514 435862 391750
rect 436098 391514 436182 391750
rect 436418 391514 436502 391750
rect 436738 391514 436822 391750
rect 437058 391514 437142 391750
rect 437378 391514 437462 391750
rect 437698 391514 437782 391750
rect 438018 391514 438102 391750
rect 438338 391514 438422 391750
rect 438658 391514 438742 391750
rect 438978 391514 439062 391750
rect 439298 391514 439382 391750
rect 439618 391514 439740 391750
rect 435740 361114 439740 391514
rect 435740 360878 435862 361114
rect 436098 360878 436182 361114
rect 436418 360878 436502 361114
rect 436738 360878 436822 361114
rect 437058 360878 437142 361114
rect 437378 360878 437462 361114
rect 437698 360878 437782 361114
rect 438018 360878 438102 361114
rect 438338 360878 438422 361114
rect 438658 360878 438742 361114
rect 438978 360878 439062 361114
rect 439298 360878 439382 361114
rect 439618 360878 439740 361114
rect 435740 330478 439740 360878
rect 435740 330242 435862 330478
rect 436098 330242 436182 330478
rect 436418 330242 436502 330478
rect 436738 330242 436822 330478
rect 437058 330242 437142 330478
rect 437378 330242 437462 330478
rect 437698 330242 437782 330478
rect 438018 330242 438102 330478
rect 438338 330242 438422 330478
rect 438658 330242 438742 330478
rect 438978 330242 439062 330478
rect 439298 330242 439382 330478
rect 439618 330242 439740 330478
rect 339499 327436 339565 327437
rect 339499 327372 339500 327436
rect 339564 327372 339565 327436
rect 339499 327371 339565 327372
rect 340971 327436 341037 327437
rect 340971 327372 340972 327436
rect 341036 327372 341037 327436
rect 340971 327371 341037 327372
rect 339502 314653 339562 327371
rect 340974 314925 341034 327371
rect 340971 314924 341037 314925
rect 340971 314860 340972 314924
rect 341036 314860 341037 314924
rect 340971 314859 341037 314860
rect 351827 314924 351893 314925
rect 351827 314860 351828 314924
rect 351892 314860 351893 314924
rect 351827 314859 351893 314860
rect 339499 314652 339565 314653
rect 339499 314588 339500 314652
rect 339564 314588 339565 314652
rect 339499 314587 339565 314588
rect 323126 289085 323186 289206
rect 323123 289084 323189 289085
rect 323123 289020 323124 289084
rect 323188 289020 323189 289084
rect 323123 289019 323189 289020
rect 84662 285005 84722 285126
rect 84659 285004 84725 285005
rect 84659 284940 84660 285004
rect 84724 284940 84725 285004
rect 84659 284939 84725 284940
rect 104534 284566 104594 286086
rect 351830 285362 351890 314859
rect 352563 314516 352629 314517
rect 352563 314452 352564 314516
rect 352628 314452 352629 314516
rect 352563 314451 352629 314452
rect 352566 305674 352626 314451
rect 352014 305614 352626 305674
rect 352014 293434 352074 305614
rect 435740 299842 439740 330242
rect 435740 299606 435862 299842
rect 436098 299606 436182 299842
rect 436418 299606 436502 299842
rect 436738 299606 436822 299842
rect 437058 299606 437142 299842
rect 437378 299606 437462 299842
rect 437698 299606 437782 299842
rect 438018 299606 438102 299842
rect 438338 299606 438422 299842
rect 438658 299606 438742 299842
rect 438978 299606 439062 299842
rect 439298 299606 439382 299842
rect 439618 299606 439740 299842
rect 352014 293374 352626 293434
rect 352566 286634 352626 293374
rect 352382 286574 352626 286634
rect 134894 284869 134954 285126
rect 134891 284868 134957 284869
rect 134891 284804 134892 284868
rect 134956 284804 134957 284868
rect 134891 284803 134957 284804
rect 351830 284594 351890 285126
rect 104464 284524 104784 284566
rect 104464 284288 104506 284524
rect 104742 284288 104784 284524
rect 104464 284246 104784 284288
rect 198464 284524 198784 284566
rect 198464 284288 198506 284524
rect 198742 284288 198784 284524
rect 198464 284246 198784 284288
rect 292464 284524 292784 284566
rect 351830 284534 352074 284594
rect 292464 284288 292506 284524
rect 292742 284288 292784 284524
rect 292464 284246 292784 284288
rect 104534 283562 104594 284246
rect 84475 282828 84541 282829
rect 84475 282764 84476 282828
rect 84540 282764 84541 282828
rect 84475 282763 84541 282764
rect 84478 282642 84538 282763
rect 352014 281194 352074 284534
rect 351830 281134 352074 281194
rect 138387 279428 138453 279429
rect 138387 279364 138388 279428
rect 138452 279364 138453 279428
rect 138387 279363 138453 279364
rect 138390 279293 138450 279363
rect 138387 279292 138453 279293
rect 138387 279228 138388 279292
rect 138452 279228 138453 279292
rect 138387 279227 138453 279228
rect 149059 274940 149125 274941
rect 149059 274876 149060 274940
rect 149124 274876 149125 274940
rect 149059 274875 149125 274876
rect 136915 273852 136981 273853
rect 136915 273788 136916 273852
rect 136980 273788 136981 273852
rect 136915 273787 136981 273788
rect 75459 263652 75525 263653
rect 75459 263588 75460 263652
rect 75524 263588 75525 263652
rect 75459 263587 75525 263588
rect 74539 263516 74605 263517
rect 74539 263452 74540 263516
rect 74604 263452 74605 263516
rect 74539 263451 74605 263452
rect 74542 257394 74602 263451
rect 74723 263380 74789 263381
rect 74723 263316 74724 263380
rect 74788 263316 74789 263380
rect 74723 263315 74789 263316
rect 74726 260114 74786 263315
rect 74726 260054 75154 260114
rect 75094 259522 75154 260054
rect 75462 259434 75522 263587
rect 75462 259374 76074 259434
rect 74542 257334 74786 257394
rect 74174 256654 74602 256714
rect 73990 255974 74234 256034
rect 74174 254762 74234 255974
rect 74174 253994 74234 254526
rect 74542 253994 74602 256654
rect 73990 253934 74234 253994
rect 74358 253934 74602 253994
rect 73990 245154 74050 253934
rect 74358 251954 74418 253934
rect 74358 251894 74602 251954
rect 74542 249914 74602 251894
rect 74174 249854 74602 249914
rect 74174 248554 74234 249854
rect 74174 248494 74418 248554
rect 74358 245922 74418 248494
rect 73990 245094 74602 245154
rect 74174 240394 74234 244326
rect 73806 240334 74050 240394
rect 74174 240334 74418 240394
rect 73990 239034 74050 240334
rect 73990 238974 74234 239034
rect 73987 236180 74053 236181
rect 73987 236116 73988 236180
rect 74052 236116 74053 236180
rect 73987 236115 74053 236116
rect 73619 236044 73685 236045
rect 73619 235980 73620 236044
rect 73684 235980 73685 236044
rect 73619 235979 73685 235980
rect 73435 213740 73501 213741
rect 73435 213676 73436 213740
rect 73500 213676 73501 213740
rect 73435 213675 73501 213676
rect 72147 204764 72213 204765
rect 72147 204700 72148 204764
rect 72212 204700 72213 204764
rect 72147 204699 72213 204700
rect 72150 202178 72210 204699
rect 72150 202118 72394 202178
rect 72334 192661 72394 202118
rect 72331 192660 72397 192661
rect 72331 192596 72332 192660
rect 72396 192596 72397 192660
rect 72331 192595 72397 192596
rect 72699 192524 72765 192525
rect 72699 192460 72700 192524
rect 72764 192460 72765 192524
rect 72699 192459 72765 192460
rect 72702 185317 72762 192459
rect 71963 185316 72029 185317
rect 71963 185252 71964 185316
rect 72028 185252 72029 185316
rect 71963 185251 72029 185252
rect 72699 185316 72765 185317
rect 72699 185252 72700 185316
rect 72764 185252 72765 185316
rect 72699 185251 72765 185252
rect 71966 176477 72026 185251
rect 71963 176476 72029 176477
rect 71963 176412 71964 176476
rect 72028 176412 72029 176476
rect 71963 176411 72029 176412
rect 71966 175933 72026 176411
rect 71963 175932 72029 175933
rect 71963 175868 71964 175932
rect 72028 175868 72029 175932
rect 71963 175867 72029 175868
rect 72331 175932 72397 175933
rect 72331 175868 72332 175932
rect 72396 175868 72397 175932
rect 72331 175867 72397 175868
rect 55587 172940 55653 172941
rect 55587 172876 55588 172940
rect 55652 172876 55653 172940
rect 55587 172875 55653 172876
rect 55403 172804 55469 172805
rect 55403 172740 55404 172804
rect 55468 172740 55469 172804
rect 55403 172739 55469 172740
rect 72334 169269 72394 175867
rect 73438 169541 73498 213675
rect 73622 204493 73682 235979
rect 73803 234140 73869 234141
rect 73803 234076 73804 234140
rect 73868 234076 73869 234140
rect 73803 234075 73869 234076
rect 73806 224349 73866 234075
rect 73990 228834 74050 236115
rect 74174 233869 74234 238974
rect 74358 235637 74418 240334
rect 74542 236453 74602 245094
rect 74539 236452 74605 236453
rect 74539 236388 74540 236452
rect 74604 236388 74605 236452
rect 74539 236387 74605 236388
rect 74726 236317 74786 257334
rect 75094 246514 75154 259286
rect 76014 258162 76074 259374
rect 75462 252042 75522 254526
rect 75094 246454 75338 246514
rect 74723 236316 74789 236317
rect 74723 236252 74724 236316
rect 74788 236252 74789 236316
rect 74723 236251 74789 236252
rect 74355 235636 74421 235637
rect 74355 235572 74356 235636
rect 74420 235572 74421 235636
rect 74355 235571 74421 235572
rect 74171 233868 74237 233869
rect 74171 233804 74172 233868
rect 74236 233804 74237 233868
rect 74171 233803 74237 233804
rect 73990 228774 74234 228834
rect 73803 224348 73869 224349
rect 73803 224284 73804 224348
rect 73868 224284 73869 224348
rect 73803 224283 73869 224284
rect 73803 224212 73869 224213
rect 73803 224148 73804 224212
rect 73868 224148 73869 224212
rect 73803 224147 73869 224148
rect 73806 224077 73866 224147
rect 73803 224076 73869 224077
rect 73803 224012 73804 224076
rect 73868 224012 73869 224076
rect 73803 224011 73869 224012
rect 73803 223940 73869 223941
rect 73803 223876 73804 223940
rect 73868 223876 73869 223940
rect 73803 223875 73869 223876
rect 73806 205037 73866 223875
rect 73803 205036 73869 205037
rect 73803 204972 73804 205036
rect 73868 204972 73869 205036
rect 73803 204971 73869 204972
rect 73803 204900 73869 204901
rect 73803 204836 73804 204900
rect 73868 204836 73869 204900
rect 73803 204835 73869 204836
rect 73619 204492 73685 204493
rect 73619 204428 73620 204492
rect 73684 204428 73685 204492
rect 73619 204427 73685 204428
rect 73622 203541 73682 204427
rect 73619 203540 73685 203541
rect 73619 203476 73620 203540
rect 73684 203476 73685 203540
rect 73619 203475 73685 203476
rect 73619 202180 73685 202181
rect 73619 202116 73620 202180
rect 73684 202116 73685 202180
rect 73619 202115 73685 202116
rect 73622 177973 73682 202115
rect 73619 177972 73685 177973
rect 73619 177908 73620 177972
rect 73684 177908 73685 177972
rect 73619 177907 73685 177908
rect 73806 169541 73866 204835
rect 73987 204764 74053 204765
rect 73987 204700 73988 204764
rect 74052 204700 74053 204764
rect 73987 204699 74053 204700
rect 73990 191301 74050 204699
rect 74174 195245 74234 228774
rect 74358 202181 74418 235571
rect 74539 235500 74605 235501
rect 74539 235436 74540 235500
rect 74604 235436 74605 235500
rect 74539 235435 74605 235436
rect 74542 224213 74602 235435
rect 75278 235093 75338 246454
rect 76566 241162 76626 242286
rect 75459 236452 75525 236453
rect 75459 236388 75460 236452
rect 75524 236388 75525 236452
rect 75459 236387 75525 236388
rect 75462 235501 75522 236387
rect 76014 236045 76074 240246
rect 76379 236316 76445 236317
rect 76379 236252 76380 236316
rect 76444 236252 76445 236316
rect 76379 236251 76445 236252
rect 76011 236044 76077 236045
rect 76011 235980 76012 236044
rect 76076 235980 76077 236044
rect 76011 235979 76077 235980
rect 75643 235908 75709 235909
rect 75643 235844 75644 235908
rect 75708 235844 75709 235908
rect 75643 235843 75709 235844
rect 75459 235500 75525 235501
rect 75459 235436 75460 235500
rect 75524 235436 75525 235500
rect 75459 235435 75525 235436
rect 75275 235092 75341 235093
rect 75275 235028 75276 235092
rect 75340 235028 75341 235092
rect 75275 235027 75341 235028
rect 75646 234141 75706 235843
rect 76382 235722 76442 236251
rect 76566 236181 76626 240926
rect 76934 239802 76994 243646
rect 136918 241842 136978 273787
rect 138571 269908 138637 269909
rect 138571 269844 138572 269908
rect 138636 269844 138637 269908
rect 138571 269843 138637 269844
rect 138574 269637 138634 269843
rect 138571 269636 138637 269637
rect 138571 269572 138572 269636
rect 138636 269572 138637 269636
rect 138571 269571 138637 269572
rect 138755 269636 138821 269637
rect 138755 269572 138756 269636
rect 138820 269572 138821 269636
rect 138755 269571 138821 269572
rect 138758 259981 138818 269571
rect 149062 262242 149122 274875
rect 168931 274804 168997 274805
rect 168931 274740 168932 274804
rect 168996 274740 168997 274804
rect 168931 274739 168997 274740
rect 262035 274804 262101 274805
rect 262035 274740 262036 274804
rect 262100 274740 262101 274804
rect 262035 274739 262101 274740
rect 168563 274668 168629 274669
rect 168563 274604 168564 274668
rect 168628 274604 168629 274668
rect 168563 274603 168629 274604
rect 167827 274532 167893 274533
rect 167827 274468 167828 274532
rect 167892 274468 167893 274532
rect 167827 274467 167893 274468
rect 154579 273852 154645 273853
rect 154579 273788 154580 273852
rect 154644 273788 154645 273852
rect 154579 273787 154645 273788
rect 154582 262922 154642 273787
rect 138755 259980 138821 259981
rect 138755 259916 138756 259980
rect 138820 259916 138821 259980
rect 138755 259915 138821 259916
rect 138755 250460 138821 250461
rect 138755 250396 138756 250460
rect 138820 250396 138821 250460
rect 138755 250395 138821 250396
rect 138758 245565 138818 250395
rect 144094 247962 144154 256566
rect 138755 245564 138821 245565
rect 138755 245500 138756 245564
rect 138820 245500 138821 245564
rect 138755 245499 138821 245500
rect 96067 241756 96133 241757
rect 96067 241692 96068 241756
rect 96132 241692 96133 241756
rect 96067 241691 96133 241692
rect 104899 241756 104965 241757
rect 104899 241692 104900 241756
rect 104964 241692 104965 241756
rect 104899 241691 104965 241692
rect 96070 241162 96130 241691
rect 104902 240482 104962 241691
rect 137066 241694 137346 241754
rect 76563 236180 76629 236181
rect 76563 236116 76564 236180
rect 76628 236116 76629 236180
rect 76563 236115 76629 236116
rect 76934 235909 76994 239566
rect 92571 239444 92637 239445
rect 92571 239380 92572 239444
rect 92636 239380 92637 239444
rect 92571 239379 92637 239380
rect 81350 236453 81410 236846
rect 81347 236452 81413 236453
rect 81347 236388 81348 236452
rect 81412 236388 81413 236452
rect 81347 236387 81413 236388
rect 76931 235908 76997 235909
rect 76931 235844 76932 235908
rect 76996 235844 76997 235908
rect 76931 235843 76997 235844
rect 75643 234140 75709 234141
rect 75643 234076 75644 234140
rect 75708 234076 75709 234140
rect 75643 234075 75709 234076
rect 74907 233868 74973 233869
rect 74907 233804 74908 233868
rect 74972 233804 74973 233868
rect 74907 233803 74973 233804
rect 74910 233733 74970 233803
rect 74907 233732 74973 233733
rect 74907 233668 74908 233732
rect 74972 233668 74973 233732
rect 74907 233667 74973 233668
rect 92574 226525 92634 239379
rect 100115 237948 100181 237949
rect 100115 237884 100116 237948
rect 100180 237884 100181 237948
rect 100115 237883 100181 237884
rect 100118 237762 100178 237883
rect 100118 236997 100178 237526
rect 100115 236996 100181 236997
rect 100115 236932 100116 236996
rect 100180 236932 100181 236996
rect 100115 236931 100181 236932
rect 105086 235773 105146 236166
rect 116123 235908 116189 235909
rect 116123 235844 116124 235908
rect 116188 235844 116189 235908
rect 116123 235843 116189 235844
rect 105083 235772 105149 235773
rect 105083 235708 105084 235772
rect 105148 235708 105149 235772
rect 116126 235722 116186 235843
rect 105083 235707 105149 235708
rect 133974 235637 134034 236166
rect 133971 235636 134037 235637
rect 133971 235572 133972 235636
rect 134036 235572 134037 235636
rect 133971 235571 134037 235572
rect 136366 235093 136426 236166
rect 136363 235092 136429 235093
rect 136363 235028 136364 235092
rect 136428 235028 136429 235092
rect 137286 235042 137346 241694
rect 138387 240804 138453 240805
rect 138387 240740 138388 240804
rect 138452 240740 138453 240804
rect 138387 240739 138453 240740
rect 138390 239802 138450 240739
rect 141150 239802 141210 244326
rect 141150 237677 141210 239566
rect 141147 237676 141213 237677
rect 141147 237612 141148 237676
rect 141212 237612 141213 237676
rect 141147 237611 141213 237612
rect 142990 237082 143050 245686
rect 143171 237676 143237 237677
rect 143171 237612 143172 237676
rect 143236 237674 143237 237676
rect 143236 237614 145994 237674
rect 143236 237612 143237 237614
rect 143171 237611 143237 237612
rect 145934 237082 145994 237614
rect 145198 235365 145258 236846
rect 147774 236045 147834 237526
rect 147771 236044 147837 236045
rect 147771 235980 147772 236044
rect 147836 235980 147837 236044
rect 147771 235979 147837 235980
rect 148694 235909 148754 236846
rect 167830 236181 167890 274467
rect 168195 274396 168261 274397
rect 168195 274332 168196 274396
rect 168260 274332 168261 274396
rect 168195 274331 168261 274332
rect 168198 240482 168258 274331
rect 167827 236180 167893 236181
rect 148691 235908 148757 235909
rect 148691 235844 148692 235908
rect 148756 235844 148757 235908
rect 148691 235843 148757 235844
rect 152003 235636 152069 235637
rect 152003 235572 152004 235636
rect 152068 235572 152069 235636
rect 152003 235571 152069 235572
rect 145195 235364 145261 235365
rect 145195 235300 145196 235364
rect 145260 235300 145261 235364
rect 145195 235299 145261 235300
rect 136363 235027 136429 235028
rect 137286 234764 137346 234806
rect 152006 234362 152066 235571
rect 156790 233733 156850 236166
rect 167827 236116 167828 236180
rect 167892 236116 167893 236180
rect 167827 236115 167893 236116
rect 167830 235773 167890 236115
rect 168198 236045 168258 240246
rect 168195 236044 168261 236045
rect 168195 235980 168196 236044
rect 168260 235980 168261 236044
rect 168195 235979 168261 235980
rect 167827 235772 167893 235773
rect 167827 235708 167828 235772
rect 167892 235708 167893 235772
rect 167827 235707 167893 235708
rect 158811 235636 158877 235637
rect 158811 235572 158812 235636
rect 158876 235572 158877 235636
rect 158811 235571 158877 235572
rect 158814 235042 158874 235571
rect 168566 235042 168626 274603
rect 168934 236402 168994 274739
rect 261667 274396 261733 274397
rect 261667 274332 261668 274396
rect 261732 274332 261733 274396
rect 261667 274331 261733 274332
rect 247867 273988 247933 273989
rect 247867 273924 247868 273988
rect 247932 273924 247933 273988
rect 247867 273923 247933 273924
rect 242347 273852 242413 273853
rect 242347 273788 242348 273852
rect 242412 273788 242413 273852
rect 242347 273787 242413 273788
rect 242350 272354 242410 273787
rect 242350 272294 242594 272354
rect 242534 271674 242594 272294
rect 242534 271614 242778 271674
rect 182915 269500 182981 269501
rect 182915 269436 182916 269500
rect 182980 269436 182981 269500
rect 182915 269435 182981 269436
rect 177030 236181 177090 236846
rect 177027 236180 177093 236181
rect 177027 236116 177028 236180
rect 177092 236116 177093 236180
rect 177027 236115 177093 236116
rect 156787 233732 156853 233733
rect 156787 233668 156788 233732
rect 156852 233668 156853 233732
rect 156787 233667 156853 233668
rect 174083 226932 174149 226933
rect 174083 226868 174084 226932
rect 174148 226868 174149 226932
rect 174083 226867 174149 226868
rect 116123 226796 116189 226797
rect 109134 226734 109562 226794
rect 109134 226525 109194 226734
rect 109502 226525 109562 226734
rect 116123 226732 116124 226796
rect 116188 226732 116189 226796
rect 116123 226731 116189 226732
rect 135443 226796 135509 226797
rect 135443 226732 135444 226796
rect 135508 226732 135509 226796
rect 135443 226731 135509 226732
rect 116126 226525 116186 226731
rect 135446 226525 135506 226731
rect 154763 226660 154829 226661
rect 154763 226596 154764 226660
rect 154828 226596 154829 226660
rect 154763 226595 154829 226596
rect 92571 226524 92637 226525
rect 92571 226460 92572 226524
rect 92636 226460 92637 226524
rect 92571 226459 92637 226460
rect 109131 226524 109197 226525
rect 109131 226460 109132 226524
rect 109196 226460 109197 226524
rect 109131 226459 109197 226460
rect 109499 226524 109565 226525
rect 109499 226460 109500 226524
rect 109564 226460 109565 226524
rect 109499 226459 109565 226460
rect 116123 226524 116189 226525
rect 116123 226460 116124 226524
rect 116188 226460 116189 226524
rect 116123 226459 116189 226460
rect 135443 226524 135509 226525
rect 135443 226460 135444 226524
rect 135508 226460 135509 226524
rect 135443 226459 135509 226460
rect 154766 226389 154826 226595
rect 174086 226525 174146 226867
rect 182918 226525 182978 269435
rect 219715 268412 219781 268413
rect 219715 268348 219716 268412
rect 219780 268348 219781 268412
rect 219715 268347 219781 268348
rect 193219 262156 193285 262157
rect 193219 262092 193220 262156
rect 193284 262092 193285 262156
rect 193219 262091 193285 262092
rect 193222 260882 193282 262091
rect 212542 260797 212602 262006
rect 212539 260796 212605 260797
rect 212539 260732 212540 260796
rect 212604 260732 212605 260796
rect 212539 260731 212605 260732
rect 192115 239444 192181 239445
rect 192115 239380 192116 239444
rect 192180 239380 192181 239444
rect 192115 239379 192181 239380
rect 192118 235722 192178 239379
rect 198923 238492 198989 238493
rect 198923 238428 198924 238492
rect 198988 238428 198989 238492
rect 198923 238427 198989 238428
rect 198926 236997 198986 238427
rect 219718 237813 219778 268347
rect 242718 263925 242778 271614
rect 241427 263924 241493 263925
rect 241427 263860 241428 263924
rect 241492 263860 241493 263924
rect 241427 263859 241493 263860
rect 242715 263924 242781 263925
rect 242715 263860 242716 263924
rect 242780 263860 242781 263924
rect 242715 263859 242781 263860
rect 224870 260882 224930 263366
rect 241430 262242 241490 263859
rect 247870 262242 247930 273923
rect 251179 263516 251245 263517
rect 251179 263452 251180 263516
rect 251244 263452 251245 263516
rect 251179 263451 251245 263452
rect 251182 262242 251242 263451
rect 237750 248642 237810 255206
rect 238118 246602 238178 259286
rect 231859 237948 231925 237949
rect 231859 237884 231860 237948
rect 231924 237884 231925 237948
rect 231859 237883 231925 237884
rect 219715 237812 219781 237813
rect 219715 237748 219716 237812
rect 219780 237748 219781 237812
rect 219715 237747 219781 237748
rect 231862 237082 231922 237883
rect 237750 237762 237810 239566
rect 238118 237082 238178 245686
rect 261670 237762 261730 274331
rect 262038 240482 262098 274739
rect 262403 274668 262469 274669
rect 262403 274604 262404 274668
rect 262468 274604 262469 274668
rect 262403 274603 262469 274604
rect 198923 236996 198989 236997
rect 198923 236932 198924 236996
rect 198988 236932 198989 236996
rect 198923 236931 198989 236932
rect 247134 236402 247194 237526
rect 244187 236116 244188 236166
rect 244252 236116 244253 236166
rect 244187 236115 244253 236116
rect 247134 235909 247194 236166
rect 247131 235908 247197 235909
rect 247131 235844 247132 235908
rect 247196 235844 247197 235908
rect 247131 235843 247197 235844
rect 246211 235636 246277 235637
rect 246211 235572 246212 235636
rect 246276 235572 246277 235636
rect 246211 235571 246277 235572
rect 246214 235042 246274 235571
rect 207206 234413 207266 234806
rect 207203 234412 207269 234413
rect 207203 234348 207204 234412
rect 207268 234348 207269 234412
rect 207203 234347 207269 234348
rect 246214 234274 246274 234806
rect 245626 234214 246274 234274
rect 230755 234076 230756 234126
rect 230820 234076 230821 234126
rect 230755 234075 230821 234076
rect 249894 233461 249954 234126
rect 261670 233733 261730 237526
rect 261667 233732 261733 233733
rect 261667 233668 261668 233732
rect 261732 233668 261733 233732
rect 261667 233667 261733 233668
rect 249891 233460 249957 233461
rect 249891 233396 249892 233460
rect 249956 233396 249957 233460
rect 249891 233395 249957 233396
rect 262038 233325 262098 240246
rect 262406 235042 262466 274603
rect 262587 274532 262653 274533
rect 262587 274468 262588 274532
rect 262652 274468 262653 274532
rect 262587 274467 262653 274468
rect 262590 235773 262650 274467
rect 351830 266781 351890 281134
rect 352382 280514 352442 286574
rect 352198 280454 352442 280514
rect 352198 279698 352258 280454
rect 352747 279700 352813 279701
rect 352747 279698 352748 279700
rect 352198 279638 352748 279698
rect 352198 272354 352258 279638
rect 352747 279636 352748 279638
rect 352812 279636 352813 279700
rect 352747 279635 352813 279636
rect 352014 272294 352258 272354
rect 351827 266780 351893 266781
rect 351827 266716 351828 266780
rect 351892 266716 351893 266780
rect 351827 266715 351893 266716
rect 352014 266645 352074 272294
rect 435740 269206 439740 299606
rect 435740 268970 435862 269206
rect 436098 268970 436182 269206
rect 436418 268970 436502 269206
rect 436738 268970 436822 269206
rect 437058 268970 437142 269206
rect 437378 268970 437462 269206
rect 437698 268970 437782 269206
rect 438018 268970 438102 269206
rect 438338 268970 438422 269206
rect 438658 268970 438742 269206
rect 438978 268970 439062 269206
rect 439298 268970 439382 269206
rect 439618 268970 439740 269206
rect 352011 266644 352077 266645
rect 352011 266580 352012 266644
rect 352076 266580 352077 266644
rect 352011 266579 352077 266580
rect 356394 261414 358330 261474
rect 295523 239852 295589 239853
rect 295523 239802 295524 239852
rect 295588 239802 295589 239852
rect 283195 239444 283261 239445
rect 283195 239380 283196 239444
rect 283260 239380 283261 239444
rect 283195 239379 283261 239380
rect 264798 236997 264858 237526
rect 264795 236996 264861 236997
rect 264795 236932 264796 236996
rect 264860 236932 264861 236996
rect 264795 236931 264861 236932
rect 262587 235772 262653 235773
rect 262587 235708 262588 235772
rect 262652 235708 262653 235772
rect 262587 235707 262653 235708
rect 283198 234413 283258 239379
rect 290003 238492 290069 238493
rect 290003 238428 290004 238492
rect 290068 238428 290069 238492
rect 290003 238427 290069 238428
rect 290006 237082 290066 238427
rect 295526 235722 295586 239566
rect 283195 234412 283261 234413
rect 283195 234362 283196 234412
rect 283260 234362 283261 234412
rect 262035 233324 262101 233325
rect 262035 233260 262036 233324
rect 262100 233260 262101 233324
rect 262035 233259 262101 233260
rect 239587 232508 239653 232509
rect 239587 232444 239588 232508
rect 239652 232444 239653 232508
rect 239587 232443 239653 232444
rect 351643 232508 351709 232509
rect 351643 232444 351644 232508
rect 351708 232444 351709 232508
rect 351643 232443 351709 232444
rect 351827 232508 351893 232509
rect 351827 232444 351828 232508
rect 351892 232444 351893 232508
rect 351827 232443 351893 232444
rect 185859 227068 185925 227069
rect 185859 227004 185860 227068
rect 185924 227004 185925 227068
rect 185859 227003 185925 227004
rect 193035 227068 193101 227069
rect 193035 227004 193036 227068
rect 193100 227004 193101 227068
rect 193035 227003 193101 227004
rect 185862 226661 185922 227003
rect 185859 226660 185925 226661
rect 185859 226596 185860 226660
rect 185924 226596 185925 226660
rect 185859 226595 185925 226596
rect 174083 226524 174149 226525
rect 174083 226460 174084 226524
rect 174148 226460 174149 226524
rect 174083 226459 174149 226460
rect 178683 226524 178749 226525
rect 178683 226460 178684 226524
rect 178748 226460 178749 226524
rect 178683 226459 178749 226460
rect 182915 226524 182981 226525
rect 182915 226460 182916 226524
rect 182980 226460 182981 226524
rect 182915 226459 182981 226460
rect 154763 226388 154829 226389
rect 154763 226324 154764 226388
rect 154828 226324 154829 226388
rect 154763 226323 154829 226324
rect 74539 224212 74605 224213
rect 74539 224148 74540 224212
rect 74604 224148 74605 224212
rect 74539 224147 74605 224148
rect 74539 224076 74605 224077
rect 74539 224012 74540 224076
rect 74604 224012 74605 224076
rect 74539 224011 74605 224012
rect 74542 204901 74602 224011
rect 104464 223252 104784 223294
rect 104464 223016 104506 223252
rect 104742 223016 104784 223252
rect 104464 222974 104784 223016
rect 178686 214642 178746 226459
rect 193038 226114 193098 227003
rect 193219 226524 193285 226525
rect 193219 226460 193220 226524
rect 193284 226460 193285 226524
rect 193219 226459 193285 226460
rect 193222 226114 193282 226459
rect 193038 226054 193282 226114
rect 198464 223252 198784 223294
rect 198464 223016 198506 223252
rect 198742 223016 198784 223252
rect 198464 222974 198784 223016
rect 147035 208300 147101 208301
rect 147035 208236 147036 208300
rect 147100 208236 147101 208300
rect 147035 208235 147101 208236
rect 89104 207934 89424 207976
rect 89104 207698 89146 207934
rect 89382 207698 89424 207934
rect 89104 207656 89424 207698
rect 74539 204900 74605 204901
rect 74539 204836 74540 204900
rect 74604 204836 74605 204900
rect 74539 204835 74605 204836
rect 134707 204836 134708 204886
rect 134772 204836 134773 204886
rect 134707 204835 134773 204836
rect 74539 204764 74605 204765
rect 74539 204700 74540 204764
rect 74604 204700 74605 204764
rect 74539 204699 74605 204700
rect 74355 202180 74421 202181
rect 74355 202116 74356 202180
rect 74420 202116 74421 202180
rect 74355 202115 74421 202116
rect 74542 199189 74602 204699
rect 84659 204492 84725 204493
rect 84659 204442 84660 204492
rect 84724 204442 84725 204492
rect 74539 199188 74605 199189
rect 74539 199124 74540 199188
rect 74604 199124 74605 199188
rect 74539 199123 74605 199124
rect 74542 195245 74602 199123
rect 136918 198237 136978 198766
rect 136915 198236 136981 198237
rect 136915 198172 136916 198236
rect 136980 198172 136981 198236
rect 136915 198171 136981 198172
rect 74171 195244 74237 195245
rect 74171 195180 74172 195244
rect 74236 195180 74237 195244
rect 74171 195179 74237 195180
rect 74539 195244 74605 195245
rect 74539 195180 74540 195244
rect 74604 195180 74605 195244
rect 74539 195179 74605 195180
rect 74355 195108 74421 195109
rect 74355 195044 74356 195108
rect 74420 195044 74421 195108
rect 74355 195043 74421 195044
rect 74539 195108 74605 195109
rect 74539 195044 74540 195108
rect 74604 195044 74605 195108
rect 74539 195043 74605 195044
rect 73987 191300 74053 191301
rect 73987 191236 73988 191300
rect 74052 191236 74053 191300
rect 73987 191235 74053 191236
rect 73990 185589 74050 191235
rect 73987 185588 74053 185589
rect 73987 185524 73988 185588
rect 74052 185524 74053 185588
rect 73987 185523 74053 185524
rect 73987 185452 74053 185453
rect 73987 185388 73988 185452
rect 74052 185388 74053 185452
rect 73987 185387 74053 185388
rect 73435 169540 73501 169541
rect 73435 169476 73436 169540
rect 73500 169476 73501 169540
rect 73435 169475 73501 169476
rect 73803 169540 73869 169541
rect 73803 169476 73804 169540
rect 73868 169476 73869 169540
rect 73803 169475 73869 169476
rect 72331 169268 72397 169269
rect 72331 169204 72332 169268
rect 72396 169204 72397 169268
rect 72331 169203 72397 169204
rect 73438 168314 73498 169475
rect 73438 168254 73682 168314
rect 48966 162605 49026 162726
rect 48963 162604 49029 162605
rect 48963 162540 48964 162604
rect 49028 162540 49029 162604
rect 48963 162539 49029 162540
rect 49147 158388 49213 158389
rect 49147 158324 49148 158388
rect 49212 158324 49213 158388
rect 49147 158323 49213 158324
rect 49150 158202 49210 158323
rect 49147 152948 49213 152949
rect 49147 152884 49148 152948
rect 49212 152884 49213 152948
rect 49147 152883 49213 152884
rect 49150 152762 49210 152883
rect 49147 149004 49213 149005
rect 49147 148940 49148 149004
rect 49212 148940 49213 149004
rect 49147 148939 49213 148940
rect 49150 148682 49210 148939
rect 5000 146426 5122 146662
rect 5358 146426 5442 146662
rect 5678 146426 5762 146662
rect 5998 146426 6082 146662
rect 6318 146426 6402 146662
rect 6638 146426 6722 146662
rect 6958 146426 7042 146662
rect 7278 146426 7362 146662
rect 7598 146426 7682 146662
rect 7918 146426 8002 146662
rect 8238 146426 8322 146662
rect 8558 146426 8642 146662
rect 8878 146426 9000 146662
rect 5000 116026 9000 146426
rect 73622 143834 73682 168254
rect 73438 143774 73682 143834
rect 52643 139620 52709 139621
rect 52643 139556 52644 139620
rect 52708 139556 52709 139620
rect 52643 139555 52709 139556
rect 54851 139620 54917 139621
rect 54851 139556 54852 139620
rect 54916 139556 54917 139620
rect 54851 139555 54917 139556
rect 5000 115790 5122 116026
rect 5358 115790 5442 116026
rect 5678 115790 5762 116026
rect 5998 115790 6082 116026
rect 6318 115790 6402 116026
rect 6638 115790 6722 116026
rect 6958 115790 7042 116026
rect 7278 115790 7362 116026
rect 7598 115790 7682 116026
rect 7918 115790 8002 116026
rect 8238 115790 8322 116026
rect 8558 115790 8642 116026
rect 8878 115790 9000 116026
rect 5000 85390 9000 115790
rect 52646 113101 52706 139555
rect 54667 122076 54733 122077
rect 54667 122012 54668 122076
rect 54732 122012 54733 122076
rect 54667 122011 54733 122012
rect 52643 113100 52709 113101
rect 52643 113036 52644 113100
rect 52708 113036 52709 113100
rect 52643 113035 52709 113036
rect 5000 85154 5122 85390
rect 5358 85154 5442 85390
rect 5678 85154 5762 85390
rect 5998 85154 6082 85390
rect 6318 85154 6402 85390
rect 6638 85154 6722 85390
rect 6958 85154 7042 85390
rect 7278 85154 7362 85390
rect 7598 85154 7682 85390
rect 7918 85154 8002 85390
rect 8238 85154 8322 85390
rect 8558 85154 8642 85390
rect 8878 85154 9000 85390
rect 5000 54754 9000 85154
rect 52646 77877 52706 113035
rect 54670 77877 54730 122011
rect 54854 117181 54914 139555
rect 73438 139485 73498 143774
rect 73806 143154 73866 169475
rect 73990 168314 74050 185387
rect 74171 173756 74237 173757
rect 74171 173692 74172 173756
rect 74236 173692 74237 173756
rect 74358 173754 74418 195043
rect 74542 185725 74602 195043
rect 138019 194700 138085 194701
rect 138019 194636 138020 194700
rect 138084 194636 138085 194700
rect 138019 194635 138085 194636
rect 138022 194242 138082 194635
rect 104464 192616 104784 192658
rect 104464 192380 104506 192616
rect 104742 192380 104784 192616
rect 104464 192338 104784 192380
rect 74539 185724 74605 185725
rect 74539 185660 74540 185724
rect 74604 185660 74605 185724
rect 74539 185659 74605 185660
rect 74539 185588 74605 185589
rect 74539 185524 74540 185588
rect 74604 185524 74605 185588
rect 74539 185523 74605 185524
rect 74542 174434 74602 185523
rect 147038 181237 147098 208235
rect 164883 198916 164949 198917
rect 164883 198914 164884 198916
rect 164518 198854 164884 198914
rect 164518 197642 164578 198854
rect 164883 198852 164884 198854
rect 164948 198852 164949 198916
rect 164883 198851 164949 198852
rect 176659 198916 176725 198917
rect 176659 198852 176660 198916
rect 176724 198852 176725 198916
rect 176659 198851 176725 198852
rect 176662 198322 176722 198851
rect 178686 195602 178746 211006
rect 183104 207934 183424 207976
rect 183104 207698 183146 207934
rect 183382 207698 183424 207934
rect 183104 207656 183424 207698
rect 239590 204442 239650 232443
rect 292464 223252 292784 223294
rect 292464 223016 292506 223252
rect 292742 223016 292784 223252
rect 292464 222974 292784 223016
rect 322758 216597 322818 217806
rect 322755 216596 322821 216597
rect 322755 216532 322756 216596
rect 322820 216532 322821 216596
rect 322755 216531 322821 216532
rect 277104 207934 277424 207976
rect 277104 207698 277146 207934
rect 277382 207698 277424 207934
rect 277104 207656 277424 207698
rect 242715 204628 242781 204629
rect 242715 204564 242716 204628
rect 242780 204564 242781 204628
rect 242715 204563 242781 204564
rect 237379 204356 237445 204357
rect 237379 204292 237380 204356
rect 237444 204292 237445 204356
rect 237379 204291 237445 204292
rect 230758 197557 230818 198766
rect 230755 197556 230821 197557
rect 230755 197492 230756 197556
rect 230820 197492 230821 197556
rect 230755 197491 230821 197492
rect 230755 194972 230821 194973
rect 230755 194908 230756 194972
rect 230820 194908 230821 194972
rect 230755 194907 230821 194908
rect 178686 186082 178746 194686
rect 230758 194242 230818 194907
rect 198464 192616 198784 192658
rect 198464 192380 198506 192616
rect 198742 192380 198784 192616
rect 198464 192338 198784 192380
rect 174819 182052 174885 182053
rect 174819 181988 174820 182052
rect 174884 181988 174885 182052
rect 174819 181987 174885 181988
rect 147035 181236 147101 181237
rect 147035 181172 147036 181236
rect 147100 181172 147101 181236
rect 147035 181171 147101 181172
rect 169115 181100 169181 181101
rect 169115 181036 169116 181100
rect 169180 181036 169181 181100
rect 169115 181035 169181 181036
rect 168563 180964 168629 180965
rect 168563 180900 168564 180964
rect 168628 180900 168629 180964
rect 168563 180899 168629 180900
rect 167643 180828 167709 180829
rect 167643 180764 167644 180828
rect 167708 180764 167709 180828
rect 167643 180763 167709 180764
rect 147955 180556 148021 180557
rect 147955 180492 147956 180556
rect 148020 180492 148021 180556
rect 147955 180491 148021 180492
rect 75459 177972 75525 177973
rect 75459 177908 75460 177972
rect 75524 177908 75525 177972
rect 75459 177907 75525 177908
rect 74542 174374 74786 174434
rect 74358 173694 74602 173754
rect 74171 173691 74237 173692
rect 74174 169677 74234 173691
rect 74171 169676 74237 169677
rect 74171 169612 74172 169676
rect 74236 169612 74237 169676
rect 74171 169611 74237 169612
rect 74542 168314 74602 173694
rect 74726 169405 74786 174374
rect 75462 169813 75522 177907
rect 75459 169812 75525 169813
rect 75459 169748 75460 169812
rect 75524 169748 75525 169812
rect 75459 169747 75525 169748
rect 76747 169812 76813 169813
rect 76747 169748 76748 169812
rect 76812 169748 76813 169812
rect 76747 169747 76813 169748
rect 76379 169676 76445 169677
rect 76379 169612 76380 169676
rect 76444 169612 76445 169676
rect 76379 169611 76445 169612
rect 75459 169540 75525 169541
rect 75459 169476 75460 169540
rect 75524 169476 75525 169540
rect 75459 169475 75525 169476
rect 74723 169404 74789 169405
rect 74723 169340 74724 169404
rect 74788 169340 74789 169404
rect 74723 169339 74789 169340
rect 73990 168254 74234 168314
rect 74542 168254 74970 168314
rect 74174 156842 74234 168254
rect 74910 163554 74970 168254
rect 75462 165594 75522 169475
rect 75643 169404 75709 169405
rect 75643 169340 75644 169404
rect 75708 169340 75709 169404
rect 75643 169339 75709 169340
rect 75646 166274 75706 169339
rect 75827 169268 75893 169269
rect 75827 169204 75828 169268
rect 75892 169204 75893 169268
rect 75827 169203 75893 169204
rect 75830 167634 75890 169203
rect 75830 167574 76074 167634
rect 76014 166954 76074 167574
rect 76014 166894 76258 166954
rect 75646 166214 76074 166274
rect 75462 165534 75890 165594
rect 74726 163494 74970 163554
rect 74726 156074 74786 163494
rect 75462 161514 75522 164766
rect 74910 161454 75522 161514
rect 74910 159474 74970 161454
rect 75830 160834 75890 165534
rect 75462 160774 75890 160834
rect 75462 160242 75522 160774
rect 76014 159474 76074 166214
rect 74910 159414 75338 159474
rect 75278 158202 75338 159414
rect 75646 159414 76074 159474
rect 75646 157434 75706 159414
rect 76198 158794 76258 166894
rect 74358 156014 74786 156074
rect 74910 157374 75706 157434
rect 75830 158734 76258 158794
rect 74910 156074 74970 157374
rect 74910 156014 75338 156074
rect 74358 152762 74418 156014
rect 74358 151994 74418 152526
rect 75278 151994 75338 156014
rect 73990 151934 74418 151994
rect 74726 151934 75338 151994
rect 73990 143834 74050 151934
rect 74726 151314 74786 151934
rect 75462 151314 75522 156606
rect 74542 151254 74786 151314
rect 74910 151254 75522 151314
rect 74542 150634 74602 151254
rect 74910 150634 74970 151254
rect 74358 150574 74602 150634
rect 74726 150574 74970 150634
rect 74358 146554 74418 150574
rect 74726 148682 74786 150574
rect 75830 149954 75890 158734
rect 76382 158114 76442 169611
rect 76750 165002 76810 169747
rect 147958 169269 148018 180491
rect 144091 169268 144157 169269
rect 144091 169204 144092 169268
rect 144156 169204 144157 169268
rect 144091 169203 144157 169204
rect 147955 169268 148021 169269
rect 147955 169204 147956 169268
rect 148020 169204 148021 169268
rect 147955 169203 148021 169204
rect 76750 160242 76810 162726
rect 144094 160922 144154 169203
rect 76382 158054 76626 158114
rect 76566 157573 76626 158054
rect 76563 157572 76629 157573
rect 76563 157508 76564 157572
rect 76628 157508 76629 157572
rect 76563 157507 76629 157508
rect 76747 157164 76813 157165
rect 76747 157100 76748 157164
rect 76812 157100 76813 157164
rect 76747 157099 76813 157100
rect 76382 156074 76442 156606
rect 75278 149894 75890 149954
rect 76014 156014 76442 156074
rect 76014 149954 76074 156014
rect 76750 154802 76810 157099
rect 76014 149894 76442 149954
rect 74726 146554 74786 148446
rect 75278 146554 75338 149894
rect 76382 148594 76442 149894
rect 76563 148596 76629 148597
rect 76563 148594 76564 148596
rect 76382 148534 76564 148594
rect 76563 148532 76564 148534
rect 76628 148532 76629 148596
rect 76563 148531 76629 148532
rect 74358 146494 74602 146554
rect 74726 146494 74970 146554
rect 75278 146494 75706 146554
rect 74542 145962 74602 146494
rect 74910 145874 74970 146494
rect 74910 145814 75338 145874
rect 74910 144514 74970 145046
rect 74542 144454 74970 144514
rect 73990 143774 74418 143834
rect 73806 143094 74004 143154
rect 73803 142476 73869 142477
rect 73803 142412 73804 142476
rect 73868 142412 73869 142476
rect 73803 142411 73869 142412
rect 73435 139484 73501 139485
rect 73435 139420 73436 139484
rect 73500 139420 73501 139484
rect 73435 139419 73501 139420
rect 73619 137172 73685 137173
rect 73619 137108 73620 137172
rect 73684 137108 73685 137172
rect 73619 137107 73685 137108
rect 55219 134452 55285 134453
rect 55219 134388 55220 134452
rect 55284 134388 55285 134452
rect 55219 134387 55285 134388
rect 55035 122076 55101 122077
rect 55035 122012 55036 122076
rect 55100 122074 55101 122076
rect 55222 122074 55282 134387
rect 55403 132412 55469 132413
rect 55403 132348 55404 132412
rect 55468 132348 55469 132412
rect 55403 132347 55469 132348
rect 55406 127245 55466 132347
rect 73622 128194 73682 137107
rect 73806 137034 73866 142411
rect 73944 142069 74004 143094
rect 74358 142477 74418 143774
rect 74355 142476 74421 142477
rect 74355 142412 74356 142476
rect 74420 142412 74421 142476
rect 74355 142411 74421 142412
rect 74542 142205 74602 144454
rect 74910 142477 74970 143686
rect 74907 142476 74973 142477
rect 74907 142412 74908 142476
rect 74972 142412 74973 142476
rect 74907 142411 74973 142412
rect 74539 142204 74605 142205
rect 74539 142140 74540 142204
rect 74604 142140 74605 142204
rect 74539 142139 74605 142140
rect 75278 142069 75338 145814
rect 75646 142205 75706 146494
rect 77118 145282 77178 153206
rect 98275 144244 98341 144245
rect 98275 144180 98276 144244
rect 98340 144180 98341 144244
rect 98275 144179 98341 144180
rect 142251 144244 142317 144245
rect 142251 144180 142252 144244
rect 142316 144180 142317 144244
rect 142251 144179 142317 144180
rect 76931 144108 76997 144109
rect 76931 144044 76932 144108
rect 76996 144044 76997 144108
rect 76931 144043 76997 144044
rect 75643 142204 75709 142205
rect 75643 142140 75644 142204
rect 75708 142140 75709 142204
rect 75643 142139 75709 142140
rect 73944 142068 74053 142069
rect 73944 142006 73988 142068
rect 73987 142004 73988 142006
rect 74052 142004 74053 142068
rect 73987 142003 74053 142004
rect 74539 142068 74605 142069
rect 74539 142004 74540 142068
rect 74604 142004 74605 142068
rect 74539 142003 74605 142004
rect 75275 142068 75341 142069
rect 75275 142004 75276 142068
rect 75340 142004 75341 142068
rect 75275 142003 75341 142004
rect 74355 141796 74421 141797
rect 74355 141732 74356 141796
rect 74420 141732 74421 141796
rect 74355 141731 74421 141732
rect 73806 136974 74050 137034
rect 73254 128134 73682 128194
rect 55403 127244 55469 127245
rect 55403 127180 55404 127244
rect 55468 127180 55469 127244
rect 55403 127179 55469 127180
rect 55100 122014 55282 122074
rect 55100 122012 55101 122014
rect 55035 122011 55101 122012
rect 54851 117180 54917 117181
rect 54851 117116 54852 117180
rect 54916 117116 54917 117180
rect 54851 117115 54917 117116
rect 54854 78013 54914 117115
rect 54851 78012 54917 78013
rect 54851 77948 54852 78012
rect 54916 77948 54917 78012
rect 54851 77947 54917 77948
rect 55406 77877 55466 127179
rect 73254 124797 73314 128134
rect 73251 124796 73317 124797
rect 73251 124732 73252 124796
rect 73316 124732 73317 124796
rect 73251 124731 73317 124732
rect 73251 124660 73317 124661
rect 73251 124596 73252 124660
rect 73316 124596 73317 124660
rect 73251 124595 73317 124596
rect 73254 117314 73314 124595
rect 73990 117994 74050 136974
rect 73990 117934 74188 117994
rect 73803 117724 73869 117725
rect 73803 117660 73804 117724
rect 73868 117660 73869 117724
rect 74128 117722 74188 117934
rect 74358 117725 74418 141731
rect 74355 117724 74421 117725
rect 74128 117662 74234 117722
rect 73803 117659 73869 117660
rect 73254 117254 73682 117314
rect 73622 98277 73682 117254
rect 73806 109565 73866 117659
rect 73803 109564 73869 109565
rect 73803 109500 73804 109564
rect 73868 109500 73869 109564
rect 73803 109499 73869 109500
rect 74174 102085 74234 117662
rect 74355 117660 74356 117724
rect 74420 117660 74421 117724
rect 74355 117659 74421 117660
rect 74542 112829 74602 142003
rect 76014 141933 76074 143006
rect 76011 141932 76077 141933
rect 76011 141868 76012 141932
rect 76076 141868 76077 141932
rect 76011 141867 76077 141868
rect 76934 141797 76994 144043
rect 98278 143922 98338 144179
rect 142067 144108 142133 144109
rect 142067 144044 142068 144108
rect 142132 144044 142133 144108
rect 142067 144043 142133 144044
rect 110419 143292 110485 143293
rect 110419 143242 110420 143292
rect 110484 143242 110485 143292
rect 136915 143292 136981 143293
rect 136915 143242 136916 143292
rect 136980 143242 136981 143292
rect 89627 142884 89693 142885
rect 89627 142820 89628 142884
rect 89692 142820 89693 142884
rect 89627 142819 89693 142820
rect 76931 141796 76997 141797
rect 76931 141732 76932 141796
rect 76996 141732 76997 141796
rect 76931 141731 76997 141732
rect 89630 131594 89690 142819
rect 142070 142069 142130 144043
rect 142254 142205 142314 144179
rect 142438 142341 142498 144366
rect 142435 142340 142501 142341
rect 142435 142276 142436 142340
rect 142500 142276 142501 142340
rect 142435 142275 142501 142276
rect 144094 142205 144154 150486
rect 151822 142341 151882 143006
rect 151819 142340 151885 142341
rect 151819 142276 151820 142340
rect 151884 142276 151885 142340
rect 151819 142275 151885 142276
rect 167646 142205 167706 180763
rect 167827 180556 167893 180557
rect 167827 180492 167828 180556
rect 167892 180492 167893 180556
rect 167827 180491 167893 180492
rect 142251 142204 142317 142205
rect 142251 142140 142252 142204
rect 142316 142140 142317 142204
rect 142251 142139 142317 142140
rect 144091 142204 144157 142205
rect 144091 142140 144092 142204
rect 144156 142140 144157 142204
rect 144091 142139 144157 142140
rect 167643 142204 167709 142205
rect 167643 142140 167644 142204
rect 167708 142140 167709 142204
rect 167643 142139 167709 142140
rect 142067 142068 142133 142069
rect 142067 142004 142068 142068
rect 142132 142004 142133 142068
rect 142067 142003 142133 142004
rect 105083 141932 105149 141933
rect 105083 141882 105084 141932
rect 105148 141882 105149 141932
rect 167830 141797 167890 180491
rect 168566 143154 168626 180899
rect 168566 143094 168994 143154
rect 167827 141796 167893 141797
rect 167827 141732 167828 141796
rect 167892 141732 167893 141796
rect 167827 141731 167893 141732
rect 168934 141114 168994 143094
rect 168714 141054 168994 141114
rect 169118 142474 169178 181035
rect 169483 180692 169549 180693
rect 169483 180628 169484 180692
rect 169548 180628 169549 180692
rect 169483 180627 169549 180628
rect 169486 145282 169546 180627
rect 174822 179962 174882 181987
rect 178318 178245 178378 182446
rect 228915 182052 228981 182053
rect 228915 181988 228916 182052
rect 228980 181988 228981 182052
rect 228915 181987 228981 181988
rect 228918 181322 228978 181987
rect 178315 178244 178381 178245
rect 178315 178180 178316 178244
rect 178380 178180 178381 178244
rect 178315 178179 178381 178180
rect 182915 175796 182981 175797
rect 182915 175732 182916 175796
rect 182980 175732 182981 175796
rect 182915 175731 182981 175732
rect 169486 143242 169546 145046
rect 169854 143094 170134 143154
rect 169854 142474 169914 143094
rect 169118 142414 169914 142474
rect 137283 140236 137284 140286
rect 137348 140236 137349 140286
rect 137283 140235 137349 140236
rect 169118 139893 169178 142414
rect 147771 139892 147837 139893
rect 147771 139828 147772 139892
rect 147836 139828 147837 139892
rect 147771 139827 147837 139828
rect 148507 139892 148573 139893
rect 148507 139828 148508 139892
rect 148572 139828 148573 139892
rect 148507 139827 148573 139828
rect 169115 139892 169181 139893
rect 169115 139828 169116 139892
rect 169180 139828 169181 139892
rect 169115 139827 169181 139828
rect 84662 131534 89690 131594
rect 84662 127517 84722 131534
rect 84659 127516 84725 127517
rect 84659 127452 84660 127516
rect 84724 127452 84725 127516
rect 84659 127451 84725 127452
rect 89104 116026 89424 116068
rect 89104 115790 89146 116026
rect 89382 115790 89424 116026
rect 89104 115748 89424 115790
rect 147774 113237 147834 139827
rect 148510 117402 148570 139827
rect 182918 132549 182978 175731
rect 219715 175524 219781 175525
rect 219715 175460 219716 175524
rect 219780 175460 219781 175524
rect 219715 175459 219781 175460
rect 187147 145196 187213 145197
rect 187147 145132 187148 145196
rect 187212 145132 187213 145196
rect 187147 145131 187213 145132
rect 187150 144602 187210 145131
rect 197635 144652 197701 144653
rect 197635 144588 197636 144652
rect 197700 144588 197701 144652
rect 197635 144587 197701 144588
rect 197638 143973 197698 144587
rect 197635 143972 197701 143973
rect 197635 143908 197636 143972
rect 197700 143908 197701 143972
rect 197635 143907 197701 143908
rect 219718 142069 219778 175459
rect 237011 167092 237077 167093
rect 237011 167028 237012 167092
rect 237076 167028 237077 167092
rect 237011 167027 237077 167028
rect 237014 166954 237074 167027
rect 237382 166954 237442 204291
rect 239590 204164 239650 204206
rect 242718 202045 242778 204563
rect 322755 204156 322756 204206
rect 322820 204156 322821 204206
rect 322755 204155 322821 204156
rect 242715 202044 242781 202045
rect 242715 201980 242716 202044
rect 242780 201980 242781 202044
rect 242715 201979 242781 201980
rect 322755 198716 322756 198766
rect 322820 198716 322821 198766
rect 322755 198715 322821 198716
rect 270502 197557 270562 198086
rect 270499 197556 270565 197557
rect 270499 197492 270500 197556
rect 270564 197492 270565 197556
rect 270499 197491 270565 197492
rect 322755 194564 322821 194565
rect 322755 194500 322756 194564
rect 322820 194500 322821 194564
rect 322755 194499 322821 194500
rect 322758 194242 322818 194499
rect 292464 192616 292784 192658
rect 242531 192524 242597 192525
rect 242531 192460 242532 192524
rect 242596 192460 242597 192524
rect 242531 192459 242597 192460
rect 242534 185994 242594 192459
rect 292464 192380 292506 192616
rect 292742 192380 292784 192616
rect 292464 192338 292784 192380
rect 242534 185934 242778 185994
rect 242718 183141 242778 185934
rect 351646 184093 351706 232443
rect 351830 191434 351890 232443
rect 358270 216461 358330 261414
rect 435740 238570 439740 268970
rect 435740 238334 435862 238570
rect 436098 238334 436182 238570
rect 436418 238334 436502 238570
rect 436738 238334 436822 238570
rect 437058 238334 437142 238570
rect 437378 238334 437462 238570
rect 437698 238334 437782 238570
rect 438018 238334 438102 238570
rect 438338 238334 438422 238570
rect 438658 238334 438742 238570
rect 438978 238334 439062 238570
rect 439298 238334 439382 238570
rect 439618 238334 439740 238570
rect 380840 223252 381160 223294
rect 380840 223016 380882 223252
rect 381118 223016 381160 223252
rect 380840 222974 381160 223016
rect 358267 216460 358333 216461
rect 358267 216396 358268 216460
rect 358332 216396 358333 216460
rect 358267 216395 358333 216396
rect 435740 207934 439740 238334
rect 435740 207698 435862 207934
rect 436098 207698 436182 207934
rect 436418 207698 436502 207934
rect 436738 207698 436822 207934
rect 437058 207698 437142 207934
rect 437378 207698 437462 207934
rect 437698 207698 437782 207934
rect 438018 207698 438102 207934
rect 438338 207698 438422 207934
rect 438658 207698 438742 207934
rect 438978 207698 439062 207934
rect 439298 207698 439382 207934
rect 439618 207698 439740 207934
rect 352747 191436 352813 191437
rect 352747 191434 352748 191436
rect 351830 191374 352748 191434
rect 351643 184092 351709 184093
rect 351643 184028 351644 184092
rect 351708 184028 351709 184092
rect 351643 184027 351709 184028
rect 242715 183140 242781 183141
rect 242715 183076 242716 183140
rect 242780 183076 242781 183140
rect 242715 183075 242781 183076
rect 271422 182189 271482 182446
rect 322942 182189 323002 183126
rect 271419 182188 271485 182189
rect 271419 182124 271420 182188
rect 271484 182124 271485 182188
rect 271419 182123 271485 182124
rect 322939 182188 323005 182189
rect 322939 182124 322940 182188
rect 323004 182124 323005 182188
rect 322939 182123 323005 182124
rect 271419 182052 271485 182053
rect 271419 181988 271420 182052
rect 271484 181988 271485 182052
rect 322939 182052 323005 182053
rect 322939 182002 322940 182052
rect 323004 182002 323005 182052
rect 271419 181987 271485 181988
rect 261667 180828 261733 180829
rect 261667 180764 261668 180828
rect 261732 180764 261733 180828
rect 261667 180763 261733 180764
rect 242347 180692 242413 180693
rect 242347 180628 242348 180692
rect 242412 180628 242413 180692
rect 242347 180627 242413 180628
rect 241795 180148 241861 180149
rect 241795 180084 241796 180148
rect 241860 180084 241861 180148
rect 241795 180083 241861 180084
rect 241798 169082 241858 180083
rect 242350 168402 242410 180627
rect 242899 180012 242965 180013
rect 242899 179948 242900 180012
rect 242964 179948 242965 180012
rect 242899 179947 242965 179948
rect 242902 169674 242962 179947
rect 242902 169614 243330 169674
rect 243270 168402 243330 169614
rect 237014 166894 237442 166954
rect 237382 160922 237442 164086
rect 237750 156842 237810 164766
rect 238118 157522 238178 165446
rect 236830 147917 236890 153206
rect 237382 149894 238178 149954
rect 237382 148682 237442 149894
rect 236827 147916 236893 147917
rect 236827 147852 236828 147916
rect 236892 147852 236893 147916
rect 236827 147851 236893 147852
rect 237195 147916 237261 147917
rect 237195 147852 237196 147916
rect 237260 147914 237261 147916
rect 238118 147914 238178 149894
rect 237260 147854 237994 147914
rect 238118 147854 238362 147914
rect 237260 147852 237261 147854
rect 237195 147851 237261 147852
rect 237934 147234 237994 147854
rect 237934 147174 238178 147234
rect 236091 144108 236157 144109
rect 236091 144044 236092 144108
rect 236156 144044 236157 144108
rect 237566 144106 237626 147086
rect 237566 144046 237810 144106
rect 236091 144043 236157 144044
rect 219715 142068 219781 142069
rect 219715 142004 219716 142068
rect 219780 142004 219781 142068
rect 219715 142003 219781 142004
rect 230755 141932 230821 141933
rect 230755 141868 230756 141932
rect 230820 141868 230821 141932
rect 236094 141882 236154 144043
rect 237750 141882 237810 144046
rect 238118 142205 238178 147174
rect 238302 142477 238362 147854
rect 238299 142476 238365 142477
rect 238299 142412 238300 142476
rect 238364 142412 238365 142476
rect 238299 142411 238365 142412
rect 242531 142476 242597 142477
rect 242531 142412 242532 142476
rect 242596 142412 242597 142476
rect 242531 142411 242597 142412
rect 238115 142204 238181 142205
rect 238115 142140 238116 142204
rect 238180 142140 238181 142204
rect 238115 142139 238181 142140
rect 230755 141867 230821 141868
rect 230758 140522 230818 141867
rect 241979 141796 242045 141797
rect 241979 141732 241980 141796
rect 242044 141732 242045 141796
rect 241979 141731 242045 141732
rect 230758 140029 230818 140286
rect 230755 140028 230821 140029
rect 230755 139964 230756 140028
rect 230820 139964 230821 140028
rect 230755 139963 230821 139964
rect 198555 135132 198621 135133
rect 198555 135068 198556 135132
rect 198620 135068 198621 135132
rect 198555 135067 198621 135068
rect 198558 132549 198618 135067
rect 178683 132548 178749 132549
rect 178683 132484 178684 132548
rect 178748 132484 178749 132548
rect 178683 132483 178749 132484
rect 182915 132548 182981 132549
rect 182915 132484 182916 132548
rect 182980 132484 182981 132548
rect 182915 132483 182981 132484
rect 198555 132548 198621 132549
rect 198555 132484 198556 132548
rect 198620 132484 198621 132548
rect 198555 132483 198621 132484
rect 199291 132548 199357 132549
rect 199291 132484 199292 132548
rect 199356 132484 199357 132548
rect 199291 132483 199357 132484
rect 178686 124882 178746 132483
rect 199294 131002 199354 132483
rect 241982 129557 242042 141731
rect 242534 139757 242594 142411
rect 261670 142205 261730 180763
rect 262403 180692 262469 180693
rect 262403 180628 262404 180692
rect 262468 180628 262469 180692
rect 262403 180627 262469 180628
rect 261667 142204 261733 142205
rect 261667 142140 261668 142204
rect 261732 142140 261733 142204
rect 261667 142139 261733 142140
rect 262406 141202 262466 180627
rect 262955 180556 263021 180557
rect 262955 180492 262956 180556
rect 263020 180492 263021 180556
rect 262955 180491 263021 180492
rect 262958 143242 263018 180491
rect 271422 179962 271482 181987
rect 287427 179332 287493 179333
rect 287427 179282 287428 179332
rect 287492 179282 287493 179332
rect 289451 179332 289517 179333
rect 289451 179282 289452 179332
rect 289516 179282 289517 179332
rect 310979 179332 311045 179333
rect 310979 179282 310980 179332
rect 311044 179282 311045 179332
rect 317051 179332 317117 179333
rect 317051 179282 317052 179332
rect 317116 179282 317117 179332
rect 351646 172669 351706 184027
rect 351830 172669 351890 191374
rect 352747 191372 352748 191374
rect 352812 191372 352813 191436
rect 352747 191371 352813 191372
rect 435740 177298 439740 207698
rect 435740 177062 435862 177298
rect 436098 177062 436182 177298
rect 436418 177062 436502 177298
rect 436738 177062 436822 177298
rect 437058 177062 437142 177298
rect 437378 177062 437462 177298
rect 437698 177062 437782 177298
rect 438018 177062 438102 177298
rect 438338 177062 438422 177298
rect 438658 177062 438742 177298
rect 438978 177062 439062 177298
rect 439298 177062 439382 177298
rect 439618 177062 439740 177298
rect 351643 172668 351709 172669
rect 351643 172604 351644 172668
rect 351708 172604 351709 172668
rect 351643 172603 351709 172604
rect 351827 172668 351893 172669
rect 351827 172604 351828 172668
rect 351892 172604 351893 172668
rect 351827 172603 351893 172604
rect 435740 146662 439740 177062
rect 435740 146426 435862 146662
rect 436098 146426 436182 146662
rect 436418 146426 436502 146662
rect 436738 146426 436822 146662
rect 437058 146426 437142 146662
rect 437378 146426 437462 146662
rect 437698 146426 437782 146662
rect 438018 146426 438102 146662
rect 438338 146426 438422 146662
rect 438658 146426 438742 146662
rect 438978 146426 439062 146662
rect 439298 146426 439382 146662
rect 439618 146426 439740 146662
rect 290003 144516 290069 144517
rect 290003 144452 290004 144516
rect 290068 144452 290069 144516
rect 290003 144451 290069 144452
rect 243086 139893 243146 140286
rect 243083 139892 243149 139893
rect 243083 139828 243084 139892
rect 243148 139828 243149 139892
rect 243083 139827 243149 139828
rect 251366 139757 251426 140286
rect 262958 139893 263018 143006
rect 290006 141882 290066 144451
rect 262955 139892 263021 139893
rect 262955 139828 262956 139892
rect 263020 139828 263021 139892
rect 262955 139827 263021 139828
rect 242531 139756 242597 139757
rect 242531 139692 242532 139756
rect 242596 139692 242597 139756
rect 242531 139691 242597 139692
rect 251363 139756 251429 139757
rect 251363 139692 251364 139756
rect 251428 139692 251429 139756
rect 251363 139691 251429 139692
rect 351643 139620 351709 139621
rect 351643 139556 351644 139620
rect 351708 139556 351709 139620
rect 351643 139555 351709 139556
rect 351827 139620 351893 139621
rect 351827 139556 351828 139620
rect 351892 139556 351893 139620
rect 351827 139555 351893 139556
rect 252651 138532 252717 138533
rect 252651 138468 252652 138532
rect 252716 138468 252717 138532
rect 252651 138467 252717 138468
rect 249707 138396 249773 138397
rect 249707 138332 249708 138396
rect 249772 138332 249773 138396
rect 249707 138331 249773 138332
rect 249155 134452 249221 134453
rect 249155 134388 249156 134452
rect 249220 134388 249221 134452
rect 249155 134387 249221 134388
rect 246211 130236 246277 130237
rect 246211 130172 246212 130236
rect 246276 130172 246277 130236
rect 246211 130171 246277 130172
rect 241979 129556 242045 129557
rect 241979 129492 241980 129556
rect 242044 129492 242045 129556
rect 241979 129491 242045 129492
rect 242163 124796 242229 124797
rect 242163 124732 242164 124796
rect 242228 124732 242229 124796
rect 242163 124731 242229 124732
rect 148691 122348 148757 122349
rect 148691 122284 148692 122348
rect 148756 122284 148757 122348
rect 148691 122283 148757 122284
rect 148694 122074 148754 122283
rect 148875 122212 148941 122213
rect 148875 122148 148876 122212
rect 148940 122148 148941 122212
rect 148875 122147 148941 122148
rect 148878 122074 148938 122147
rect 148694 122014 148938 122074
rect 163782 115362 163842 117846
rect 147771 113236 147837 113237
rect 147771 113172 147772 113236
rect 147836 113172 147837 113236
rect 147771 113171 147837 113172
rect 74539 112828 74605 112829
rect 74539 112764 74540 112828
rect 74604 112764 74605 112828
rect 74539 112763 74605 112764
rect 148694 109094 148938 109154
rect 148694 108885 148754 109094
rect 148878 108885 148938 109094
rect 148691 108884 148757 108885
rect 148691 108820 148692 108884
rect 148756 108820 148757 108884
rect 148691 108819 148757 108820
rect 148875 108884 148941 108885
rect 148875 108820 148876 108884
rect 148940 108820 148941 108884
rect 148875 108819 148941 108820
rect 137467 106844 137533 106845
rect 137467 106780 137468 106844
rect 137532 106780 137533 106844
rect 137467 106779 137533 106780
rect 74171 102084 74237 102085
rect 74171 102020 74172 102084
rect 74236 102020 74237 102084
rect 74171 102019 74237 102020
rect 137470 101762 137530 106779
rect 104464 100708 104784 100750
rect 104464 100472 104506 100708
rect 104742 100472 104784 100708
rect 104464 100430 104784 100472
rect 145747 99908 145813 99909
rect 145747 99844 145748 99908
rect 145812 99844 145813 99908
rect 145747 99843 145813 99844
rect 145750 99722 145810 99843
rect 73619 98276 73685 98277
rect 73619 98212 73620 98276
rect 73684 98212 73685 98276
rect 73619 98211 73685 98212
rect 148875 95556 148941 95557
rect 148875 95492 148876 95556
rect 148940 95492 148941 95556
rect 148875 95491 148941 95492
rect 74539 93924 74605 93925
rect 74539 93860 74540 93924
rect 74604 93860 74605 93924
rect 74539 93859 74605 93860
rect 74542 93602 74602 93859
rect 148878 90117 148938 95491
rect 152190 90117 152250 113766
rect 163782 105842 163842 114446
rect 178686 108562 178746 123966
rect 242166 119442 242226 124731
rect 242314 119294 242594 119354
rect 229286 116637 229346 117846
rect 229283 116636 229349 116637
rect 229283 116572 229284 116636
rect 229348 116572 229349 116636
rect 229283 116571 229349 116572
rect 183104 116026 183424 116068
rect 183104 115790 183146 116026
rect 183382 115790 183424 116026
rect 183104 115748 183424 115790
rect 230755 112964 230821 112965
rect 230755 112900 230756 112964
rect 230820 112900 230821 112964
rect 230755 112899 230821 112900
rect 230758 112642 230818 112899
rect 242534 110245 242594 119294
rect 245478 116722 245538 123286
rect 241979 110244 242045 110245
rect 241979 110180 241980 110244
rect 242044 110180 242045 110244
rect 241979 110179 242045 110180
rect 242531 110244 242597 110245
rect 242531 110180 242532 110244
rect 242596 110180 242597 110244
rect 242531 110179 242597 110180
rect 230755 107932 230821 107933
rect 230755 107868 230756 107932
rect 230820 107868 230821 107932
rect 230755 107867 230821 107868
rect 163782 94282 163842 104926
rect 164886 100725 164946 104246
rect 177030 102357 177090 102886
rect 171323 102356 171389 102357
rect 171323 102292 171324 102356
rect 171388 102292 171389 102356
rect 171323 102291 171389 102292
rect 177027 102356 177093 102357
rect 177027 102292 177028 102356
rect 177092 102292 177093 102356
rect 177027 102291 177093 102292
rect 171326 101762 171386 102291
rect 164883 100724 164949 100725
rect 164883 100660 164884 100724
rect 164948 100660 164949 100724
rect 164883 100659 164949 100660
rect 164883 98684 164949 98685
rect 164883 98620 164884 98684
rect 164948 98620 164949 98684
rect 164883 98619 164949 98620
rect 164886 98362 164946 98619
rect 177950 96322 178010 106966
rect 228731 103988 228797 103989
rect 228731 103924 228732 103988
rect 228796 103924 228797 103988
rect 228731 103923 228797 103924
rect 178686 100725 178746 103566
rect 228734 102354 228794 103923
rect 228734 102294 229014 102354
rect 230758 101762 230818 107867
rect 178683 100724 178749 100725
rect 178683 100660 178684 100724
rect 178748 100660 178749 100724
rect 178683 100659 178749 100660
rect 198464 100708 198784 100750
rect 241982 100725 242042 110179
rect 245478 105162 245538 116486
rect 245846 114002 245906 123966
rect 198464 100472 198506 100708
rect 198742 100472 198784 100708
rect 241979 100724 242045 100725
rect 241979 100660 241980 100724
rect 242044 100660 242045 100724
rect 241979 100659 242045 100660
rect 198464 100430 198784 100472
rect 178683 100044 178749 100045
rect 178683 99980 178684 100044
rect 178748 99980 178749 100044
rect 178683 99979 178749 99980
rect 228731 100044 228797 100045
rect 228731 99980 228732 100044
rect 228796 99980 228797 100044
rect 228731 99979 228797 99980
rect 178686 99042 178746 99979
rect 228734 98362 228794 99979
rect 242715 99908 242781 99909
rect 242715 99844 242716 99908
rect 242780 99844 242781 99908
rect 242715 99843 242781 99844
rect 242718 99722 242778 99843
rect 245478 96322 245538 103566
rect 241979 95828 242045 95829
rect 241979 95764 241980 95828
rect 242044 95764 242045 95828
rect 241979 95763 242045 95764
rect 155466 90734 155746 90794
rect 148875 90116 148941 90117
rect 148875 90052 148876 90116
rect 148940 90052 148941 90116
rect 148875 90051 148941 90052
rect 152187 90116 152253 90117
rect 152187 90052 152188 90116
rect 152252 90052 152253 90116
rect 152187 90051 152253 90052
rect 155499 90116 155565 90117
rect 155499 90052 155500 90116
rect 155564 90052 155565 90116
rect 155499 90051 155565 90052
rect 74171 89844 74237 89845
rect 74171 89780 74172 89844
rect 74236 89780 74237 89844
rect 74171 89779 74237 89780
rect 74174 87533 74234 89779
rect 155502 88893 155562 90051
rect 155686 88893 155746 90734
rect 241982 89029 242042 95763
rect 245846 89165 245906 113766
rect 245843 89164 245909 89165
rect 245843 89100 245844 89164
rect 245908 89100 245909 89164
rect 245843 89099 245909 89100
rect 241979 89028 242045 89029
rect 241979 88964 241980 89028
rect 242044 88964 242045 89028
rect 241979 88963 242045 88964
rect 155499 88892 155565 88893
rect 155499 88828 155500 88892
rect 155564 88828 155565 88892
rect 155499 88827 155565 88828
rect 155683 88892 155749 88893
rect 155683 88828 155684 88892
rect 155748 88828 155749 88892
rect 241979 88892 242045 88893
rect 155683 88827 155749 88828
rect 241979 88828 241980 88892
rect 242044 88828 242045 88892
rect 241979 88827 242045 88828
rect 74171 87532 74237 87533
rect 74171 87468 74172 87532
rect 74236 87468 74237 87532
rect 74171 87467 74237 87468
rect 72883 86308 72949 86309
rect 72883 86244 72884 86308
rect 72948 86244 72949 86308
rect 72883 86243 72949 86244
rect 72699 86172 72765 86173
rect 72699 86108 72700 86172
rect 72764 86108 72765 86172
rect 72699 86107 72765 86108
rect 52643 77876 52709 77877
rect 52643 77812 52644 77876
rect 52708 77812 52709 77876
rect 52643 77811 52709 77812
rect 54667 77876 54733 77877
rect 54667 77812 54668 77876
rect 54732 77812 54733 77876
rect 54667 77811 54733 77812
rect 55403 77876 55469 77877
rect 55403 77812 55404 77876
rect 55468 77812 55469 77876
rect 55403 77811 55469 77812
rect 72702 73794 72762 86107
rect 72886 75154 72946 86243
rect 73987 86172 74053 86173
rect 73987 86108 73988 86172
rect 74052 86108 74053 86172
rect 73987 86107 74053 86108
rect 72886 75094 73866 75154
rect 72702 73734 73498 73794
rect 5000 54518 5122 54754
rect 5358 54518 5442 54754
rect 5678 54518 5762 54754
rect 5998 54518 6082 54754
rect 6318 54518 6402 54754
rect 6638 54518 6722 54754
rect 6958 54518 7042 54754
rect 7278 54518 7362 54754
rect 7598 54518 7682 54754
rect 7918 54518 8002 54754
rect 8238 54518 8322 54754
rect 8558 54518 8642 54754
rect 8878 54518 9000 54754
rect 5000 24118 9000 54518
rect 73438 49314 73498 73734
rect 72886 49254 73498 49314
rect 67918 48093 67978 48486
rect 67915 48092 67981 48093
rect 67915 48028 67916 48092
rect 67980 48028 67981 48092
rect 67915 48027 67981 48028
rect 72886 47413 72946 49254
rect 73806 48634 73866 75094
rect 73402 48574 73866 48634
rect 73990 48093 74050 86107
rect 73987 48092 74053 48093
rect 73987 48028 73988 48092
rect 74052 48028 74053 48092
rect 73987 48027 74053 48028
rect 72883 47412 72949 47413
rect 72883 47348 72884 47412
rect 72948 47348 72949 47412
rect 72883 47347 72949 47348
rect 74174 46189 74234 87467
rect 156051 87396 156117 87397
rect 156051 87332 156052 87396
rect 156116 87332 156117 87396
rect 156051 87331 156117 87332
rect 167643 87396 167709 87397
rect 167643 87332 167644 87396
rect 167708 87332 167709 87396
rect 167643 87331 167709 87332
rect 148507 87260 148573 87261
rect 148507 87196 148508 87260
rect 148572 87196 148573 87260
rect 148507 87195 148573 87196
rect 74539 86444 74605 86445
rect 74539 86380 74540 86444
rect 74604 86380 74605 86444
rect 74539 86379 74605 86380
rect 74542 49402 74602 86379
rect 148510 73882 148570 87195
rect 156054 73882 156114 87331
rect 144646 64362 144706 72966
rect 113915 53124 113981 53125
rect 113915 53060 113916 53124
rect 113980 53060 113981 53124
rect 113915 53059 113981 53060
rect 118699 53124 118765 53125
rect 118699 53060 118700 53124
rect 118764 53060 118765 53124
rect 118699 53059 118765 53060
rect 107475 50268 107541 50269
rect 107475 50204 107476 50268
rect 107540 50204 107541 50268
rect 107475 50203 107541 50204
rect 109315 50268 109381 50269
rect 109315 50204 109316 50268
rect 109380 50204 109381 50268
rect 109315 50203 109381 50204
rect 74171 46188 74237 46189
rect 74171 46124 74172 46188
rect 74236 46124 74237 46188
rect 74171 46123 74237 46124
rect 74542 45917 74602 49166
rect 107478 47413 107538 50203
rect 107475 47412 107541 47413
rect 107475 47348 107476 47412
rect 107540 47348 107541 47412
rect 107475 47347 107541 47348
rect 107478 46682 107538 47347
rect 109318 47277 109378 50203
rect 109315 47276 109381 47277
rect 109315 47212 109316 47276
rect 109380 47212 109381 47276
rect 109315 47211 109381 47212
rect 74539 45916 74605 45917
rect 74539 45852 74540 45916
rect 74604 45852 74605 45916
rect 74539 45851 74605 45852
rect 113918 43333 113978 53059
rect 118702 46189 118762 53059
rect 142438 51085 142498 51206
rect 142435 51084 142501 51085
rect 142435 51020 142436 51084
rect 142500 51020 142501 51084
rect 142435 51019 142501 51020
rect 144830 49314 144890 63446
rect 144830 49254 145478 49314
rect 145566 47957 145626 49166
rect 147958 48093 148018 49166
rect 167646 48722 167706 87331
rect 168747 87124 168813 87125
rect 168747 87060 168748 87124
rect 168812 87060 168813 87124
rect 168747 87059 168813 87060
rect 168011 86852 168077 86853
rect 168011 86788 168012 86852
rect 168076 86788 168077 86852
rect 168011 86787 168077 86788
rect 168014 49402 168074 86787
rect 154766 48093 154826 48486
rect 147955 48092 148021 48093
rect 147955 48028 147956 48092
rect 148020 48028 148021 48092
rect 147955 48027 148021 48028
rect 154763 48092 154829 48093
rect 154763 48028 154764 48092
rect 154828 48028 154829 48092
rect 154763 48027 154829 48028
rect 145563 47956 145629 47957
rect 145563 47892 145564 47956
rect 145628 47892 145629 47956
rect 145563 47891 145629 47892
rect 147955 47956 148021 47957
rect 147955 47892 147956 47956
rect 148020 47892 148021 47956
rect 147955 47891 148021 47892
rect 118699 46188 118765 46189
rect 118699 46124 118700 46188
rect 118764 46124 118765 46188
rect 118699 46123 118765 46124
rect 147958 45781 148018 47891
rect 168014 47549 168074 49166
rect 168750 47957 168810 87059
rect 169299 86988 169365 86989
rect 169299 86924 169300 86988
rect 169364 86924 169365 86988
rect 169299 86923 169365 86924
rect 169115 86716 169181 86717
rect 169115 86652 169116 86716
rect 169180 86652 169181 86716
rect 169115 86651 169181 86652
rect 169118 48042 169178 86651
rect 169302 48634 169362 86923
rect 178686 84269 178746 88606
rect 241982 86714 242042 88827
rect 246214 87533 246274 130171
rect 249158 127602 249218 134387
rect 249710 126837 249770 138331
rect 252654 137853 252714 138467
rect 252651 137852 252717 137853
rect 252651 137788 252652 137852
rect 252716 137788 252717 137852
rect 252651 137787 252717 137788
rect 298099 137852 298165 137853
rect 298099 137788 298100 137852
rect 298164 137788 298165 137852
rect 298099 137787 298165 137788
rect 252654 127517 252714 137787
rect 298102 132549 298162 137787
rect 298099 132548 298165 132549
rect 298099 132484 298100 132548
rect 298164 132484 298165 132548
rect 298099 132483 298165 132484
rect 252651 127516 252717 127517
rect 252651 127452 252652 127516
rect 252716 127452 252717 127516
rect 252651 127451 252717 127452
rect 259643 127516 259709 127517
rect 259643 127452 259644 127516
rect 259708 127452 259709 127516
rect 259643 127451 259709 127452
rect 249707 126836 249773 126837
rect 249707 126772 249708 126836
rect 249772 126772 249773 126836
rect 249707 126771 249773 126772
rect 258726 100725 258786 103566
rect 258723 100724 258789 100725
rect 258723 100660 258724 100724
rect 258788 100660 258789 100724
rect 258723 100659 258789 100660
rect 258723 100044 258789 100045
rect 258723 99980 258724 100044
rect 258788 99980 258789 100044
rect 258723 99979 258789 99980
rect 258726 99722 258786 99979
rect 249526 88893 249586 89966
rect 249523 88892 249589 88893
rect 249523 88842 249524 88892
rect 249588 88842 249589 88892
rect 251731 88620 251797 88621
rect 251731 88556 251732 88620
rect 251796 88556 251797 88620
rect 251731 88555 251797 88556
rect 251734 88162 251794 88555
rect 259646 88162 259706 127451
rect 277104 116026 277424 116068
rect 277104 115790 277146 116026
rect 277382 115790 277424 116026
rect 277104 115748 277424 115790
rect 324595 106844 324661 106845
rect 324595 106780 324596 106844
rect 324660 106780 324661 106844
rect 324595 106779 324661 106780
rect 322755 103988 322821 103989
rect 322755 103924 322756 103988
rect 322820 103924 322821 103988
rect 322755 103923 322821 103924
rect 270499 103036 270565 103037
rect 270499 102972 270500 103036
rect 270564 102972 270565 103036
rect 270499 102971 270565 102972
rect 270502 101762 270562 102971
rect 322758 102354 322818 103923
rect 322758 102294 323038 102354
rect 272710 100725 272770 102206
rect 324598 101762 324658 106779
rect 272707 100724 272773 100725
rect 272707 100660 272708 100724
rect 272772 100660 272773 100724
rect 272707 100659 272773 100660
rect 292464 100708 292784 100750
rect 292464 100472 292506 100708
rect 292742 100472 292784 100708
rect 292464 100430 292784 100472
rect 322755 100452 322821 100453
rect 322755 100388 322756 100452
rect 322820 100388 322821 100452
rect 322755 100387 322821 100388
rect 272707 100044 272773 100045
rect 272707 99980 272708 100044
rect 272772 99980 272773 100044
rect 272707 99979 272773 99980
rect 272710 99722 272770 99979
rect 322758 98362 322818 100387
rect 351646 90117 351706 139555
rect 351830 134317 351890 139555
rect 351827 134316 351893 134317
rect 351827 134252 351828 134316
rect 351892 134252 351893 134316
rect 351827 134251 351893 134252
rect 352563 134180 352629 134181
rect 352563 134116 352564 134180
rect 352628 134116 352629 134180
rect 352563 134115 352629 134116
rect 352566 124794 352626 134115
rect 352198 124734 352626 124794
rect 352198 117314 352258 124734
rect 351830 117254 352258 117314
rect 351830 108474 351890 117254
rect 435740 116026 439740 146426
rect 435740 115790 435862 116026
rect 436098 115790 436182 116026
rect 436418 115790 436502 116026
rect 436738 115790 436822 116026
rect 437058 115790 437142 116026
rect 437378 115790 437462 116026
rect 437698 115790 437782 116026
rect 438018 115790 438102 116026
rect 438338 115790 438422 116026
rect 438658 115790 438742 116026
rect 438978 115790 439062 116026
rect 439298 115790 439382 116026
rect 439618 115790 439740 116026
rect 351830 108414 352810 108474
rect 352750 97869 352810 108414
rect 352747 97868 352813 97869
rect 352747 97804 352748 97868
rect 352812 97804 352813 97868
rect 352747 97803 352813 97804
rect 352750 97594 352810 97803
rect 352014 97534 352810 97594
rect 351643 90116 351709 90117
rect 351643 90052 351644 90116
rect 351708 90052 351709 90116
rect 351643 90051 351709 90052
rect 246211 87532 246277 87533
rect 246211 87468 246212 87532
rect 246276 87468 246277 87532
rect 246211 87467 246277 87468
rect 251179 87396 251245 87397
rect 251179 87332 251180 87396
rect 251244 87332 251245 87396
rect 251179 87331 251245 87332
rect 241982 86654 242226 86714
rect 178683 84268 178749 84269
rect 178683 84204 178684 84268
rect 178748 84204 178749 84268
rect 178683 84203 178749 84204
rect 242166 83453 242226 86654
rect 251182 86309 251242 87331
rect 251179 86308 251245 86309
rect 251179 86244 251180 86308
rect 251244 86244 251245 86308
rect 251179 86243 251245 86244
rect 249891 86172 249957 86173
rect 249891 86108 249892 86172
rect 249956 86108 249957 86172
rect 249891 86107 249957 86108
rect 242163 83452 242229 83453
rect 242163 83388 242164 83452
rect 242228 83388 242229 83452
rect 242163 83387 242229 83388
rect 242899 83452 242965 83453
rect 242899 83388 242900 83452
rect 242964 83388 242965 83452
rect 242899 83387 242965 83388
rect 242902 75429 242962 83387
rect 238667 75428 238733 75429
rect 238667 75364 238668 75428
rect 238732 75364 238733 75428
rect 238667 75363 238733 75364
rect 242899 75428 242965 75429
rect 242899 75364 242900 75428
rect 242964 75364 242965 75428
rect 242899 75363 242965 75364
rect 170038 52714 170098 73646
rect 238670 60282 238730 75363
rect 249894 73882 249954 86107
rect 251182 75429 251242 86243
rect 251179 75428 251245 75429
rect 251179 75364 251180 75428
rect 251244 75364 251245 75428
rect 251179 75363 251245 75364
rect 237382 54074 237442 59366
rect 237382 54014 237810 54074
rect 212539 53124 212605 53125
rect 212539 53060 212540 53124
rect 212604 53060 212605 53124
rect 212539 53059 212605 53060
rect 170038 52654 170466 52714
rect 170406 50674 170466 52654
rect 191379 51628 191445 51629
rect 191379 51564 191380 51628
rect 191444 51564 191445 51628
rect 191379 51563 191445 51564
rect 204259 51628 204325 51629
rect 204259 51564 204260 51628
rect 204324 51564 204325 51628
rect 204259 51563 204325 51564
rect 170587 50676 170653 50677
rect 170587 50674 170588 50676
rect 170406 50614 170588 50674
rect 170587 50612 170588 50614
rect 170652 50612 170653 50676
rect 170587 50611 170653 50612
rect 191382 48722 191442 51563
rect 169302 48574 169730 48634
rect 168747 47956 168813 47957
rect 168747 47892 168748 47956
rect 168812 47892 168813 47956
rect 168747 47891 168813 47892
rect 168011 47548 168077 47549
rect 168011 47484 168012 47548
rect 168076 47484 168077 47548
rect 168011 47483 168077 47484
rect 157526 45917 157586 46446
rect 158998 46053 159058 47126
rect 169670 46053 169730 48574
rect 181811 46732 181877 46733
rect 181811 46682 181812 46732
rect 181876 46682 181877 46732
rect 204262 46682 204322 51563
rect 207755 51356 207821 51357
rect 207755 51292 207756 51356
rect 207820 51292 207821 51356
rect 207755 51291 207821 51292
rect 158995 46052 159061 46053
rect 158995 45988 158996 46052
rect 159060 45988 159061 46052
rect 158995 45987 159061 45988
rect 169667 46052 169733 46053
rect 169667 45988 169668 46052
rect 169732 45988 169733 46052
rect 169667 45987 169733 45988
rect 157523 45916 157589 45917
rect 157523 45852 157524 45916
rect 157588 45852 157589 45916
rect 157523 45851 157589 45852
rect 147955 45780 148021 45781
rect 147955 45716 147956 45780
rect 148020 45716 148021 45780
rect 147955 45715 148021 45716
rect 204262 45373 204322 46446
rect 204259 45372 204325 45373
rect 204259 45308 204260 45372
rect 204324 45308 204325 45372
rect 204259 45307 204325 45308
rect 113915 43332 113981 43333
rect 113915 43268 113916 43332
rect 113980 43268 113981 43332
rect 113915 43267 113981 43268
rect 207758 37757 207818 51291
rect 212542 47413 212602 53059
rect 237750 50762 237810 54014
rect 238670 48093 238730 51206
rect 238667 48092 238733 48093
rect 238667 48028 238668 48092
rect 238732 48028 238733 48092
rect 238667 48027 238733 48028
rect 212539 47412 212605 47413
rect 212539 47348 212540 47412
rect 212604 47348 212605 47412
rect 212539 47347 212605 47348
rect 248974 46053 249034 48486
rect 261670 47957 261730 87926
rect 262403 86852 262469 86853
rect 262403 86788 262404 86852
rect 262468 86788 262469 86852
rect 262403 86787 262469 86788
rect 261851 75428 261917 75429
rect 261851 75364 261852 75428
rect 261916 75364 261917 75428
rect 261851 75363 261917 75364
rect 261854 48093 261914 75363
rect 262406 48093 262466 86787
rect 262587 86716 262653 86717
rect 262587 86652 262588 86716
rect 262652 86652 262653 86716
rect 262587 86651 262653 86652
rect 261851 48092 261917 48093
rect 261851 48028 261852 48092
rect 261916 48028 261917 48092
rect 261851 48027 261917 48028
rect 262403 48092 262469 48093
rect 262403 48028 262404 48092
rect 262468 48028 262469 48092
rect 262403 48027 262469 48028
rect 261667 47956 261733 47957
rect 261667 47892 261668 47956
rect 261732 47892 261733 47956
rect 261667 47891 261733 47892
rect 261854 46682 261914 48027
rect 248971 46052 249037 46053
rect 248971 45988 248972 46052
rect 249036 45988 249037 46052
rect 248971 45987 249037 45988
rect 252838 45917 252898 46446
rect 262590 46053 262650 86651
rect 263878 49314 263938 88606
rect 336371 86716 336437 86717
rect 336371 86652 336372 86716
rect 336436 86652 336437 86716
rect 336371 86651 336437 86652
rect 263510 49254 263938 49314
rect 263510 47954 263570 49254
rect 264246 48722 264306 73646
rect 301595 53124 301661 53125
rect 301595 53060 301596 53124
rect 301660 53060 301661 53124
rect 301595 53059 301661 53060
rect 306563 53124 306629 53125
rect 306563 53060 306564 53124
rect 306628 53060 306629 53124
rect 306563 53059 306629 53060
rect 270686 51357 270746 51886
rect 270683 51356 270749 51357
rect 270683 51292 270684 51356
rect 270748 51292 270749 51356
rect 270683 51291 270749 51292
rect 264246 48093 264306 48486
rect 264243 48092 264309 48093
rect 264243 48028 264244 48092
rect 264308 48028 264309 48092
rect 264243 48027 264309 48028
rect 263510 47894 263938 47954
rect 263878 47413 263938 47894
rect 263875 47412 263941 47413
rect 263875 47362 263876 47412
rect 263940 47362 263941 47412
rect 262587 46052 262653 46053
rect 262587 45988 262588 46052
rect 262652 45988 262653 46052
rect 262587 45987 262653 45988
rect 252835 45916 252901 45917
rect 252835 45852 252836 45916
rect 252900 45852 252901 45916
rect 252835 45851 252901 45852
rect 301598 37757 301658 53059
rect 306566 47413 306626 53059
rect 306563 47412 306629 47413
rect 306563 47348 306564 47412
rect 306628 47348 306629 47412
rect 306563 47347 306629 47348
rect 336374 46053 336434 86651
rect 351646 77877 351706 90051
rect 352014 79234 352074 97534
rect 351830 79174 352074 79234
rect 435740 85390 439740 115790
rect 435740 85154 435862 85390
rect 436098 85154 436182 85390
rect 436418 85154 436502 85390
rect 436738 85154 436822 85390
rect 437058 85154 437142 85390
rect 437378 85154 437462 85390
rect 437698 85154 437782 85390
rect 438018 85154 438102 85390
rect 438338 85154 438422 85390
rect 438658 85154 438742 85390
rect 438978 85154 439062 85390
rect 439298 85154 439382 85390
rect 439618 85154 439740 85390
rect 351830 77877 351890 79174
rect 351643 77876 351709 77877
rect 351643 77812 351644 77876
rect 351708 77812 351709 77876
rect 351643 77811 351709 77812
rect 351827 77876 351893 77877
rect 351827 77812 351828 77876
rect 351892 77812 351893 77876
rect 351827 77811 351893 77812
rect 435740 54754 439740 85154
rect 435740 54518 435862 54754
rect 436098 54518 436182 54754
rect 436418 54518 436502 54754
rect 436738 54518 436822 54754
rect 437058 54518 437142 54754
rect 437378 54518 437462 54754
rect 437698 54518 437782 54754
rect 438018 54518 438102 54754
rect 438338 54518 438422 54754
rect 438658 54518 438742 54754
rect 438978 54518 439062 54754
rect 439298 54518 439382 54754
rect 439618 54518 439740 54754
rect 358451 50404 358517 50405
rect 358451 50340 358452 50404
rect 358516 50340 358517 50404
rect 358451 50339 358517 50340
rect 358454 47549 358514 50339
rect 358451 47548 358517 47549
rect 358451 47484 358452 47548
rect 358516 47484 358517 47548
rect 358451 47483 358517 47484
rect 336371 46052 336437 46053
rect 336371 45988 336372 46052
rect 336436 45988 336437 46052
rect 336371 45987 336437 45988
rect 207755 37756 207821 37757
rect 207755 37692 207756 37756
rect 207820 37692 207821 37756
rect 207755 37691 207821 37692
rect 301595 37756 301661 37757
rect 301595 37692 301596 37756
rect 301660 37692 301661 37756
rect 301595 37691 301661 37692
rect 5000 23882 5122 24118
rect 5358 23882 5442 24118
rect 5678 23882 5762 24118
rect 5998 23882 6082 24118
rect 6318 23882 6402 24118
rect 6638 23882 6722 24118
rect 6958 23882 7042 24118
rect 7278 23882 7362 24118
rect 7598 23882 7682 24118
rect 7918 23882 8002 24118
rect 8238 23882 8322 24118
rect 8558 23882 8642 24118
rect 8878 23882 9000 24118
rect 5000 8878 9000 23882
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 9000 8878
rect 5000 8558 9000 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 9000 8558
rect 5000 8238 9000 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 9000 8238
rect 5000 7918 9000 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 9000 7918
rect 5000 7598 9000 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 9000 7598
rect 5000 7278 9000 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 9000 7278
rect 5000 6958 9000 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 9000 6958
rect 5000 6638 9000 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 9000 6638
rect 5000 6318 9000 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 9000 6318
rect 5000 5998 9000 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 9000 5998
rect 5000 5678 9000 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 9000 5678
rect 5000 5358 9000 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 9000 5358
rect 5000 5000 9000 5122
rect 435740 24118 439740 54518
rect 435740 23882 435862 24118
rect 436098 23882 436182 24118
rect 436418 23882 436502 24118
rect 436738 23882 436822 24118
rect 437058 23882 437142 24118
rect 437378 23882 437462 24118
rect 437698 23882 437782 24118
rect 438018 23882 438102 24118
rect 438338 23882 438422 24118
rect 438658 23882 438742 24118
rect 438978 23882 439062 24118
rect 439298 23882 439382 24118
rect 439618 23882 439740 24118
rect 435740 8878 439740 23882
rect 435740 8642 435862 8878
rect 436098 8642 436182 8878
rect 436418 8642 436502 8878
rect 436738 8642 436822 8878
rect 437058 8642 437142 8878
rect 437378 8642 437462 8878
rect 437698 8642 437782 8878
rect 438018 8642 438102 8878
rect 438338 8642 438422 8878
rect 438658 8642 438742 8878
rect 438978 8642 439062 8878
rect 439298 8642 439382 8878
rect 439618 8642 439740 8878
rect 435740 8558 439740 8642
rect 435740 8322 435862 8558
rect 436098 8322 436182 8558
rect 436418 8322 436502 8558
rect 436738 8322 436822 8558
rect 437058 8322 437142 8558
rect 437378 8322 437462 8558
rect 437698 8322 437782 8558
rect 438018 8322 438102 8558
rect 438338 8322 438422 8558
rect 438658 8322 438742 8558
rect 438978 8322 439062 8558
rect 439298 8322 439382 8558
rect 439618 8322 439740 8558
rect 435740 8238 439740 8322
rect 435740 8002 435862 8238
rect 436098 8002 436182 8238
rect 436418 8002 436502 8238
rect 436738 8002 436822 8238
rect 437058 8002 437142 8238
rect 437378 8002 437462 8238
rect 437698 8002 437782 8238
rect 438018 8002 438102 8238
rect 438338 8002 438422 8238
rect 438658 8002 438742 8238
rect 438978 8002 439062 8238
rect 439298 8002 439382 8238
rect 439618 8002 439740 8238
rect 435740 7918 439740 8002
rect 435740 7682 435862 7918
rect 436098 7682 436182 7918
rect 436418 7682 436502 7918
rect 436738 7682 436822 7918
rect 437058 7682 437142 7918
rect 437378 7682 437462 7918
rect 437698 7682 437782 7918
rect 438018 7682 438102 7918
rect 438338 7682 438422 7918
rect 438658 7682 438742 7918
rect 438978 7682 439062 7918
rect 439298 7682 439382 7918
rect 439618 7682 439740 7918
rect 435740 7598 439740 7682
rect 435740 7362 435862 7598
rect 436098 7362 436182 7598
rect 436418 7362 436502 7598
rect 436738 7362 436822 7598
rect 437058 7362 437142 7598
rect 437378 7362 437462 7598
rect 437698 7362 437782 7598
rect 438018 7362 438102 7598
rect 438338 7362 438422 7598
rect 438658 7362 438742 7598
rect 438978 7362 439062 7598
rect 439298 7362 439382 7598
rect 439618 7362 439740 7598
rect 435740 7278 439740 7362
rect 435740 7042 435862 7278
rect 436098 7042 436182 7278
rect 436418 7042 436502 7278
rect 436738 7042 436822 7278
rect 437058 7042 437142 7278
rect 437378 7042 437462 7278
rect 437698 7042 437782 7278
rect 438018 7042 438102 7278
rect 438338 7042 438422 7278
rect 438658 7042 438742 7278
rect 438978 7042 439062 7278
rect 439298 7042 439382 7278
rect 439618 7042 439740 7278
rect 435740 6958 439740 7042
rect 435740 6722 435862 6958
rect 436098 6722 436182 6958
rect 436418 6722 436502 6958
rect 436738 6722 436822 6958
rect 437058 6722 437142 6958
rect 437378 6722 437462 6958
rect 437698 6722 437782 6958
rect 438018 6722 438102 6958
rect 438338 6722 438422 6958
rect 438658 6722 438742 6958
rect 438978 6722 439062 6958
rect 439298 6722 439382 6958
rect 439618 6722 439740 6958
rect 435740 6638 439740 6722
rect 435740 6402 435862 6638
rect 436098 6402 436182 6638
rect 436418 6402 436502 6638
rect 436738 6402 436822 6638
rect 437058 6402 437142 6638
rect 437378 6402 437462 6638
rect 437698 6402 437782 6638
rect 438018 6402 438102 6638
rect 438338 6402 438422 6638
rect 438658 6402 438742 6638
rect 438978 6402 439062 6638
rect 439298 6402 439382 6638
rect 439618 6402 439740 6638
rect 435740 6318 439740 6402
rect 435740 6082 435862 6318
rect 436098 6082 436182 6318
rect 436418 6082 436502 6318
rect 436738 6082 436822 6318
rect 437058 6082 437142 6318
rect 437378 6082 437462 6318
rect 437698 6082 437782 6318
rect 438018 6082 438102 6318
rect 438338 6082 438422 6318
rect 438658 6082 438742 6318
rect 438978 6082 439062 6318
rect 439298 6082 439382 6318
rect 439618 6082 439740 6318
rect 435740 5998 439740 6082
rect 435740 5762 435862 5998
rect 436098 5762 436182 5998
rect 436418 5762 436502 5998
rect 436738 5762 436822 5998
rect 437058 5762 437142 5998
rect 437378 5762 437462 5998
rect 437698 5762 437782 5998
rect 438018 5762 438102 5998
rect 438338 5762 438422 5998
rect 438658 5762 438742 5998
rect 438978 5762 439062 5998
rect 439298 5762 439382 5998
rect 439618 5762 439740 5998
rect 435740 5678 439740 5762
rect 435740 5442 435862 5678
rect 436098 5442 436182 5678
rect 436418 5442 436502 5678
rect 436738 5442 436822 5678
rect 437058 5442 437142 5678
rect 437378 5442 437462 5678
rect 437698 5442 437782 5678
rect 438018 5442 438102 5678
rect 438338 5442 438422 5678
rect 438658 5442 438742 5678
rect 438978 5442 439062 5678
rect 439298 5442 439382 5678
rect 439618 5442 439740 5678
rect 435740 5358 439740 5442
rect 435740 5122 435862 5358
rect 436098 5122 436182 5358
rect 436418 5122 436502 5358
rect 436738 5122 436822 5358
rect 437058 5122 437142 5358
rect 437378 5122 437462 5358
rect 437698 5122 437782 5358
rect 438018 5122 438102 5358
rect 438338 5122 438422 5358
rect 438658 5122 438742 5358
rect 438978 5122 439062 5358
rect 439298 5122 439382 5358
rect 439618 5122 439740 5358
rect 435740 5000 439740 5122
rect 440740 376432 444740 401642
rect 440740 376196 440862 376432
rect 441098 376196 441182 376432
rect 441418 376196 441502 376432
rect 441738 376196 441822 376432
rect 442058 376196 442142 376432
rect 442378 376196 442462 376432
rect 442698 376196 442782 376432
rect 443018 376196 443102 376432
rect 443338 376196 443422 376432
rect 443658 376196 443742 376432
rect 443978 376196 444062 376432
rect 444298 376196 444382 376432
rect 444618 376196 444740 376432
rect 440740 345796 444740 376196
rect 440740 345560 440862 345796
rect 441098 345560 441182 345796
rect 441418 345560 441502 345796
rect 441738 345560 441822 345796
rect 442058 345560 442142 345796
rect 442378 345560 442462 345796
rect 442698 345560 442782 345796
rect 443018 345560 443102 345796
rect 443338 345560 443422 345796
rect 443658 345560 443742 345796
rect 443978 345560 444062 345796
rect 444298 345560 444382 345796
rect 444618 345560 444740 345796
rect 440740 315160 444740 345560
rect 440740 314924 440862 315160
rect 441098 314924 441182 315160
rect 441418 314924 441502 315160
rect 441738 314924 441822 315160
rect 442058 314924 442142 315160
rect 442378 314924 442462 315160
rect 442698 314924 442782 315160
rect 443018 314924 443102 315160
rect 443338 314924 443422 315160
rect 443658 314924 443742 315160
rect 443978 314924 444062 315160
rect 444298 314924 444382 315160
rect 444618 314924 444740 315160
rect 440740 284524 444740 314924
rect 440740 284288 440862 284524
rect 441098 284288 441182 284524
rect 441418 284288 441502 284524
rect 441738 284288 441822 284524
rect 442058 284288 442142 284524
rect 442378 284288 442462 284524
rect 442698 284288 442782 284524
rect 443018 284288 443102 284524
rect 443338 284288 443422 284524
rect 443658 284288 443742 284524
rect 443978 284288 444062 284524
rect 444298 284288 444382 284524
rect 444618 284288 444740 284524
rect 440740 253888 444740 284288
rect 440740 253652 440862 253888
rect 441098 253652 441182 253888
rect 441418 253652 441502 253888
rect 441738 253652 441822 253888
rect 442058 253652 442142 253888
rect 442378 253652 442462 253888
rect 442698 253652 442782 253888
rect 443018 253652 443102 253888
rect 443338 253652 443422 253888
rect 443658 253652 443742 253888
rect 443978 253652 444062 253888
rect 444298 253652 444382 253888
rect 444618 253652 444740 253888
rect 440740 223252 444740 253652
rect 440740 223016 440862 223252
rect 441098 223016 441182 223252
rect 441418 223016 441502 223252
rect 441738 223016 441822 223252
rect 442058 223016 442142 223252
rect 442378 223016 442462 223252
rect 442698 223016 442782 223252
rect 443018 223016 443102 223252
rect 443338 223016 443422 223252
rect 443658 223016 443742 223252
rect 443978 223016 444062 223252
rect 444298 223016 444382 223252
rect 444618 223016 444740 223252
rect 440740 192616 444740 223016
rect 440740 192380 440862 192616
rect 441098 192380 441182 192616
rect 441418 192380 441502 192616
rect 441738 192380 441822 192616
rect 442058 192380 442142 192616
rect 442378 192380 442462 192616
rect 442698 192380 442782 192616
rect 443018 192380 443102 192616
rect 443338 192380 443422 192616
rect 443658 192380 443742 192616
rect 443978 192380 444062 192616
rect 444298 192380 444382 192616
rect 444618 192380 444740 192616
rect 440740 161980 444740 192380
rect 440740 161744 440862 161980
rect 441098 161744 441182 161980
rect 441418 161744 441502 161980
rect 441738 161744 441822 161980
rect 442058 161744 442142 161980
rect 442378 161744 442462 161980
rect 442698 161744 442782 161980
rect 443018 161744 443102 161980
rect 443338 161744 443422 161980
rect 443658 161744 443742 161980
rect 443978 161744 444062 161980
rect 444298 161744 444382 161980
rect 444618 161744 444740 161980
rect 440740 131344 444740 161744
rect 440740 131108 440862 131344
rect 441098 131108 441182 131344
rect 441418 131108 441502 131344
rect 441738 131108 441822 131344
rect 442058 131108 442142 131344
rect 442378 131108 442462 131344
rect 442698 131108 442782 131344
rect 443018 131108 443102 131344
rect 443338 131108 443422 131344
rect 443658 131108 443742 131344
rect 443978 131108 444062 131344
rect 444298 131108 444382 131344
rect 444618 131108 444740 131344
rect 440740 100708 444740 131108
rect 440740 100472 440862 100708
rect 441098 100472 441182 100708
rect 441418 100472 441502 100708
rect 441738 100472 441822 100708
rect 442058 100472 442142 100708
rect 442378 100472 442462 100708
rect 442698 100472 442782 100708
rect 443018 100472 443102 100708
rect 443338 100472 443422 100708
rect 443658 100472 443742 100708
rect 443978 100472 444062 100708
rect 444298 100472 444382 100708
rect 444618 100472 444740 100708
rect 440740 70072 444740 100472
rect 440740 69836 440862 70072
rect 441098 69836 441182 70072
rect 441418 69836 441502 70072
rect 441738 69836 441822 70072
rect 442058 69836 442142 70072
rect 442378 69836 442462 70072
rect 442698 69836 442782 70072
rect 443018 69836 443102 70072
rect 443338 69836 443422 70072
rect 443658 69836 443742 70072
rect 443978 69836 444062 70072
rect 444298 69836 444382 70072
rect 444618 69836 444740 70072
rect 440740 39436 444740 69836
rect 440740 39200 440862 39436
rect 441098 39200 441182 39436
rect 441418 39200 441502 39436
rect 441738 39200 441822 39436
rect 442058 39200 442142 39436
rect 442378 39200 442462 39436
rect 442698 39200 442782 39436
rect 443018 39200 443102 39436
rect 443338 39200 443422 39436
rect 443658 39200 443742 39436
rect 443978 39200 444062 39436
rect 444298 39200 444382 39436
rect 444618 39200 444740 39436
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 4000 3878
rect 0 3558 4000 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 4000 3558
rect 0 3238 4000 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 4000 3238
rect 0 2918 4000 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 4000 2918
rect 0 2598 4000 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 4000 2598
rect 0 2278 4000 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 4000 2278
rect 0 1958 4000 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 4000 1958
rect 0 1638 4000 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 4000 1638
rect 0 1318 4000 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 4000 1318
rect 0 998 4000 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 4000 998
rect 0 678 4000 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 4000 678
rect 0 358 4000 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 4000 358
rect 0 0 4000 122
rect 440740 3878 444740 39200
rect 440740 3642 440862 3878
rect 441098 3642 441182 3878
rect 441418 3642 441502 3878
rect 441738 3642 441822 3878
rect 442058 3642 442142 3878
rect 442378 3642 442462 3878
rect 442698 3642 442782 3878
rect 443018 3642 443102 3878
rect 443338 3642 443422 3878
rect 443658 3642 443742 3878
rect 443978 3642 444062 3878
rect 444298 3642 444382 3878
rect 444618 3642 444740 3878
rect 440740 3558 444740 3642
rect 440740 3322 440862 3558
rect 441098 3322 441182 3558
rect 441418 3322 441502 3558
rect 441738 3322 441822 3558
rect 442058 3322 442142 3558
rect 442378 3322 442462 3558
rect 442698 3322 442782 3558
rect 443018 3322 443102 3558
rect 443338 3322 443422 3558
rect 443658 3322 443742 3558
rect 443978 3322 444062 3558
rect 444298 3322 444382 3558
rect 444618 3322 444740 3558
rect 440740 3238 444740 3322
rect 440740 3002 440862 3238
rect 441098 3002 441182 3238
rect 441418 3002 441502 3238
rect 441738 3002 441822 3238
rect 442058 3002 442142 3238
rect 442378 3002 442462 3238
rect 442698 3002 442782 3238
rect 443018 3002 443102 3238
rect 443338 3002 443422 3238
rect 443658 3002 443742 3238
rect 443978 3002 444062 3238
rect 444298 3002 444382 3238
rect 444618 3002 444740 3238
rect 440740 2918 444740 3002
rect 440740 2682 440862 2918
rect 441098 2682 441182 2918
rect 441418 2682 441502 2918
rect 441738 2682 441822 2918
rect 442058 2682 442142 2918
rect 442378 2682 442462 2918
rect 442698 2682 442782 2918
rect 443018 2682 443102 2918
rect 443338 2682 443422 2918
rect 443658 2682 443742 2918
rect 443978 2682 444062 2918
rect 444298 2682 444382 2918
rect 444618 2682 444740 2918
rect 440740 2598 444740 2682
rect 440740 2362 440862 2598
rect 441098 2362 441182 2598
rect 441418 2362 441502 2598
rect 441738 2362 441822 2598
rect 442058 2362 442142 2598
rect 442378 2362 442462 2598
rect 442698 2362 442782 2598
rect 443018 2362 443102 2598
rect 443338 2362 443422 2598
rect 443658 2362 443742 2598
rect 443978 2362 444062 2598
rect 444298 2362 444382 2598
rect 444618 2362 444740 2598
rect 440740 2278 444740 2362
rect 440740 2042 440862 2278
rect 441098 2042 441182 2278
rect 441418 2042 441502 2278
rect 441738 2042 441822 2278
rect 442058 2042 442142 2278
rect 442378 2042 442462 2278
rect 442698 2042 442782 2278
rect 443018 2042 443102 2278
rect 443338 2042 443422 2278
rect 443658 2042 443742 2278
rect 443978 2042 444062 2278
rect 444298 2042 444382 2278
rect 444618 2042 444740 2278
rect 440740 1958 444740 2042
rect 440740 1722 440862 1958
rect 441098 1722 441182 1958
rect 441418 1722 441502 1958
rect 441738 1722 441822 1958
rect 442058 1722 442142 1958
rect 442378 1722 442462 1958
rect 442698 1722 442782 1958
rect 443018 1722 443102 1958
rect 443338 1722 443422 1958
rect 443658 1722 443742 1958
rect 443978 1722 444062 1958
rect 444298 1722 444382 1958
rect 444618 1722 444740 1958
rect 440740 1638 444740 1722
rect 440740 1402 440862 1638
rect 441098 1402 441182 1638
rect 441418 1402 441502 1638
rect 441738 1402 441822 1638
rect 442058 1402 442142 1638
rect 442378 1402 442462 1638
rect 442698 1402 442782 1638
rect 443018 1402 443102 1638
rect 443338 1402 443422 1638
rect 443658 1402 443742 1638
rect 443978 1402 444062 1638
rect 444298 1402 444382 1638
rect 444618 1402 444740 1638
rect 440740 1318 444740 1402
rect 440740 1082 440862 1318
rect 441098 1082 441182 1318
rect 441418 1082 441502 1318
rect 441738 1082 441822 1318
rect 442058 1082 442142 1318
rect 442378 1082 442462 1318
rect 442698 1082 442782 1318
rect 443018 1082 443102 1318
rect 443338 1082 443422 1318
rect 443658 1082 443742 1318
rect 443978 1082 444062 1318
rect 444298 1082 444382 1318
rect 444618 1082 444740 1318
rect 440740 998 444740 1082
rect 440740 762 440862 998
rect 441098 762 441182 998
rect 441418 762 441502 998
rect 441738 762 441822 998
rect 442058 762 442142 998
rect 442378 762 442462 998
rect 442698 762 442782 998
rect 443018 762 443102 998
rect 443338 762 443422 998
rect 443658 762 443742 998
rect 443978 762 444062 998
rect 444298 762 444382 998
rect 444618 762 444740 998
rect 440740 678 444740 762
rect 440740 442 440862 678
rect 441098 442 441182 678
rect 441418 442 441502 678
rect 441738 442 441822 678
rect 442058 442 442142 678
rect 442378 442 442462 678
rect 442698 442 442782 678
rect 443018 442 443102 678
rect 443338 442 443422 678
rect 443658 442 443742 678
rect 443978 442 444062 678
rect 444298 442 444382 678
rect 444618 442 444740 678
rect 440740 358 444740 442
rect 440740 122 440862 358
rect 441098 122 441182 358
rect 441418 122 441502 358
rect 441738 122 441822 358
rect 442058 122 442142 358
rect 442378 122 442462 358
rect 442698 122 442782 358
rect 443018 122 443102 358
rect 443338 122 443422 358
rect 443658 122 443742 358
rect 443978 122 444062 358
rect 444298 122 444382 358
rect 444618 122 444740 358
rect 440740 0 444740 122
<< via4 >>
rect 122 405162 358 405398
rect 442 405162 678 405398
rect 762 405162 998 405398
rect 1082 405162 1318 405398
rect 1402 405162 1638 405398
rect 1722 405162 1958 405398
rect 2042 405162 2278 405398
rect 2362 405162 2598 405398
rect 2682 405162 2918 405398
rect 3002 405162 3238 405398
rect 3322 405162 3558 405398
rect 3642 405162 3878 405398
rect 122 404842 358 405078
rect 442 404842 678 405078
rect 762 404842 998 405078
rect 1082 404842 1318 405078
rect 1402 404842 1638 405078
rect 1722 404842 1958 405078
rect 2042 404842 2278 405078
rect 2362 404842 2598 405078
rect 2682 404842 2918 405078
rect 3002 404842 3238 405078
rect 3322 404842 3558 405078
rect 3642 404842 3878 405078
rect 122 404522 358 404758
rect 442 404522 678 404758
rect 762 404522 998 404758
rect 1082 404522 1318 404758
rect 1402 404522 1638 404758
rect 1722 404522 1958 404758
rect 2042 404522 2278 404758
rect 2362 404522 2598 404758
rect 2682 404522 2918 404758
rect 3002 404522 3238 404758
rect 3322 404522 3558 404758
rect 3642 404522 3878 404758
rect 122 404202 358 404438
rect 442 404202 678 404438
rect 762 404202 998 404438
rect 1082 404202 1318 404438
rect 1402 404202 1638 404438
rect 1722 404202 1958 404438
rect 2042 404202 2278 404438
rect 2362 404202 2598 404438
rect 2682 404202 2918 404438
rect 3002 404202 3238 404438
rect 3322 404202 3558 404438
rect 3642 404202 3878 404438
rect 122 403882 358 404118
rect 442 403882 678 404118
rect 762 403882 998 404118
rect 1082 403882 1318 404118
rect 1402 403882 1638 404118
rect 1722 403882 1958 404118
rect 2042 403882 2278 404118
rect 2362 403882 2598 404118
rect 2682 403882 2918 404118
rect 3002 403882 3238 404118
rect 3322 403882 3558 404118
rect 3642 403882 3878 404118
rect 122 403562 358 403798
rect 442 403562 678 403798
rect 762 403562 998 403798
rect 1082 403562 1318 403798
rect 1402 403562 1638 403798
rect 1722 403562 1958 403798
rect 2042 403562 2278 403798
rect 2362 403562 2598 403798
rect 2682 403562 2918 403798
rect 3002 403562 3238 403798
rect 3322 403562 3558 403798
rect 3642 403562 3878 403798
rect 122 403242 358 403478
rect 442 403242 678 403478
rect 762 403242 998 403478
rect 1082 403242 1318 403478
rect 1402 403242 1638 403478
rect 1722 403242 1958 403478
rect 2042 403242 2278 403478
rect 2362 403242 2598 403478
rect 2682 403242 2918 403478
rect 3002 403242 3238 403478
rect 3322 403242 3558 403478
rect 3642 403242 3878 403478
rect 122 402922 358 403158
rect 442 402922 678 403158
rect 762 402922 998 403158
rect 1082 402922 1318 403158
rect 1402 402922 1638 403158
rect 1722 402922 1958 403158
rect 2042 402922 2278 403158
rect 2362 402922 2598 403158
rect 2682 402922 2918 403158
rect 3002 402922 3238 403158
rect 3322 402922 3558 403158
rect 3642 402922 3878 403158
rect 122 402602 358 402838
rect 442 402602 678 402838
rect 762 402602 998 402838
rect 1082 402602 1318 402838
rect 1402 402602 1638 402838
rect 1722 402602 1958 402838
rect 2042 402602 2278 402838
rect 2362 402602 2598 402838
rect 2682 402602 2918 402838
rect 3002 402602 3238 402838
rect 3322 402602 3558 402838
rect 3642 402602 3878 402838
rect 122 402282 358 402518
rect 442 402282 678 402518
rect 762 402282 998 402518
rect 1082 402282 1318 402518
rect 1402 402282 1638 402518
rect 1722 402282 1958 402518
rect 2042 402282 2278 402518
rect 2362 402282 2598 402518
rect 2682 402282 2918 402518
rect 3002 402282 3238 402518
rect 3322 402282 3558 402518
rect 3642 402282 3878 402518
rect 122 401962 358 402198
rect 442 401962 678 402198
rect 762 401962 998 402198
rect 1082 401962 1318 402198
rect 1402 401962 1638 402198
rect 1722 401962 1958 402198
rect 2042 401962 2278 402198
rect 2362 401962 2598 402198
rect 2682 401962 2918 402198
rect 3002 401962 3238 402198
rect 3322 401962 3558 402198
rect 3642 401962 3878 402198
rect 122 401642 358 401878
rect 442 401642 678 401878
rect 762 401642 998 401878
rect 1082 401642 1318 401878
rect 1402 401642 1638 401878
rect 1722 401642 1958 401878
rect 2042 401642 2278 401878
rect 2362 401642 2598 401878
rect 2682 401642 2918 401878
rect 3002 401642 3238 401878
rect 3322 401642 3558 401878
rect 3642 401642 3878 401878
rect 440862 405162 441098 405398
rect 441182 405162 441418 405398
rect 441502 405162 441738 405398
rect 441822 405162 442058 405398
rect 442142 405162 442378 405398
rect 442462 405162 442698 405398
rect 442782 405162 443018 405398
rect 443102 405162 443338 405398
rect 443422 405162 443658 405398
rect 443742 405162 443978 405398
rect 444062 405162 444298 405398
rect 444382 405162 444618 405398
rect 440862 404842 441098 405078
rect 441182 404842 441418 405078
rect 441502 404842 441738 405078
rect 441822 404842 442058 405078
rect 442142 404842 442378 405078
rect 442462 404842 442698 405078
rect 442782 404842 443018 405078
rect 443102 404842 443338 405078
rect 443422 404842 443658 405078
rect 443742 404842 443978 405078
rect 444062 404842 444298 405078
rect 444382 404842 444618 405078
rect 440862 404522 441098 404758
rect 441182 404522 441418 404758
rect 441502 404522 441738 404758
rect 441822 404522 442058 404758
rect 442142 404522 442378 404758
rect 442462 404522 442698 404758
rect 442782 404522 443018 404758
rect 443102 404522 443338 404758
rect 443422 404522 443658 404758
rect 443742 404522 443978 404758
rect 444062 404522 444298 404758
rect 444382 404522 444618 404758
rect 440862 404202 441098 404438
rect 441182 404202 441418 404438
rect 441502 404202 441738 404438
rect 441822 404202 442058 404438
rect 442142 404202 442378 404438
rect 442462 404202 442698 404438
rect 442782 404202 443018 404438
rect 443102 404202 443338 404438
rect 443422 404202 443658 404438
rect 443742 404202 443978 404438
rect 444062 404202 444298 404438
rect 444382 404202 444618 404438
rect 440862 403882 441098 404118
rect 441182 403882 441418 404118
rect 441502 403882 441738 404118
rect 441822 403882 442058 404118
rect 442142 403882 442378 404118
rect 442462 403882 442698 404118
rect 442782 403882 443018 404118
rect 443102 403882 443338 404118
rect 443422 403882 443658 404118
rect 443742 403882 443978 404118
rect 444062 403882 444298 404118
rect 444382 403882 444618 404118
rect 440862 403562 441098 403798
rect 441182 403562 441418 403798
rect 441502 403562 441738 403798
rect 441822 403562 442058 403798
rect 442142 403562 442378 403798
rect 442462 403562 442698 403798
rect 442782 403562 443018 403798
rect 443102 403562 443338 403798
rect 443422 403562 443658 403798
rect 443742 403562 443978 403798
rect 444062 403562 444298 403798
rect 444382 403562 444618 403798
rect 440862 403242 441098 403478
rect 441182 403242 441418 403478
rect 441502 403242 441738 403478
rect 441822 403242 442058 403478
rect 442142 403242 442378 403478
rect 442462 403242 442698 403478
rect 442782 403242 443018 403478
rect 443102 403242 443338 403478
rect 443422 403242 443658 403478
rect 443742 403242 443978 403478
rect 444062 403242 444298 403478
rect 444382 403242 444618 403478
rect 440862 402922 441098 403158
rect 441182 402922 441418 403158
rect 441502 402922 441738 403158
rect 441822 402922 442058 403158
rect 442142 402922 442378 403158
rect 442462 402922 442698 403158
rect 442782 402922 443018 403158
rect 443102 402922 443338 403158
rect 443422 402922 443658 403158
rect 443742 402922 443978 403158
rect 444062 402922 444298 403158
rect 444382 402922 444618 403158
rect 440862 402602 441098 402838
rect 441182 402602 441418 402838
rect 441502 402602 441738 402838
rect 441822 402602 442058 402838
rect 442142 402602 442378 402838
rect 442462 402602 442698 402838
rect 442782 402602 443018 402838
rect 443102 402602 443338 402838
rect 443422 402602 443658 402838
rect 443742 402602 443978 402838
rect 444062 402602 444298 402838
rect 444382 402602 444618 402838
rect 440862 402282 441098 402518
rect 441182 402282 441418 402518
rect 441502 402282 441738 402518
rect 441822 402282 442058 402518
rect 442142 402282 442378 402518
rect 442462 402282 442698 402518
rect 442782 402282 443018 402518
rect 443102 402282 443338 402518
rect 443422 402282 443658 402518
rect 443742 402282 443978 402518
rect 444062 402282 444298 402518
rect 444382 402282 444618 402518
rect 440862 401962 441098 402198
rect 441182 401962 441418 402198
rect 441502 401962 441738 402198
rect 441822 401962 442058 402198
rect 442142 401962 442378 402198
rect 442462 401962 442698 402198
rect 442782 401962 443018 402198
rect 443102 401962 443338 402198
rect 443422 401962 443658 402198
rect 443742 401962 443978 402198
rect 444062 401962 444298 402198
rect 444382 401962 444618 402198
rect 440862 401642 441098 401878
rect 441182 401642 441418 401878
rect 441502 401642 441738 401878
rect 441822 401642 442058 401878
rect 442142 401642 442378 401878
rect 442462 401642 442698 401878
rect 442782 401642 443018 401878
rect 443102 401642 443338 401878
rect 443422 401642 443658 401878
rect 443742 401642 443978 401878
rect 444062 401642 444298 401878
rect 444382 401642 444618 401878
rect 122 376196 358 376432
rect 442 376196 678 376432
rect 762 376196 998 376432
rect 1082 376196 1318 376432
rect 1402 376196 1638 376432
rect 1722 376196 1958 376432
rect 2042 376196 2278 376432
rect 2362 376196 2598 376432
rect 2682 376196 2918 376432
rect 3002 376196 3238 376432
rect 3322 376196 3558 376432
rect 3642 376196 3878 376432
rect 122 345560 358 345796
rect 442 345560 678 345796
rect 762 345560 998 345796
rect 1082 345560 1318 345796
rect 1402 345560 1638 345796
rect 1722 345560 1958 345796
rect 2042 345560 2278 345796
rect 2362 345560 2598 345796
rect 2682 345560 2918 345796
rect 3002 345560 3238 345796
rect 3322 345560 3558 345796
rect 3642 345560 3878 345796
rect 122 314924 358 315160
rect 442 314924 678 315160
rect 762 314924 998 315160
rect 1082 314924 1318 315160
rect 1402 314924 1638 315160
rect 1722 314924 1958 315160
rect 2042 314924 2278 315160
rect 2362 314924 2598 315160
rect 2682 314924 2918 315160
rect 3002 314924 3238 315160
rect 3322 314924 3558 315160
rect 3642 314924 3878 315160
rect 122 284288 358 284524
rect 442 284288 678 284524
rect 762 284288 998 284524
rect 1082 284288 1318 284524
rect 1402 284288 1638 284524
rect 1722 284288 1958 284524
rect 2042 284288 2278 284524
rect 2362 284288 2598 284524
rect 2682 284288 2918 284524
rect 3002 284288 3238 284524
rect 3322 284288 3558 284524
rect 3642 284288 3878 284524
rect 122 253652 358 253888
rect 442 253652 678 253888
rect 762 253652 998 253888
rect 1082 253652 1318 253888
rect 1402 253652 1638 253888
rect 1722 253652 1958 253888
rect 2042 253652 2278 253888
rect 2362 253652 2598 253888
rect 2682 253652 2918 253888
rect 3002 253652 3238 253888
rect 3322 253652 3558 253888
rect 3642 253652 3878 253888
rect 122 223016 358 223252
rect 442 223016 678 223252
rect 762 223016 998 223252
rect 1082 223016 1318 223252
rect 1402 223016 1638 223252
rect 1722 223016 1958 223252
rect 2042 223016 2278 223252
rect 2362 223016 2598 223252
rect 2682 223016 2918 223252
rect 3002 223016 3238 223252
rect 3322 223016 3558 223252
rect 3642 223016 3878 223252
rect 122 192380 358 192616
rect 442 192380 678 192616
rect 762 192380 998 192616
rect 1082 192380 1318 192616
rect 1402 192380 1638 192616
rect 1722 192380 1958 192616
rect 2042 192380 2278 192616
rect 2362 192380 2598 192616
rect 2682 192380 2918 192616
rect 3002 192380 3238 192616
rect 3322 192380 3558 192616
rect 3642 192380 3878 192616
rect 122 161744 358 161980
rect 442 161744 678 161980
rect 762 161744 998 161980
rect 1082 161744 1318 161980
rect 1402 161744 1638 161980
rect 1722 161744 1958 161980
rect 2042 161744 2278 161980
rect 2362 161744 2598 161980
rect 2682 161744 2918 161980
rect 3002 161744 3238 161980
rect 3322 161744 3558 161980
rect 3642 161744 3878 161980
rect 122 131108 358 131344
rect 442 131108 678 131344
rect 762 131108 998 131344
rect 1082 131108 1318 131344
rect 1402 131108 1638 131344
rect 1722 131108 1958 131344
rect 2042 131108 2278 131344
rect 2362 131108 2598 131344
rect 2682 131108 2918 131344
rect 3002 131108 3238 131344
rect 3322 131108 3558 131344
rect 3642 131108 3878 131344
rect 122 100472 358 100708
rect 442 100472 678 100708
rect 762 100472 998 100708
rect 1082 100472 1318 100708
rect 1402 100472 1638 100708
rect 1722 100472 1958 100708
rect 2042 100472 2278 100708
rect 2362 100472 2598 100708
rect 2682 100472 2918 100708
rect 3002 100472 3238 100708
rect 3322 100472 3558 100708
rect 3642 100472 3878 100708
rect 122 69836 358 70072
rect 442 69836 678 70072
rect 762 69836 998 70072
rect 1082 69836 1318 70072
rect 1402 69836 1638 70072
rect 1722 69836 1958 70072
rect 2042 69836 2278 70072
rect 2362 69836 2598 70072
rect 2682 69836 2918 70072
rect 3002 69836 3238 70072
rect 3322 69836 3558 70072
rect 3642 69836 3878 70072
rect 122 39200 358 39436
rect 442 39200 678 39436
rect 762 39200 998 39436
rect 1082 39200 1318 39436
rect 1402 39200 1638 39436
rect 1722 39200 1958 39436
rect 2042 39200 2278 39436
rect 2362 39200 2598 39436
rect 2682 39200 2918 39436
rect 3002 39200 3238 39436
rect 3322 39200 3558 39436
rect 3642 39200 3878 39436
rect 5122 400162 5358 400398
rect 5442 400162 5678 400398
rect 5762 400162 5998 400398
rect 6082 400162 6318 400398
rect 6402 400162 6638 400398
rect 6722 400162 6958 400398
rect 7042 400162 7278 400398
rect 7362 400162 7598 400398
rect 7682 400162 7918 400398
rect 8002 400162 8238 400398
rect 8322 400162 8558 400398
rect 8642 400162 8878 400398
rect 5122 399842 5358 400078
rect 5442 399842 5678 400078
rect 5762 399842 5998 400078
rect 6082 399842 6318 400078
rect 6402 399842 6638 400078
rect 6722 399842 6958 400078
rect 7042 399842 7278 400078
rect 7362 399842 7598 400078
rect 7682 399842 7918 400078
rect 8002 399842 8238 400078
rect 8322 399842 8558 400078
rect 8642 399842 8878 400078
rect 5122 399522 5358 399758
rect 5442 399522 5678 399758
rect 5762 399522 5998 399758
rect 6082 399522 6318 399758
rect 6402 399522 6638 399758
rect 6722 399522 6958 399758
rect 7042 399522 7278 399758
rect 7362 399522 7598 399758
rect 7682 399522 7918 399758
rect 8002 399522 8238 399758
rect 8322 399522 8558 399758
rect 8642 399522 8878 399758
rect 5122 399202 5358 399438
rect 5442 399202 5678 399438
rect 5762 399202 5998 399438
rect 6082 399202 6318 399438
rect 6402 399202 6638 399438
rect 6722 399202 6958 399438
rect 7042 399202 7278 399438
rect 7362 399202 7598 399438
rect 7682 399202 7918 399438
rect 8002 399202 8238 399438
rect 8322 399202 8558 399438
rect 8642 399202 8878 399438
rect 5122 398882 5358 399118
rect 5442 398882 5678 399118
rect 5762 398882 5998 399118
rect 6082 398882 6318 399118
rect 6402 398882 6638 399118
rect 6722 398882 6958 399118
rect 7042 398882 7278 399118
rect 7362 398882 7598 399118
rect 7682 398882 7918 399118
rect 8002 398882 8238 399118
rect 8322 398882 8558 399118
rect 8642 398882 8878 399118
rect 5122 398562 5358 398798
rect 5442 398562 5678 398798
rect 5762 398562 5998 398798
rect 6082 398562 6318 398798
rect 6402 398562 6638 398798
rect 6722 398562 6958 398798
rect 7042 398562 7278 398798
rect 7362 398562 7598 398798
rect 7682 398562 7918 398798
rect 8002 398562 8238 398798
rect 8322 398562 8558 398798
rect 8642 398562 8878 398798
rect 5122 398242 5358 398478
rect 5442 398242 5678 398478
rect 5762 398242 5998 398478
rect 6082 398242 6318 398478
rect 6402 398242 6638 398478
rect 6722 398242 6958 398478
rect 7042 398242 7278 398478
rect 7362 398242 7598 398478
rect 7682 398242 7918 398478
rect 8002 398242 8238 398478
rect 8322 398242 8558 398478
rect 8642 398242 8878 398478
rect 5122 397922 5358 398158
rect 5442 397922 5678 398158
rect 5762 397922 5998 398158
rect 6082 397922 6318 398158
rect 6402 397922 6638 398158
rect 6722 397922 6958 398158
rect 7042 397922 7278 398158
rect 7362 397922 7598 398158
rect 7682 397922 7918 398158
rect 8002 397922 8238 398158
rect 8322 397922 8558 398158
rect 8642 397922 8878 398158
rect 5122 397602 5358 397838
rect 5442 397602 5678 397838
rect 5762 397602 5998 397838
rect 6082 397602 6318 397838
rect 6402 397602 6638 397838
rect 6722 397602 6958 397838
rect 7042 397602 7278 397838
rect 7362 397602 7598 397838
rect 7682 397602 7918 397838
rect 8002 397602 8238 397838
rect 8322 397602 8558 397838
rect 8642 397602 8878 397838
rect 5122 397282 5358 397518
rect 5442 397282 5678 397518
rect 5762 397282 5998 397518
rect 6082 397282 6318 397518
rect 6402 397282 6638 397518
rect 6722 397282 6958 397518
rect 7042 397282 7278 397518
rect 7362 397282 7598 397518
rect 7682 397282 7918 397518
rect 8002 397282 8238 397518
rect 8322 397282 8558 397518
rect 8642 397282 8878 397518
rect 5122 396962 5358 397198
rect 5442 396962 5678 397198
rect 5762 396962 5998 397198
rect 6082 396962 6318 397198
rect 6402 396962 6638 397198
rect 6722 396962 6958 397198
rect 7042 396962 7278 397198
rect 7362 396962 7598 397198
rect 7682 396962 7918 397198
rect 8002 396962 8238 397198
rect 8322 396962 8558 397198
rect 8642 396962 8878 397198
rect 5122 396642 5358 396878
rect 5442 396642 5678 396878
rect 5762 396642 5998 396878
rect 6082 396642 6318 396878
rect 6402 396642 6638 396878
rect 6722 396642 6958 396878
rect 7042 396642 7278 396878
rect 7362 396642 7598 396878
rect 7682 396642 7918 396878
rect 8002 396642 8238 396878
rect 8322 396642 8558 396878
rect 8642 396642 8878 396878
rect 435862 400162 436098 400398
rect 436182 400162 436418 400398
rect 436502 400162 436738 400398
rect 436822 400162 437058 400398
rect 437142 400162 437378 400398
rect 437462 400162 437698 400398
rect 437782 400162 438018 400398
rect 438102 400162 438338 400398
rect 438422 400162 438658 400398
rect 438742 400162 438978 400398
rect 439062 400162 439298 400398
rect 439382 400162 439618 400398
rect 435862 399842 436098 400078
rect 436182 399842 436418 400078
rect 436502 399842 436738 400078
rect 436822 399842 437058 400078
rect 437142 399842 437378 400078
rect 437462 399842 437698 400078
rect 437782 399842 438018 400078
rect 438102 399842 438338 400078
rect 438422 399842 438658 400078
rect 438742 399842 438978 400078
rect 439062 399842 439298 400078
rect 439382 399842 439618 400078
rect 435862 399522 436098 399758
rect 436182 399522 436418 399758
rect 436502 399522 436738 399758
rect 436822 399522 437058 399758
rect 437142 399522 437378 399758
rect 437462 399522 437698 399758
rect 437782 399522 438018 399758
rect 438102 399522 438338 399758
rect 438422 399522 438658 399758
rect 438742 399522 438978 399758
rect 439062 399522 439298 399758
rect 439382 399522 439618 399758
rect 435862 399202 436098 399438
rect 436182 399202 436418 399438
rect 436502 399202 436738 399438
rect 436822 399202 437058 399438
rect 437142 399202 437378 399438
rect 437462 399202 437698 399438
rect 437782 399202 438018 399438
rect 438102 399202 438338 399438
rect 438422 399202 438658 399438
rect 438742 399202 438978 399438
rect 439062 399202 439298 399438
rect 439382 399202 439618 399438
rect 435862 398882 436098 399118
rect 436182 398882 436418 399118
rect 436502 398882 436738 399118
rect 436822 398882 437058 399118
rect 437142 398882 437378 399118
rect 437462 398882 437698 399118
rect 437782 398882 438018 399118
rect 438102 398882 438338 399118
rect 438422 398882 438658 399118
rect 438742 398882 438978 399118
rect 439062 398882 439298 399118
rect 439382 398882 439618 399118
rect 435862 398562 436098 398798
rect 436182 398562 436418 398798
rect 436502 398562 436738 398798
rect 436822 398562 437058 398798
rect 437142 398562 437378 398798
rect 437462 398562 437698 398798
rect 437782 398562 438018 398798
rect 438102 398562 438338 398798
rect 438422 398562 438658 398798
rect 438742 398562 438978 398798
rect 439062 398562 439298 398798
rect 439382 398562 439618 398798
rect 435862 398242 436098 398478
rect 436182 398242 436418 398478
rect 436502 398242 436738 398478
rect 436822 398242 437058 398478
rect 437142 398242 437378 398478
rect 437462 398242 437698 398478
rect 437782 398242 438018 398478
rect 438102 398242 438338 398478
rect 438422 398242 438658 398478
rect 438742 398242 438978 398478
rect 439062 398242 439298 398478
rect 439382 398242 439618 398478
rect 435862 397922 436098 398158
rect 436182 397922 436418 398158
rect 436502 397922 436738 398158
rect 436822 397922 437058 398158
rect 437142 397922 437378 398158
rect 437462 397922 437698 398158
rect 437782 397922 438018 398158
rect 438102 397922 438338 398158
rect 438422 397922 438658 398158
rect 438742 397922 438978 398158
rect 439062 397922 439298 398158
rect 439382 397922 439618 398158
rect 435862 397602 436098 397838
rect 436182 397602 436418 397838
rect 436502 397602 436738 397838
rect 436822 397602 437058 397838
rect 437142 397602 437378 397838
rect 437462 397602 437698 397838
rect 437782 397602 438018 397838
rect 438102 397602 438338 397838
rect 438422 397602 438658 397838
rect 438742 397602 438978 397838
rect 439062 397602 439298 397838
rect 439382 397602 439618 397838
rect 435862 397282 436098 397518
rect 436182 397282 436418 397518
rect 436502 397282 436738 397518
rect 436822 397282 437058 397518
rect 437142 397282 437378 397518
rect 437462 397282 437698 397518
rect 437782 397282 438018 397518
rect 438102 397282 438338 397518
rect 438422 397282 438658 397518
rect 438742 397282 438978 397518
rect 439062 397282 439298 397518
rect 439382 397282 439618 397518
rect 435862 396962 436098 397198
rect 436182 396962 436418 397198
rect 436502 396962 436738 397198
rect 436822 396962 437058 397198
rect 437142 396962 437378 397198
rect 437462 396962 437698 397198
rect 437782 396962 438018 397198
rect 438102 396962 438338 397198
rect 438422 396962 438658 397198
rect 438742 396962 438978 397198
rect 439062 396962 439298 397198
rect 439382 396962 439618 397198
rect 435862 396642 436098 396878
rect 436182 396642 436418 396878
rect 436502 396642 436738 396878
rect 436822 396642 437058 396878
rect 437142 396642 437378 396878
rect 437462 396642 437698 396878
rect 437782 396642 438018 396878
rect 438102 396642 438338 396878
rect 438422 396642 438658 396878
rect 438742 396642 438978 396878
rect 439062 396642 439298 396878
rect 439382 396642 439618 396878
rect 5122 391514 5358 391750
rect 5442 391514 5678 391750
rect 5762 391514 5998 391750
rect 6082 391514 6318 391750
rect 6402 391514 6638 391750
rect 6722 391514 6958 391750
rect 7042 391514 7278 391750
rect 7362 391514 7598 391750
rect 7682 391514 7918 391750
rect 8002 391514 8238 391750
rect 8322 391514 8558 391750
rect 8642 391514 8878 391750
rect 5122 360878 5358 361114
rect 5442 360878 5678 361114
rect 5762 360878 5998 361114
rect 6082 360878 6318 361114
rect 6402 360878 6638 361114
rect 6722 360878 6958 361114
rect 7042 360878 7278 361114
rect 7362 360878 7598 361114
rect 7682 360878 7918 361114
rect 8002 360878 8238 361114
rect 8322 360878 8558 361114
rect 8642 360878 8878 361114
rect 5122 330242 5358 330478
rect 5442 330242 5678 330478
rect 5762 330242 5998 330478
rect 6082 330242 6318 330478
rect 6402 330242 6638 330478
rect 6722 330242 6958 330478
rect 7042 330242 7278 330478
rect 7362 330242 7598 330478
rect 7682 330242 7918 330478
rect 8002 330242 8238 330478
rect 8322 330242 8558 330478
rect 8642 330242 8878 330478
rect 231774 333556 232010 333642
rect 231774 333492 231860 333556
rect 231860 333492 231924 333556
rect 231924 333492 232010 333556
rect 137198 332196 137434 332282
rect 137198 332132 137284 332196
rect 137284 332132 137348 332196
rect 137348 332132 137434 332196
rect 137198 332046 137434 332132
rect 168478 332046 168714 332282
rect 198654 332196 198890 332282
rect 198654 332132 198740 332196
rect 198740 332132 198804 332196
rect 198804 332132 198890 332196
rect 198654 332046 198890 332132
rect 137198 331516 137434 331602
rect 137198 331452 137284 331516
rect 137284 331452 137348 331516
rect 137348 331452 137434 331516
rect 137198 331366 137434 331452
rect 159462 331366 159698 331602
rect 161670 329476 161906 329562
rect 161670 329412 161756 329476
rect 161756 329412 161820 329476
rect 161820 329412 161906 329476
rect 161670 329326 161906 329412
rect 204358 331588 204444 331602
rect 204444 331588 204508 331602
rect 204508 331588 204594 331602
rect 204358 331366 204594 331588
rect 231774 333406 232010 333492
rect 262318 333406 262554 333642
rect 231774 332196 232010 332282
rect 231774 332132 231860 332196
rect 231860 332132 231924 332196
rect 231924 332132 232010 332196
rect 231774 332046 232010 332132
rect 231774 331516 232010 331602
rect 231774 331452 231860 331516
rect 231860 331452 231924 331516
rect 231924 331452 232010 331516
rect 231774 331366 232010 331452
rect 251462 331366 251698 331602
rect 252198 331366 252434 331602
rect 252934 331366 253170 331602
rect 212086 329326 212322 329562
rect 306110 333556 306346 333642
rect 306110 333492 306196 333556
rect 306196 333492 306260 333556
rect 306260 333492 306346 333556
rect 306110 333406 306346 333492
rect 295990 332196 296226 332282
rect 295990 332132 296076 332196
rect 296076 332132 296140 332196
rect 296140 332132 296226 332196
rect 295990 332046 296226 332132
rect 293966 331588 294052 331602
rect 294052 331588 294116 331602
rect 294116 331588 294202 331602
rect 293966 331366 294202 331588
rect 104814 319806 105050 320042
rect 5122 299606 5358 299842
rect 5442 299606 5678 299842
rect 5762 299606 5998 299842
rect 6082 299606 6318 299842
rect 6402 299606 6638 299842
rect 6722 299606 6958 299842
rect 7042 299606 7278 299842
rect 7362 299606 7598 299842
rect 7682 299606 7918 299842
rect 8002 299606 8238 299842
rect 8322 299606 8558 299842
rect 8642 299606 8878 299842
rect 5122 268970 5358 269206
rect 5442 268970 5678 269206
rect 5762 268970 5998 269206
rect 6082 268970 6318 269206
rect 6402 268970 6638 269206
rect 6722 268970 6958 269206
rect 7042 268970 7278 269206
rect 7362 268970 7598 269206
rect 7682 268970 7918 269206
rect 8002 268970 8238 269206
rect 8322 268970 8558 269206
rect 8642 268970 8878 269206
rect 104630 315726 104866 315962
rect 104506 314924 104742 315160
rect 198506 314924 198742 315160
rect 292506 314924 292742 315160
rect 104630 314366 104866 314602
rect 48878 259436 49114 259522
rect 48878 259372 48964 259436
rect 48964 259372 49028 259436
rect 49028 259372 49114 259436
rect 48878 259286 49114 259372
rect 48878 255900 49114 256122
rect 48878 255886 48964 255900
rect 48964 255886 49028 255900
rect 49028 255886 49114 255900
rect 48878 249236 49114 249322
rect 48878 249172 48964 249236
rect 48964 249172 49028 249236
rect 49028 249172 49114 249236
rect 48878 249086 49114 249172
rect 46854 242286 47090 242522
rect 49062 240926 49298 241162
rect 49062 239788 49148 239802
rect 49148 239788 49212 239802
rect 49212 239788 49298 239802
rect 49062 239566 49298 239788
rect 5122 238334 5358 238570
rect 5442 238334 5678 238570
rect 5762 238334 5998 238570
rect 6082 238334 6318 238570
rect 6402 238334 6638 238570
rect 6722 238334 6958 238570
rect 7042 238334 7278 238570
rect 7362 238334 7598 238570
rect 7682 238334 7918 238570
rect 8002 238334 8238 238570
rect 8322 238334 8558 238570
rect 8642 238334 8878 238570
rect 5122 207698 5358 207934
rect 5442 207698 5678 207934
rect 5762 207698 5998 207934
rect 6082 207698 6318 207934
rect 6402 207698 6638 207934
rect 6722 207698 6958 207934
rect 7042 207698 7278 207934
rect 7362 207698 7598 207934
rect 7682 207698 7918 207934
rect 8002 207698 8238 207934
rect 8322 207698 8558 207934
rect 8642 207698 8878 207934
rect 5122 177062 5358 177298
rect 5442 177062 5678 177298
rect 5762 177062 5998 177298
rect 6082 177062 6318 177298
rect 6402 177062 6638 177298
rect 6722 177062 6958 177298
rect 7042 177062 7278 177298
rect 7362 177062 7598 177298
rect 7682 177062 7918 177298
rect 8002 177062 8238 177298
rect 8322 177062 8558 177298
rect 8642 177062 8878 177298
rect 104630 300766 104866 301002
rect 89146 299606 89382 299842
rect 104446 299406 104682 299642
rect 183146 299606 183382 299842
rect 277146 299606 277382 299842
rect 134622 298196 134858 298282
rect 134622 298132 134708 298196
rect 134708 298132 134772 298196
rect 134772 298132 134858 298196
rect 134622 298046 134858 298132
rect 231774 295326 232010 295562
rect 136830 294796 137066 294882
rect 136830 294732 136916 294796
rect 136916 294732 136980 294796
rect 136980 294732 137066 294796
rect 136830 294646 137066 294732
rect 228646 294796 228882 294882
rect 228646 294732 228732 294796
rect 228732 294732 228796 294796
rect 228796 294732 228882 294796
rect 228646 294646 228882 294732
rect 136830 292148 136916 292162
rect 136916 292148 136980 292162
rect 136980 292148 137066 292162
rect 136830 291926 137066 292148
rect 230670 292076 230906 292162
rect 230670 292012 230756 292076
rect 230756 292012 230820 292076
rect 230820 292012 230906 292076
rect 230670 291926 230906 292012
rect 322670 291940 322906 292162
rect 322670 291926 322756 291940
rect 322756 291926 322820 291940
rect 322820 291926 322906 291940
rect 261030 290716 261266 290802
rect 261030 290652 261116 290716
rect 261116 290652 261180 290716
rect 261180 290652 261266 290716
rect 261030 290566 261266 290652
rect 435862 391514 436098 391750
rect 436182 391514 436418 391750
rect 436502 391514 436738 391750
rect 436822 391514 437058 391750
rect 437142 391514 437378 391750
rect 437462 391514 437698 391750
rect 437782 391514 438018 391750
rect 438102 391514 438338 391750
rect 438422 391514 438658 391750
rect 438742 391514 438978 391750
rect 439062 391514 439298 391750
rect 439382 391514 439618 391750
rect 435862 360878 436098 361114
rect 436182 360878 436418 361114
rect 436502 360878 436738 361114
rect 436822 360878 437058 361114
rect 437142 360878 437378 361114
rect 437462 360878 437698 361114
rect 437782 360878 438018 361114
rect 438102 360878 438338 361114
rect 438422 360878 438658 361114
rect 438742 360878 438978 361114
rect 439062 360878 439298 361114
rect 439382 360878 439618 361114
rect 435862 330242 436098 330478
rect 436182 330242 436418 330478
rect 436502 330242 436738 330478
rect 436822 330242 437058 330478
rect 437142 330242 437378 330478
rect 437462 330242 437698 330478
rect 437782 330242 438018 330478
rect 438102 330242 438338 330478
rect 438422 330242 438658 330478
rect 438742 330242 438978 330478
rect 439062 330242 439298 330478
rect 439382 330242 439618 330478
rect 323406 295476 323642 295562
rect 323406 295412 323492 295476
rect 323492 295412 323556 295476
rect 323556 295412 323642 295476
rect 323406 295326 323642 295412
rect 137934 289356 138170 289442
rect 137934 289292 138020 289356
rect 138020 289292 138084 289356
rect 138084 289292 138170 289356
rect 137934 289206 138170 289292
rect 228646 289356 228882 289442
rect 228646 289292 228732 289356
rect 228732 289292 228796 289356
rect 228796 289292 228882 289356
rect 228646 289206 228882 289292
rect 270414 289206 270650 289442
rect 323038 289206 323274 289442
rect 104446 286086 104682 286322
rect 84574 285126 84810 285362
rect 435862 299606 436098 299842
rect 436182 299606 436418 299842
rect 436502 299606 436738 299842
rect 436822 299606 437058 299842
rect 437142 299606 437378 299842
rect 437462 299606 437698 299842
rect 437782 299606 438018 299842
rect 438102 299606 438338 299842
rect 438422 299606 438658 299842
rect 438742 299606 438978 299842
rect 439062 299606 439298 299842
rect 439382 299606 439618 299842
rect 134806 285126 135042 285362
rect 351742 285126 351978 285362
rect 104506 284288 104742 284524
rect 198506 284288 198742 284524
rect 292506 284288 292742 284524
rect 104446 283326 104682 283562
rect 84390 282406 84626 282642
rect 75006 259286 75242 259522
rect 74086 254526 74322 254762
rect 74270 245686 74506 245922
rect 74086 244326 74322 244562
rect 75926 257926 76162 258162
rect 75374 254526 75610 254762
rect 75374 251806 75610 252042
rect 74822 235636 75058 235722
rect 74822 235572 74908 235636
rect 74908 235572 74972 235636
rect 74972 235572 75058 235636
rect 74822 235486 75058 235572
rect 76846 243646 77082 243882
rect 76478 242286 76714 242522
rect 76478 240926 76714 241162
rect 75926 240246 76162 240482
rect 154494 262686 154730 262922
rect 148974 262006 149210 262242
rect 144006 256566 144242 256802
rect 144006 247726 144242 247962
rect 142902 245686 143138 245922
rect 141062 244326 141298 244562
rect 84390 241076 84626 241162
rect 84390 241012 84476 241076
rect 84476 241012 84540 241076
rect 84540 241012 84626 241076
rect 84390 240926 84626 241012
rect 93774 241076 94010 241162
rect 93774 241012 93860 241076
rect 93860 241012 93924 241076
rect 93924 241012 94010 241076
rect 93774 240926 94010 241012
rect 95982 240926 96218 241162
rect 136830 241606 137066 241842
rect 104814 240246 105050 240482
rect 76846 239566 77082 239802
rect 95062 239716 95298 239802
rect 95062 239652 95148 239716
rect 95148 239652 95212 239716
rect 95212 239652 95298 239716
rect 95062 239566 95298 239652
rect 81262 236846 81498 237082
rect 89910 236996 90146 237082
rect 89910 236932 89996 236996
rect 89996 236932 90060 236996
rect 90060 236932 90146 236996
rect 89910 236846 90146 236932
rect 76294 235486 76530 235722
rect 100030 237526 100266 237762
rect 104998 236166 105234 236402
rect 133886 236166 134122 236402
rect 136278 236166 136514 236402
rect 116038 235486 116274 235722
rect 124318 235636 124554 235722
rect 124318 235572 124404 235636
rect 124404 235572 124468 235636
rect 124468 235572 124554 235636
rect 124318 235486 124554 235572
rect 138302 239566 138538 239802
rect 141062 239566 141298 239802
rect 147686 237526 147922 237762
rect 142902 236846 143138 237082
rect 145110 236846 145346 237082
rect 145846 236846 146082 237082
rect 148606 236846 148842 237082
rect 156702 236166 156938 236402
rect 168110 240246 168346 240482
rect 137198 234956 137434 235042
rect 137198 234892 137284 234956
rect 137284 234892 137348 234956
rect 137348 234892 137434 234956
rect 137198 234806 137434 234892
rect 148054 234956 148290 235042
rect 148054 234892 148140 234956
rect 148140 234892 148204 234956
rect 148204 234892 148290 234956
rect 148054 234806 148290 234892
rect 137566 234276 137802 234362
rect 137566 234212 137652 234276
rect 137652 234212 137716 234276
rect 137716 234212 137802 234276
rect 137566 234126 137802 234212
rect 151918 234126 152154 234362
rect 176942 236846 177178 237082
rect 168846 236166 169082 236402
rect 158726 234806 158962 235042
rect 168478 234806 168714 235042
rect 183750 262156 183986 262242
rect 183750 262092 183836 262156
rect 183836 262092 183900 262156
rect 183900 262092 183986 262156
rect 183750 262006 183986 262092
rect 212454 262006 212690 262242
rect 193134 260646 193370 260882
rect 203070 260796 203306 260882
rect 203070 260732 203156 260796
rect 203156 260732 203220 260796
rect 203220 260732 203306 260796
rect 203070 260646 203306 260732
rect 196078 240396 196314 240482
rect 196078 240332 196164 240396
rect 196164 240332 196228 240396
rect 196228 240332 196314 240396
rect 196078 240246 196314 240332
rect 187798 239716 188034 239802
rect 187798 239652 187884 239716
rect 187884 239652 187948 239716
rect 187948 239652 188034 239716
rect 187798 239566 188034 239652
rect 186510 236996 186746 237082
rect 186510 236932 186596 236996
rect 186596 236932 186660 236996
rect 186660 236932 186746 236996
rect 186510 236846 186746 236932
rect 224782 263366 225018 263602
rect 245022 263516 245258 263602
rect 245022 263452 245108 263516
rect 245108 263452 245172 263516
rect 245172 263452 245258 263516
rect 245022 263366 245258 263452
rect 241342 262006 241578 262242
rect 247782 262006 248018 262242
rect 251094 262006 251330 262242
rect 224782 260646 225018 260882
rect 238030 259286 238266 259522
rect 237662 255206 237898 255442
rect 237662 248406 237898 248642
rect 238030 246366 238266 246602
rect 238030 245686 238266 245922
rect 237662 239566 237898 239802
rect 237662 237526 237898 237762
rect 261950 240246 262186 240482
rect 247046 237526 247282 237762
rect 261582 237526 261818 237762
rect 231774 236846 232010 237082
rect 238030 236846 238266 237082
rect 203070 236316 203306 236402
rect 203070 236252 203156 236316
rect 203156 236252 203220 236316
rect 203220 236252 203306 236316
rect 203070 236166 203306 236252
rect 244102 236180 244338 236402
rect 244102 236166 244188 236180
rect 244188 236166 244252 236180
rect 244252 236166 244338 236180
rect 247046 236166 247282 236402
rect 192030 235486 192266 235722
rect 207118 234806 207354 235042
rect 231222 234956 231458 235042
rect 231222 234892 231308 234956
rect 231308 234892 231372 234956
rect 231372 234892 231458 234956
rect 231222 234806 231458 234892
rect 245390 234956 245626 235042
rect 245390 234892 245476 234956
rect 245476 234892 245540 234956
rect 245540 234892 245626 234956
rect 245390 234806 245626 234892
rect 246126 234806 246362 235042
rect 230670 234140 230906 234362
rect 230670 234126 230756 234140
rect 230756 234126 230820 234140
rect 230820 234126 230906 234140
rect 245390 234126 245626 234362
rect 249806 234126 250042 234362
rect 353582 285276 353818 285362
rect 353582 285212 353668 285276
rect 353668 285212 353732 285276
rect 353732 285212 353818 285276
rect 353582 285126 353818 285212
rect 435862 268970 436098 269206
rect 436182 268970 436418 269206
rect 436502 268970 436738 269206
rect 436822 268970 437058 269206
rect 437142 268970 437378 269206
rect 437462 268970 437698 269206
rect 437782 268970 438018 269206
rect 438102 268970 438338 269206
rect 438422 268970 438658 269206
rect 438742 268970 438978 269206
rect 439062 268970 439298 269206
rect 439382 268970 439618 269206
rect 278878 261476 279114 261562
rect 278878 261412 278964 261476
rect 278964 261412 279028 261476
rect 279028 261412 279114 261476
rect 278878 261326 279114 261412
rect 288446 261476 288682 261562
rect 288446 261412 288532 261476
rect 288532 261412 288596 261476
rect 288596 261412 288682 261476
rect 288446 261326 288682 261412
rect 298198 261476 298434 261562
rect 298198 261412 298284 261476
rect 298284 261412 298348 261476
rect 298348 261412 298434 261476
rect 298198 261326 298434 261412
rect 307766 261476 308002 261562
rect 307766 261412 307852 261476
rect 307852 261412 307916 261476
rect 307916 261412 308002 261476
rect 307766 261326 308002 261412
rect 317518 261476 317754 261562
rect 317518 261412 317604 261476
rect 317604 261412 317668 261476
rect 317668 261412 317754 261476
rect 317518 261326 317754 261412
rect 327086 261476 327322 261562
rect 327086 261412 327172 261476
rect 327172 261412 327236 261476
rect 327236 261412 327322 261476
rect 327086 261326 327322 261412
rect 356158 261326 356394 261562
rect 305006 240396 305242 240482
rect 305006 240332 305092 240396
rect 305092 240332 305156 240396
rect 305156 240332 305242 240396
rect 305006 240246 305242 240332
rect 295438 239788 295524 239802
rect 295524 239788 295588 239802
rect 295588 239788 295674 239802
rect 295438 239566 295674 239788
rect 324510 239716 324746 239802
rect 324510 239652 324596 239716
rect 324596 239652 324660 239716
rect 324660 239652 324746 239716
rect 324510 239566 324746 239652
rect 264710 237526 264946 237762
rect 273726 236996 273962 237082
rect 273726 236932 273812 236996
rect 273812 236932 273876 236996
rect 273876 236932 273962 236996
rect 273726 236846 273962 236932
rect 262318 234806 262554 235042
rect 289918 236846 290154 237082
rect 286790 236316 287026 236402
rect 286790 236252 286876 236316
rect 286876 236252 286940 236316
rect 286940 236252 287026 236316
rect 286790 236166 287026 236252
rect 295438 235486 295674 235722
rect 300958 234956 301194 235042
rect 300958 234892 301044 234956
rect 301044 234892 301108 234956
rect 301108 234892 301194 234956
rect 300958 234806 301194 234892
rect 283110 234348 283196 234362
rect 283196 234348 283260 234362
rect 283260 234348 283346 234362
rect 283110 234126 283346 234348
rect 104506 223016 104742 223252
rect 198506 223016 198742 223252
rect 178598 214406 178834 214642
rect 178598 211006 178834 211242
rect 89146 207698 89382 207934
rect 134622 204900 134858 205122
rect 134622 204886 134708 204900
rect 134708 204886 134772 204900
rect 134772 204886 134858 204900
rect 84574 204428 84660 204442
rect 84660 204428 84724 204442
rect 84724 204428 84810 204442
rect 84574 204206 84810 204428
rect 136830 200956 137066 201042
rect 136830 200892 136916 200956
rect 136916 200892 136980 200956
rect 136980 200892 137066 200956
rect 136830 200806 137066 200892
rect 136830 198766 137066 199002
rect 48878 162726 49114 162962
rect 49062 157966 49298 158202
rect 49062 155396 49298 155482
rect 49062 155332 49148 155396
rect 49148 155332 49212 155396
rect 49212 155332 49298 155396
rect 49062 155246 49298 155332
rect 49062 152526 49298 152762
rect 49062 148446 49298 148682
rect 5122 146426 5358 146662
rect 5442 146426 5678 146662
rect 5762 146426 5998 146662
rect 6082 146426 6318 146662
rect 6402 146426 6638 146662
rect 6722 146426 6958 146662
rect 7042 146426 7278 146662
rect 7362 146426 7598 146662
rect 7682 146426 7918 146662
rect 8002 146426 8238 146662
rect 8322 146426 8558 146662
rect 8642 146426 8878 146662
rect 49062 145876 49298 145962
rect 49062 145812 49148 145876
rect 49148 145812 49212 145876
rect 49212 145812 49298 145876
rect 49062 145726 49298 145812
rect 5122 115790 5358 116026
rect 5442 115790 5678 116026
rect 5762 115790 5998 116026
rect 6082 115790 6318 116026
rect 6402 115790 6638 116026
rect 6722 115790 6958 116026
rect 7042 115790 7278 116026
rect 7362 115790 7598 116026
rect 7682 115790 7918 116026
rect 8002 115790 8238 116026
rect 8322 115790 8558 116026
rect 8642 115790 8878 116026
rect 5122 85154 5358 85390
rect 5442 85154 5678 85390
rect 5762 85154 5998 85390
rect 6082 85154 6318 85390
rect 6402 85154 6638 85390
rect 6722 85154 6958 85390
rect 7042 85154 7278 85390
rect 7362 85154 7598 85390
rect 7682 85154 7918 85390
rect 8002 85154 8238 85390
rect 8322 85154 8558 85390
rect 8642 85154 8878 85390
rect 137934 194006 138170 194242
rect 104506 192380 104742 192616
rect 176574 198086 176810 198322
rect 164430 197406 164666 197642
rect 183146 207698 183382 207934
rect 292506 223016 292742 223252
rect 322670 217806 322906 218042
rect 242630 216596 242866 216682
rect 242630 216532 242716 216596
rect 242716 216532 242780 216596
rect 242780 216532 242866 216596
rect 242630 216446 242866 216532
rect 258822 216596 259058 216682
rect 258822 216532 258908 216596
rect 258908 216532 258972 216596
rect 258972 216532 259058 216596
rect 258822 216446 259058 216532
rect 272622 216596 272858 216682
rect 272622 216532 272708 216596
rect 272708 216532 272772 216596
rect 272772 216532 272858 216596
rect 272622 216446 272858 216532
rect 336654 216596 336890 216682
rect 336654 216532 336740 216596
rect 336740 216532 336804 216596
rect 336804 216532 336890 216596
rect 336654 216446 336890 216532
rect 277146 207698 277382 207934
rect 239502 204356 239738 204442
rect 239502 204292 239588 204356
rect 239588 204292 239652 204356
rect 239652 204292 239738 204356
rect 228646 200956 228882 201042
rect 228646 200892 228732 200956
rect 228732 200892 228796 200956
rect 228796 200892 228882 200956
rect 228646 200806 228882 200892
rect 230670 198766 230906 199002
rect 178598 195366 178834 195602
rect 178598 194686 178834 194922
rect 230670 194006 230906 194242
rect 198506 192380 198742 192616
rect 178598 185846 178834 186082
rect 178230 182446 178466 182682
rect 75374 164766 75610 165002
rect 74086 156606 74322 156842
rect 75374 160006 75610 160242
rect 75190 157966 75426 158202
rect 75374 156606 75610 156842
rect 74270 152526 74506 152762
rect 76662 164766 76898 165002
rect 76662 162726 76898 162962
rect 144006 160686 144242 160922
rect 76662 160006 76898 160242
rect 76294 156606 76530 156842
rect 76662 154566 76898 154802
rect 77030 153206 77266 153442
rect 74638 148446 74874 148682
rect 74454 145726 74690 145962
rect 74822 145046 75058 145282
rect 74822 143686 75058 143922
rect 76478 145876 76714 145962
rect 76478 145812 76564 145876
rect 76564 145812 76628 145876
rect 76628 145812 76714 145876
rect 76478 145726 76714 145812
rect 144006 150486 144242 150722
rect 77030 145046 77266 145282
rect 142350 144366 142586 144602
rect 75926 143006 76162 143242
rect 98190 143686 98426 143922
rect 110334 143228 110420 143242
rect 110420 143228 110484 143242
rect 110484 143228 110570 143242
rect 110334 143006 110570 143228
rect 136830 143228 136916 143242
rect 136916 143228 136980 143242
rect 136980 143228 137066 143242
rect 136830 143006 137066 143228
rect 78134 141796 78370 141882
rect 78134 141732 78220 141796
rect 78220 141732 78284 141796
rect 78284 141732 78370 141796
rect 78134 141646 78370 141732
rect 151734 143006 151970 143242
rect 104998 141868 105084 141882
rect 105084 141868 105148 141882
rect 105148 141868 105234 141882
rect 104998 141646 105234 141868
rect 168294 141796 168530 141882
rect 168294 141732 168380 141796
rect 168380 141732 168444 141796
rect 168444 141732 168530 141796
rect 168294 141646 168530 141732
rect 137382 141116 137618 141202
rect 137382 141052 137468 141116
rect 137468 141052 137532 141116
rect 137532 141052 137618 141116
rect 137382 140966 137618 141052
rect 148974 141116 149210 141202
rect 148974 141052 149060 141116
rect 149060 141052 149124 141116
rect 149124 141052 149210 141116
rect 148974 140966 149210 141052
rect 168478 140966 168714 141202
rect 174734 179726 174970 179962
rect 228830 181086 229066 181322
rect 169398 145046 169634 145282
rect 176206 145196 176442 145282
rect 176206 145132 176292 145196
rect 176292 145132 176356 145196
rect 176356 145132 176442 145196
rect 176206 145046 176442 145132
rect 169398 143006 169634 143242
rect 170134 143006 170370 143242
rect 137198 140300 137434 140522
rect 137198 140286 137284 140300
rect 137284 140286 137348 140300
rect 137348 140286 137434 140300
rect 151918 140436 152154 140522
rect 151918 140372 152004 140436
rect 152004 140372 152068 140436
rect 152068 140372 152154 140436
rect 151918 140286 152154 140372
rect 136830 116636 137066 116722
rect 136830 116572 136916 116636
rect 136916 116572 136980 116636
rect 136980 116572 137066 116636
rect 136830 116486 137066 116572
rect 89146 115790 89382 116026
rect 146582 113236 146818 113322
rect 187062 144366 187298 144602
rect 196078 144516 196314 144602
rect 196078 144452 196164 144516
rect 196164 144452 196228 144516
rect 196228 144452 196314 144516
rect 196078 144366 196314 144452
rect 210062 143156 210298 143242
rect 210062 143092 210148 143156
rect 210148 143092 210212 143156
rect 210212 143092 210298 143156
rect 210062 143006 210298 143092
rect 239502 204206 239738 204292
rect 322670 204220 322906 204442
rect 322670 204206 322756 204220
rect 322756 204206 322820 204220
rect 322820 204206 322906 204220
rect 322670 200956 322906 201042
rect 322670 200892 322756 200956
rect 322756 200892 322820 200956
rect 322820 200892 322906 200956
rect 322670 200806 322906 200892
rect 322670 198780 322906 199002
rect 322670 198766 322756 198780
rect 322756 198766 322820 198780
rect 322820 198766 322906 198780
rect 270414 198086 270650 198322
rect 261030 197556 261266 197642
rect 261030 197492 261116 197556
rect 261116 197492 261180 197556
rect 261180 197492 261266 197556
rect 261030 197406 261266 197492
rect 322670 194006 322906 194242
rect 292506 192380 292742 192616
rect 352662 216596 352898 216682
rect 352662 216532 352748 216596
rect 352748 216532 352812 216596
rect 352812 216532 352898 216596
rect 352662 216446 352898 216532
rect 435862 238334 436098 238570
rect 436182 238334 436418 238570
rect 436502 238334 436738 238570
rect 436822 238334 437058 238570
rect 437142 238334 437378 238570
rect 437462 238334 437698 238570
rect 437782 238334 438018 238570
rect 438102 238334 438338 238570
rect 438422 238334 438658 238570
rect 438742 238334 438978 238570
rect 439062 238334 439298 238570
rect 439382 238334 439618 238570
rect 380882 223016 381118 223252
rect 357446 215916 357682 216002
rect 357446 215852 357532 215916
rect 357532 215852 357596 215916
rect 357596 215852 357682 215916
rect 357446 215766 357682 215852
rect 405838 215916 406074 216002
rect 405838 215852 405924 215916
rect 405924 215852 405988 215916
rect 405988 215852 406074 215916
rect 405838 215766 406074 215852
rect 435862 207698 436098 207934
rect 436182 207698 436418 207934
rect 436502 207698 436738 207934
rect 436822 207698 437058 207934
rect 437142 207698 437378 207934
rect 437462 207698 437698 207934
rect 437782 207698 438018 207934
rect 438102 207698 438338 207934
rect 438422 207698 438658 207934
rect 438742 207698 438978 207934
rect 439062 207698 439298 207934
rect 439382 207698 439618 207934
rect 322854 183126 323090 183362
rect 271334 182446 271570 182682
rect 322854 181988 322940 182002
rect 322940 181988 323004 182002
rect 323004 181988 323090 182002
rect 241710 168846 241946 169082
rect 242262 168166 242498 168402
rect 243182 168166 243418 168402
rect 238030 165446 238266 165682
rect 237662 164766 237898 165002
rect 237294 164086 237530 164322
rect 237294 160686 237530 160922
rect 238030 157286 238266 157522
rect 237662 156606 237898 156842
rect 236742 153206 236978 153442
rect 237294 148446 237530 148682
rect 237478 147086 237714 147322
rect 207118 141116 207354 141202
rect 207118 141052 207204 141116
rect 207204 141052 207268 141116
rect 207268 141052 207354 141116
rect 207118 140966 207354 141052
rect 236006 141646 236242 141882
rect 237662 141796 237898 141882
rect 237662 141732 237748 141796
rect 237748 141732 237812 141796
rect 237812 141732 237898 141796
rect 237662 141646 237898 141732
rect 230670 140286 230906 140522
rect 199206 130766 199442 131002
rect 256614 141796 256850 141882
rect 256614 141732 256700 141796
rect 256700 141732 256764 141796
rect 256764 141732 256850 141796
rect 256614 141646 256850 141732
rect 322854 181766 323090 181988
rect 271334 179726 271570 179962
rect 286054 179196 286290 179282
rect 286054 179132 286140 179196
rect 286140 179132 286204 179196
rect 286204 179132 286290 179196
rect 286054 179046 286290 179132
rect 287342 179268 287428 179282
rect 287428 179268 287492 179282
rect 287492 179268 287578 179282
rect 287342 179046 287578 179268
rect 288446 179196 288682 179282
rect 288446 179132 288532 179196
rect 288532 179132 288596 179196
rect 288596 179132 288682 179196
rect 288446 179046 288682 179132
rect 289366 179268 289452 179282
rect 289452 179268 289516 179282
rect 289516 179268 289602 179282
rect 289366 179046 289602 179268
rect 309790 179196 310026 179282
rect 309790 179132 309876 179196
rect 309876 179132 309940 179196
rect 309940 179132 310026 179196
rect 309790 179046 310026 179132
rect 310894 179268 310980 179282
rect 310980 179268 311044 179282
rect 311044 179268 311130 179282
rect 310894 179046 311130 179268
rect 311814 179196 312050 179282
rect 311814 179132 311900 179196
rect 311900 179132 311964 179196
rect 311964 179132 312050 179196
rect 311814 179046 312050 179132
rect 316966 179268 317052 179282
rect 317052 179268 317116 179282
rect 317116 179268 317202 179282
rect 316966 179046 317202 179268
rect 435862 177062 436098 177298
rect 436182 177062 436418 177298
rect 436502 177062 436738 177298
rect 436822 177062 437058 177298
rect 437142 177062 437378 177298
rect 437462 177062 437698 177298
rect 437782 177062 438018 177298
rect 438102 177062 438338 177298
rect 438422 177062 438658 177298
rect 438742 177062 438978 177298
rect 439062 177062 439298 177298
rect 439382 177062 439618 177298
rect 435862 146426 436098 146662
rect 436182 146426 436418 146662
rect 436502 146426 436738 146662
rect 436822 146426 437058 146662
rect 437142 146426 437378 146662
rect 437462 146426 437698 146662
rect 437782 146426 438018 146662
rect 438102 146426 438338 146662
rect 438422 146426 438658 146662
rect 438742 146426 438978 146662
rect 439062 146426 439298 146662
rect 439382 146426 439618 146662
rect 262870 143006 263106 143242
rect 262318 140966 262554 141202
rect 242998 140286 243234 140522
rect 251278 140286 251514 140522
rect 294150 143156 294386 143242
rect 294150 143092 294236 143156
rect 294236 143092 294300 143156
rect 294300 143092 294386 143156
rect 294150 143006 294386 143092
rect 289918 141646 290154 141882
rect 296910 141116 297146 141202
rect 296910 141052 296996 141116
rect 296996 141052 297060 141116
rect 297060 141052 297146 141116
rect 296910 140966 297146 141052
rect 178598 124646 178834 124882
rect 178598 123966 178834 124202
rect 163694 117846 163930 118082
rect 148422 117166 148658 117402
rect 163694 115126 163930 115362
rect 163694 114446 163930 114682
rect 152102 113766 152338 114002
rect 146582 113172 146668 113236
rect 146668 113172 146732 113236
rect 146732 113172 146818 113236
rect 146582 113086 146818 113172
rect 84574 109836 84810 109922
rect 84574 109772 84660 109836
rect 84660 109772 84724 109836
rect 84724 109772 84810 109836
rect 84574 109686 84810 109772
rect 134622 109836 134858 109922
rect 134622 109772 134708 109836
rect 134708 109772 134772 109836
rect 134772 109772 134858 109836
rect 134622 109686 134858 109772
rect 137934 104396 138170 104482
rect 137934 104332 138020 104396
rect 138020 104332 138084 104396
rect 138084 104332 138170 104396
rect 137934 104246 138170 104332
rect 137382 101526 137618 101762
rect 104506 100472 104742 100708
rect 145662 99486 145898 99722
rect 74454 93366 74690 93602
rect 84574 93516 84810 93602
rect 84574 93452 84660 93516
rect 84660 93452 84724 93516
rect 84724 93452 84810 93516
rect 84574 93366 84810 93452
rect 245758 123966 245994 124202
rect 245390 123286 245626 123522
rect 231774 119356 232010 119442
rect 231774 119292 231860 119356
rect 231860 119292 231924 119356
rect 231924 119292 232010 119356
rect 231774 119206 232010 119292
rect 242078 119206 242314 119442
rect 229198 117846 229434 118082
rect 238766 116636 239002 116722
rect 238766 116572 238852 116636
rect 238852 116572 238916 116636
rect 238916 116572 239002 116636
rect 238766 116486 239002 116572
rect 183146 115790 183382 116026
rect 230670 112406 230906 112642
rect 245390 116486 245626 116722
rect 240054 109836 240290 109922
rect 240054 109772 240140 109836
rect 240140 109772 240204 109836
rect 240204 109772 240290 109836
rect 240054 109686 240290 109772
rect 178598 108326 178834 108562
rect 177862 106966 178098 107202
rect 163694 105606 163930 105842
rect 163694 104926 163930 105162
rect 164798 104246 165034 104482
rect 176942 102886 177178 103122
rect 171238 101526 171474 101762
rect 164798 98126 165034 98362
rect 178598 103566 178834 103802
rect 229014 102206 229250 102442
rect 231774 104396 232010 104482
rect 231774 104332 231860 104396
rect 231860 104332 231924 104396
rect 231924 104332 232010 104396
rect 231774 104246 232010 104332
rect 230670 101526 230906 101762
rect 245758 113766 245994 114002
rect 245390 104926 245626 105162
rect 245390 103566 245626 103802
rect 198506 100472 198742 100708
rect 178598 98806 178834 99042
rect 242630 99486 242866 99722
rect 228646 98126 228882 98362
rect 177862 96086 178098 96322
rect 245390 96086 245626 96322
rect 163694 94046 163930 94282
rect 155230 90646 155466 90882
rect 178598 88606 178834 88842
rect 5122 54518 5358 54754
rect 5442 54518 5678 54754
rect 5762 54518 5998 54754
rect 6082 54518 6318 54754
rect 6402 54518 6638 54754
rect 6722 54518 6958 54754
rect 7042 54518 7278 54754
rect 7362 54518 7598 54754
rect 7682 54518 7918 54754
rect 8002 54518 8238 54754
rect 8322 54518 8558 54754
rect 8642 54518 8878 54754
rect 67830 48486 68066 48722
rect 73166 48486 73402 48722
rect 148422 73646 148658 73882
rect 155966 73646 156202 73882
rect 144558 72966 144794 73202
rect 144558 64126 144794 64362
rect 144742 63446 144978 63682
rect 102422 51356 102658 51442
rect 102422 51292 102508 51356
rect 102508 51292 102572 51356
rect 102572 51292 102658 51356
rect 102422 51206 102658 51292
rect 93590 50676 93826 50762
rect 93590 50612 93676 50676
rect 93676 50612 93740 50676
rect 93740 50612 93826 50676
rect 93590 50526 93826 50612
rect 74454 49166 74690 49402
rect 88254 49316 88490 49402
rect 88254 49252 88340 49316
rect 88340 49252 88404 49316
rect 88404 49252 88490 49316
rect 88254 49166 88490 49252
rect 105182 49316 105418 49402
rect 105182 49252 105268 49316
rect 105268 49252 105332 49316
rect 105332 49252 105418 49316
rect 105182 49166 105418 49252
rect 88070 48636 88306 48722
rect 88070 48572 88156 48636
rect 88156 48572 88220 48636
rect 88220 48572 88306 48636
rect 88070 48486 88306 48572
rect 110334 47276 110570 47362
rect 110334 47212 110420 47276
rect 110420 47212 110484 47276
rect 110484 47212 110570 47276
rect 110334 47126 110570 47212
rect 107390 46446 107626 46682
rect 142350 51206 142586 51442
rect 145478 49166 145714 49402
rect 147870 49166 148106 49402
rect 167926 49166 168162 49402
rect 154678 48486 154914 48722
rect 167558 48486 167794 48722
rect 160014 47956 160250 48042
rect 160014 47892 160100 47956
rect 160100 47892 160164 47956
rect 160164 47892 160250 47956
rect 160014 47806 160250 47892
rect 249070 127366 249306 127602
rect 248518 126836 248754 126922
rect 248518 126772 248604 126836
rect 248604 126772 248668 126836
rect 248668 126772 248754 126836
rect 248518 126686 248754 126772
rect 258638 103566 258874 103802
rect 258638 99486 258874 99722
rect 249438 89966 249674 90202
rect 249438 88828 249524 88842
rect 249524 88828 249588 88842
rect 249588 88828 249674 88842
rect 249438 88606 249674 88828
rect 277146 115790 277382 116026
rect 322670 109836 322906 109922
rect 322670 109772 322756 109836
rect 322756 109772 322820 109836
rect 322820 109772 322906 109836
rect 322670 109686 322906 109772
rect 261030 103036 261266 103122
rect 261030 102972 261116 103036
rect 261116 102972 261180 103036
rect 261180 102972 261266 103036
rect 261030 102886 261266 102972
rect 272622 102206 272858 102442
rect 323038 102206 323274 102442
rect 270414 101526 270650 101762
rect 324510 101526 324746 101762
rect 292506 100472 292742 100708
rect 272622 99486 272858 99722
rect 322670 98126 322906 98362
rect 435862 115790 436098 116026
rect 436182 115790 436418 116026
rect 436502 115790 436738 116026
rect 436822 115790 437058 116026
rect 437142 115790 437378 116026
rect 437462 115790 437698 116026
rect 437782 115790 438018 116026
rect 438102 115790 438338 116026
rect 438422 115790 438658 116026
rect 438742 115790 438978 116026
rect 439062 115790 439298 116026
rect 439382 115790 439618 116026
rect 263790 88606 264026 88842
rect 251646 87926 251882 88162
rect 259558 87926 259794 88162
rect 261582 87926 261818 88162
rect 169950 73646 170186 73882
rect 249806 73646 250042 73882
rect 238582 60046 238818 60282
rect 237294 59366 237530 59602
rect 187062 50676 187298 50762
rect 187062 50612 187148 50676
rect 187148 50612 187212 50676
rect 187212 50612 187298 50676
rect 187062 50526 187298 50612
rect 181910 49316 182146 49402
rect 181910 49252 181996 49316
rect 181996 49252 182060 49316
rect 182060 49252 182146 49316
rect 181910 49166 182146 49252
rect 169030 47806 169266 48042
rect 158910 47126 159146 47362
rect 157438 46446 157674 46682
rect 162774 46596 163010 46682
rect 162774 46532 162860 46596
rect 162860 46532 162924 46596
rect 162924 46532 163010 46596
rect 162774 46446 163010 46532
rect 191294 48486 191530 48722
rect 181726 47956 181962 48042
rect 181726 47892 181812 47956
rect 181812 47892 181876 47956
rect 181876 47892 181962 47956
rect 181726 47806 181962 47892
rect 181726 46668 181812 46682
rect 181812 46668 181876 46682
rect 181876 46668 181962 46682
rect 181726 46446 181962 46668
rect 204174 46446 204410 46682
rect 238582 51206 238818 51442
rect 237662 50526 237898 50762
rect 248886 48486 249122 48722
rect 248518 47276 248754 47362
rect 248518 47212 248604 47276
rect 248604 47212 248668 47276
rect 248668 47212 248754 47276
rect 248518 47126 248754 47212
rect 250358 47956 250594 48042
rect 250358 47892 250444 47956
rect 250444 47892 250508 47956
rect 250508 47892 250594 47956
rect 250358 47806 250594 47892
rect 261030 47956 261266 48042
rect 261030 47892 261116 47956
rect 261116 47892 261180 47956
rect 261180 47892 261266 47956
rect 261030 47806 261266 47892
rect 252750 46446 252986 46682
rect 261766 46446 262002 46682
rect 264158 73646 264394 73882
rect 270598 51886 270834 52122
rect 264158 48486 264394 48722
rect 275934 47956 276170 48042
rect 275934 47892 276020 47956
rect 276020 47892 276084 47956
rect 276084 47892 276170 47956
rect 275934 47806 276170 47892
rect 263790 47348 263876 47362
rect 263876 47348 263940 47362
rect 263940 47348 264026 47362
rect 263790 47126 264026 47348
rect 275750 46596 275986 46682
rect 275750 46532 275836 46596
rect 275836 46532 275900 46596
rect 275900 46532 275986 46596
rect 275750 46446 275986 46532
rect 435862 85154 436098 85390
rect 436182 85154 436418 85390
rect 436502 85154 436738 85390
rect 436822 85154 437058 85390
rect 437142 85154 437378 85390
rect 437462 85154 437698 85390
rect 437782 85154 438018 85390
rect 438102 85154 438338 85390
rect 438422 85154 438658 85390
rect 438742 85154 438978 85390
rect 439062 85154 439298 85390
rect 439382 85154 439618 85390
rect 435862 54518 436098 54754
rect 436182 54518 436418 54754
rect 436502 54518 436738 54754
rect 436822 54518 437058 54754
rect 437142 54518 437378 54754
rect 437462 54518 437698 54754
rect 437782 54518 438018 54754
rect 438102 54518 438338 54754
rect 438422 54518 438658 54754
rect 438742 54518 438978 54754
rect 439062 54518 439298 54754
rect 439382 54518 439618 54754
rect 5122 23882 5358 24118
rect 5442 23882 5678 24118
rect 5762 23882 5998 24118
rect 6082 23882 6318 24118
rect 6402 23882 6638 24118
rect 6722 23882 6958 24118
rect 7042 23882 7278 24118
rect 7362 23882 7598 24118
rect 7682 23882 7918 24118
rect 8002 23882 8238 24118
rect 8322 23882 8558 24118
rect 8642 23882 8878 24118
rect 5122 8642 5358 8878
rect 5442 8642 5678 8878
rect 5762 8642 5998 8878
rect 6082 8642 6318 8878
rect 6402 8642 6638 8878
rect 6722 8642 6958 8878
rect 7042 8642 7278 8878
rect 7362 8642 7598 8878
rect 7682 8642 7918 8878
rect 8002 8642 8238 8878
rect 8322 8642 8558 8878
rect 8642 8642 8878 8878
rect 5122 8322 5358 8558
rect 5442 8322 5678 8558
rect 5762 8322 5998 8558
rect 6082 8322 6318 8558
rect 6402 8322 6638 8558
rect 6722 8322 6958 8558
rect 7042 8322 7278 8558
rect 7362 8322 7598 8558
rect 7682 8322 7918 8558
rect 8002 8322 8238 8558
rect 8322 8322 8558 8558
rect 8642 8322 8878 8558
rect 5122 8002 5358 8238
rect 5442 8002 5678 8238
rect 5762 8002 5998 8238
rect 6082 8002 6318 8238
rect 6402 8002 6638 8238
rect 6722 8002 6958 8238
rect 7042 8002 7278 8238
rect 7362 8002 7598 8238
rect 7682 8002 7918 8238
rect 8002 8002 8238 8238
rect 8322 8002 8558 8238
rect 8642 8002 8878 8238
rect 5122 7682 5358 7918
rect 5442 7682 5678 7918
rect 5762 7682 5998 7918
rect 6082 7682 6318 7918
rect 6402 7682 6638 7918
rect 6722 7682 6958 7918
rect 7042 7682 7278 7918
rect 7362 7682 7598 7918
rect 7682 7682 7918 7918
rect 8002 7682 8238 7918
rect 8322 7682 8558 7918
rect 8642 7682 8878 7918
rect 5122 7362 5358 7598
rect 5442 7362 5678 7598
rect 5762 7362 5998 7598
rect 6082 7362 6318 7598
rect 6402 7362 6638 7598
rect 6722 7362 6958 7598
rect 7042 7362 7278 7598
rect 7362 7362 7598 7598
rect 7682 7362 7918 7598
rect 8002 7362 8238 7598
rect 8322 7362 8558 7598
rect 8642 7362 8878 7598
rect 5122 7042 5358 7278
rect 5442 7042 5678 7278
rect 5762 7042 5998 7278
rect 6082 7042 6318 7278
rect 6402 7042 6638 7278
rect 6722 7042 6958 7278
rect 7042 7042 7278 7278
rect 7362 7042 7598 7278
rect 7682 7042 7918 7278
rect 8002 7042 8238 7278
rect 8322 7042 8558 7278
rect 8642 7042 8878 7278
rect 5122 6722 5358 6958
rect 5442 6722 5678 6958
rect 5762 6722 5998 6958
rect 6082 6722 6318 6958
rect 6402 6722 6638 6958
rect 6722 6722 6958 6958
rect 7042 6722 7278 6958
rect 7362 6722 7598 6958
rect 7682 6722 7918 6958
rect 8002 6722 8238 6958
rect 8322 6722 8558 6958
rect 8642 6722 8878 6958
rect 5122 6402 5358 6638
rect 5442 6402 5678 6638
rect 5762 6402 5998 6638
rect 6082 6402 6318 6638
rect 6402 6402 6638 6638
rect 6722 6402 6958 6638
rect 7042 6402 7278 6638
rect 7362 6402 7598 6638
rect 7682 6402 7918 6638
rect 8002 6402 8238 6638
rect 8322 6402 8558 6638
rect 8642 6402 8878 6638
rect 5122 6082 5358 6318
rect 5442 6082 5678 6318
rect 5762 6082 5998 6318
rect 6082 6082 6318 6318
rect 6402 6082 6638 6318
rect 6722 6082 6958 6318
rect 7042 6082 7278 6318
rect 7362 6082 7598 6318
rect 7682 6082 7918 6318
rect 8002 6082 8238 6318
rect 8322 6082 8558 6318
rect 8642 6082 8878 6318
rect 5122 5762 5358 5998
rect 5442 5762 5678 5998
rect 5762 5762 5998 5998
rect 6082 5762 6318 5998
rect 6402 5762 6638 5998
rect 6722 5762 6958 5998
rect 7042 5762 7278 5998
rect 7362 5762 7598 5998
rect 7682 5762 7918 5998
rect 8002 5762 8238 5998
rect 8322 5762 8558 5998
rect 8642 5762 8878 5998
rect 5122 5442 5358 5678
rect 5442 5442 5678 5678
rect 5762 5442 5998 5678
rect 6082 5442 6318 5678
rect 6402 5442 6638 5678
rect 6722 5442 6958 5678
rect 7042 5442 7278 5678
rect 7362 5442 7598 5678
rect 7682 5442 7918 5678
rect 8002 5442 8238 5678
rect 8322 5442 8558 5678
rect 8642 5442 8878 5678
rect 5122 5122 5358 5358
rect 5442 5122 5678 5358
rect 5762 5122 5998 5358
rect 6082 5122 6318 5358
rect 6402 5122 6638 5358
rect 6722 5122 6958 5358
rect 7042 5122 7278 5358
rect 7362 5122 7598 5358
rect 7682 5122 7918 5358
rect 8002 5122 8238 5358
rect 8322 5122 8558 5358
rect 8642 5122 8878 5358
rect 435862 23882 436098 24118
rect 436182 23882 436418 24118
rect 436502 23882 436738 24118
rect 436822 23882 437058 24118
rect 437142 23882 437378 24118
rect 437462 23882 437698 24118
rect 437782 23882 438018 24118
rect 438102 23882 438338 24118
rect 438422 23882 438658 24118
rect 438742 23882 438978 24118
rect 439062 23882 439298 24118
rect 439382 23882 439618 24118
rect 435862 8642 436098 8878
rect 436182 8642 436418 8878
rect 436502 8642 436738 8878
rect 436822 8642 437058 8878
rect 437142 8642 437378 8878
rect 437462 8642 437698 8878
rect 437782 8642 438018 8878
rect 438102 8642 438338 8878
rect 438422 8642 438658 8878
rect 438742 8642 438978 8878
rect 439062 8642 439298 8878
rect 439382 8642 439618 8878
rect 435862 8322 436098 8558
rect 436182 8322 436418 8558
rect 436502 8322 436738 8558
rect 436822 8322 437058 8558
rect 437142 8322 437378 8558
rect 437462 8322 437698 8558
rect 437782 8322 438018 8558
rect 438102 8322 438338 8558
rect 438422 8322 438658 8558
rect 438742 8322 438978 8558
rect 439062 8322 439298 8558
rect 439382 8322 439618 8558
rect 435862 8002 436098 8238
rect 436182 8002 436418 8238
rect 436502 8002 436738 8238
rect 436822 8002 437058 8238
rect 437142 8002 437378 8238
rect 437462 8002 437698 8238
rect 437782 8002 438018 8238
rect 438102 8002 438338 8238
rect 438422 8002 438658 8238
rect 438742 8002 438978 8238
rect 439062 8002 439298 8238
rect 439382 8002 439618 8238
rect 435862 7682 436098 7918
rect 436182 7682 436418 7918
rect 436502 7682 436738 7918
rect 436822 7682 437058 7918
rect 437142 7682 437378 7918
rect 437462 7682 437698 7918
rect 437782 7682 438018 7918
rect 438102 7682 438338 7918
rect 438422 7682 438658 7918
rect 438742 7682 438978 7918
rect 439062 7682 439298 7918
rect 439382 7682 439618 7918
rect 435862 7362 436098 7598
rect 436182 7362 436418 7598
rect 436502 7362 436738 7598
rect 436822 7362 437058 7598
rect 437142 7362 437378 7598
rect 437462 7362 437698 7598
rect 437782 7362 438018 7598
rect 438102 7362 438338 7598
rect 438422 7362 438658 7598
rect 438742 7362 438978 7598
rect 439062 7362 439298 7598
rect 439382 7362 439618 7598
rect 435862 7042 436098 7278
rect 436182 7042 436418 7278
rect 436502 7042 436738 7278
rect 436822 7042 437058 7278
rect 437142 7042 437378 7278
rect 437462 7042 437698 7278
rect 437782 7042 438018 7278
rect 438102 7042 438338 7278
rect 438422 7042 438658 7278
rect 438742 7042 438978 7278
rect 439062 7042 439298 7278
rect 439382 7042 439618 7278
rect 435862 6722 436098 6958
rect 436182 6722 436418 6958
rect 436502 6722 436738 6958
rect 436822 6722 437058 6958
rect 437142 6722 437378 6958
rect 437462 6722 437698 6958
rect 437782 6722 438018 6958
rect 438102 6722 438338 6958
rect 438422 6722 438658 6958
rect 438742 6722 438978 6958
rect 439062 6722 439298 6958
rect 439382 6722 439618 6958
rect 435862 6402 436098 6638
rect 436182 6402 436418 6638
rect 436502 6402 436738 6638
rect 436822 6402 437058 6638
rect 437142 6402 437378 6638
rect 437462 6402 437698 6638
rect 437782 6402 438018 6638
rect 438102 6402 438338 6638
rect 438422 6402 438658 6638
rect 438742 6402 438978 6638
rect 439062 6402 439298 6638
rect 439382 6402 439618 6638
rect 435862 6082 436098 6318
rect 436182 6082 436418 6318
rect 436502 6082 436738 6318
rect 436822 6082 437058 6318
rect 437142 6082 437378 6318
rect 437462 6082 437698 6318
rect 437782 6082 438018 6318
rect 438102 6082 438338 6318
rect 438422 6082 438658 6318
rect 438742 6082 438978 6318
rect 439062 6082 439298 6318
rect 439382 6082 439618 6318
rect 435862 5762 436098 5998
rect 436182 5762 436418 5998
rect 436502 5762 436738 5998
rect 436822 5762 437058 5998
rect 437142 5762 437378 5998
rect 437462 5762 437698 5998
rect 437782 5762 438018 5998
rect 438102 5762 438338 5998
rect 438422 5762 438658 5998
rect 438742 5762 438978 5998
rect 439062 5762 439298 5998
rect 439382 5762 439618 5998
rect 435862 5442 436098 5678
rect 436182 5442 436418 5678
rect 436502 5442 436738 5678
rect 436822 5442 437058 5678
rect 437142 5442 437378 5678
rect 437462 5442 437698 5678
rect 437782 5442 438018 5678
rect 438102 5442 438338 5678
rect 438422 5442 438658 5678
rect 438742 5442 438978 5678
rect 439062 5442 439298 5678
rect 439382 5442 439618 5678
rect 435862 5122 436098 5358
rect 436182 5122 436418 5358
rect 436502 5122 436738 5358
rect 436822 5122 437058 5358
rect 437142 5122 437378 5358
rect 437462 5122 437698 5358
rect 437782 5122 438018 5358
rect 438102 5122 438338 5358
rect 438422 5122 438658 5358
rect 438742 5122 438978 5358
rect 439062 5122 439298 5358
rect 439382 5122 439618 5358
rect 440862 376196 441098 376432
rect 441182 376196 441418 376432
rect 441502 376196 441738 376432
rect 441822 376196 442058 376432
rect 442142 376196 442378 376432
rect 442462 376196 442698 376432
rect 442782 376196 443018 376432
rect 443102 376196 443338 376432
rect 443422 376196 443658 376432
rect 443742 376196 443978 376432
rect 444062 376196 444298 376432
rect 444382 376196 444618 376432
rect 440862 345560 441098 345796
rect 441182 345560 441418 345796
rect 441502 345560 441738 345796
rect 441822 345560 442058 345796
rect 442142 345560 442378 345796
rect 442462 345560 442698 345796
rect 442782 345560 443018 345796
rect 443102 345560 443338 345796
rect 443422 345560 443658 345796
rect 443742 345560 443978 345796
rect 444062 345560 444298 345796
rect 444382 345560 444618 345796
rect 440862 314924 441098 315160
rect 441182 314924 441418 315160
rect 441502 314924 441738 315160
rect 441822 314924 442058 315160
rect 442142 314924 442378 315160
rect 442462 314924 442698 315160
rect 442782 314924 443018 315160
rect 443102 314924 443338 315160
rect 443422 314924 443658 315160
rect 443742 314924 443978 315160
rect 444062 314924 444298 315160
rect 444382 314924 444618 315160
rect 440862 284288 441098 284524
rect 441182 284288 441418 284524
rect 441502 284288 441738 284524
rect 441822 284288 442058 284524
rect 442142 284288 442378 284524
rect 442462 284288 442698 284524
rect 442782 284288 443018 284524
rect 443102 284288 443338 284524
rect 443422 284288 443658 284524
rect 443742 284288 443978 284524
rect 444062 284288 444298 284524
rect 444382 284288 444618 284524
rect 440862 253652 441098 253888
rect 441182 253652 441418 253888
rect 441502 253652 441738 253888
rect 441822 253652 442058 253888
rect 442142 253652 442378 253888
rect 442462 253652 442698 253888
rect 442782 253652 443018 253888
rect 443102 253652 443338 253888
rect 443422 253652 443658 253888
rect 443742 253652 443978 253888
rect 444062 253652 444298 253888
rect 444382 253652 444618 253888
rect 440862 223016 441098 223252
rect 441182 223016 441418 223252
rect 441502 223016 441738 223252
rect 441822 223016 442058 223252
rect 442142 223016 442378 223252
rect 442462 223016 442698 223252
rect 442782 223016 443018 223252
rect 443102 223016 443338 223252
rect 443422 223016 443658 223252
rect 443742 223016 443978 223252
rect 444062 223016 444298 223252
rect 444382 223016 444618 223252
rect 440862 192380 441098 192616
rect 441182 192380 441418 192616
rect 441502 192380 441738 192616
rect 441822 192380 442058 192616
rect 442142 192380 442378 192616
rect 442462 192380 442698 192616
rect 442782 192380 443018 192616
rect 443102 192380 443338 192616
rect 443422 192380 443658 192616
rect 443742 192380 443978 192616
rect 444062 192380 444298 192616
rect 444382 192380 444618 192616
rect 440862 161744 441098 161980
rect 441182 161744 441418 161980
rect 441502 161744 441738 161980
rect 441822 161744 442058 161980
rect 442142 161744 442378 161980
rect 442462 161744 442698 161980
rect 442782 161744 443018 161980
rect 443102 161744 443338 161980
rect 443422 161744 443658 161980
rect 443742 161744 443978 161980
rect 444062 161744 444298 161980
rect 444382 161744 444618 161980
rect 440862 131108 441098 131344
rect 441182 131108 441418 131344
rect 441502 131108 441738 131344
rect 441822 131108 442058 131344
rect 442142 131108 442378 131344
rect 442462 131108 442698 131344
rect 442782 131108 443018 131344
rect 443102 131108 443338 131344
rect 443422 131108 443658 131344
rect 443742 131108 443978 131344
rect 444062 131108 444298 131344
rect 444382 131108 444618 131344
rect 440862 100472 441098 100708
rect 441182 100472 441418 100708
rect 441502 100472 441738 100708
rect 441822 100472 442058 100708
rect 442142 100472 442378 100708
rect 442462 100472 442698 100708
rect 442782 100472 443018 100708
rect 443102 100472 443338 100708
rect 443422 100472 443658 100708
rect 443742 100472 443978 100708
rect 444062 100472 444298 100708
rect 444382 100472 444618 100708
rect 440862 69836 441098 70072
rect 441182 69836 441418 70072
rect 441502 69836 441738 70072
rect 441822 69836 442058 70072
rect 442142 69836 442378 70072
rect 442462 69836 442698 70072
rect 442782 69836 443018 70072
rect 443102 69836 443338 70072
rect 443422 69836 443658 70072
rect 443742 69836 443978 70072
rect 444062 69836 444298 70072
rect 444382 69836 444618 70072
rect 440862 39200 441098 39436
rect 441182 39200 441418 39436
rect 441502 39200 441738 39436
rect 441822 39200 442058 39436
rect 442142 39200 442378 39436
rect 442462 39200 442698 39436
rect 442782 39200 443018 39436
rect 443102 39200 443338 39436
rect 443422 39200 443658 39436
rect 443742 39200 443978 39436
rect 444062 39200 444298 39436
rect 444382 39200 444618 39436
rect 122 3642 358 3878
rect 442 3642 678 3878
rect 762 3642 998 3878
rect 1082 3642 1318 3878
rect 1402 3642 1638 3878
rect 1722 3642 1958 3878
rect 2042 3642 2278 3878
rect 2362 3642 2598 3878
rect 2682 3642 2918 3878
rect 3002 3642 3238 3878
rect 3322 3642 3558 3878
rect 3642 3642 3878 3878
rect 122 3322 358 3558
rect 442 3322 678 3558
rect 762 3322 998 3558
rect 1082 3322 1318 3558
rect 1402 3322 1638 3558
rect 1722 3322 1958 3558
rect 2042 3322 2278 3558
rect 2362 3322 2598 3558
rect 2682 3322 2918 3558
rect 3002 3322 3238 3558
rect 3322 3322 3558 3558
rect 3642 3322 3878 3558
rect 122 3002 358 3238
rect 442 3002 678 3238
rect 762 3002 998 3238
rect 1082 3002 1318 3238
rect 1402 3002 1638 3238
rect 1722 3002 1958 3238
rect 2042 3002 2278 3238
rect 2362 3002 2598 3238
rect 2682 3002 2918 3238
rect 3002 3002 3238 3238
rect 3322 3002 3558 3238
rect 3642 3002 3878 3238
rect 122 2682 358 2918
rect 442 2682 678 2918
rect 762 2682 998 2918
rect 1082 2682 1318 2918
rect 1402 2682 1638 2918
rect 1722 2682 1958 2918
rect 2042 2682 2278 2918
rect 2362 2682 2598 2918
rect 2682 2682 2918 2918
rect 3002 2682 3238 2918
rect 3322 2682 3558 2918
rect 3642 2682 3878 2918
rect 122 2362 358 2598
rect 442 2362 678 2598
rect 762 2362 998 2598
rect 1082 2362 1318 2598
rect 1402 2362 1638 2598
rect 1722 2362 1958 2598
rect 2042 2362 2278 2598
rect 2362 2362 2598 2598
rect 2682 2362 2918 2598
rect 3002 2362 3238 2598
rect 3322 2362 3558 2598
rect 3642 2362 3878 2598
rect 122 2042 358 2278
rect 442 2042 678 2278
rect 762 2042 998 2278
rect 1082 2042 1318 2278
rect 1402 2042 1638 2278
rect 1722 2042 1958 2278
rect 2042 2042 2278 2278
rect 2362 2042 2598 2278
rect 2682 2042 2918 2278
rect 3002 2042 3238 2278
rect 3322 2042 3558 2278
rect 3642 2042 3878 2278
rect 122 1722 358 1958
rect 442 1722 678 1958
rect 762 1722 998 1958
rect 1082 1722 1318 1958
rect 1402 1722 1638 1958
rect 1722 1722 1958 1958
rect 2042 1722 2278 1958
rect 2362 1722 2598 1958
rect 2682 1722 2918 1958
rect 3002 1722 3238 1958
rect 3322 1722 3558 1958
rect 3642 1722 3878 1958
rect 122 1402 358 1638
rect 442 1402 678 1638
rect 762 1402 998 1638
rect 1082 1402 1318 1638
rect 1402 1402 1638 1638
rect 1722 1402 1958 1638
rect 2042 1402 2278 1638
rect 2362 1402 2598 1638
rect 2682 1402 2918 1638
rect 3002 1402 3238 1638
rect 3322 1402 3558 1638
rect 3642 1402 3878 1638
rect 122 1082 358 1318
rect 442 1082 678 1318
rect 762 1082 998 1318
rect 1082 1082 1318 1318
rect 1402 1082 1638 1318
rect 1722 1082 1958 1318
rect 2042 1082 2278 1318
rect 2362 1082 2598 1318
rect 2682 1082 2918 1318
rect 3002 1082 3238 1318
rect 3322 1082 3558 1318
rect 3642 1082 3878 1318
rect 122 762 358 998
rect 442 762 678 998
rect 762 762 998 998
rect 1082 762 1318 998
rect 1402 762 1638 998
rect 1722 762 1958 998
rect 2042 762 2278 998
rect 2362 762 2598 998
rect 2682 762 2918 998
rect 3002 762 3238 998
rect 3322 762 3558 998
rect 3642 762 3878 998
rect 122 442 358 678
rect 442 442 678 678
rect 762 442 998 678
rect 1082 442 1318 678
rect 1402 442 1638 678
rect 1722 442 1958 678
rect 2042 442 2278 678
rect 2362 442 2598 678
rect 2682 442 2918 678
rect 3002 442 3238 678
rect 3322 442 3558 678
rect 3642 442 3878 678
rect 122 122 358 358
rect 442 122 678 358
rect 762 122 998 358
rect 1082 122 1318 358
rect 1402 122 1638 358
rect 1722 122 1958 358
rect 2042 122 2278 358
rect 2362 122 2598 358
rect 2682 122 2918 358
rect 3002 122 3238 358
rect 3322 122 3558 358
rect 3642 122 3878 358
rect 440862 3642 441098 3878
rect 441182 3642 441418 3878
rect 441502 3642 441738 3878
rect 441822 3642 442058 3878
rect 442142 3642 442378 3878
rect 442462 3642 442698 3878
rect 442782 3642 443018 3878
rect 443102 3642 443338 3878
rect 443422 3642 443658 3878
rect 443742 3642 443978 3878
rect 444062 3642 444298 3878
rect 444382 3642 444618 3878
rect 440862 3322 441098 3558
rect 441182 3322 441418 3558
rect 441502 3322 441738 3558
rect 441822 3322 442058 3558
rect 442142 3322 442378 3558
rect 442462 3322 442698 3558
rect 442782 3322 443018 3558
rect 443102 3322 443338 3558
rect 443422 3322 443658 3558
rect 443742 3322 443978 3558
rect 444062 3322 444298 3558
rect 444382 3322 444618 3558
rect 440862 3002 441098 3238
rect 441182 3002 441418 3238
rect 441502 3002 441738 3238
rect 441822 3002 442058 3238
rect 442142 3002 442378 3238
rect 442462 3002 442698 3238
rect 442782 3002 443018 3238
rect 443102 3002 443338 3238
rect 443422 3002 443658 3238
rect 443742 3002 443978 3238
rect 444062 3002 444298 3238
rect 444382 3002 444618 3238
rect 440862 2682 441098 2918
rect 441182 2682 441418 2918
rect 441502 2682 441738 2918
rect 441822 2682 442058 2918
rect 442142 2682 442378 2918
rect 442462 2682 442698 2918
rect 442782 2682 443018 2918
rect 443102 2682 443338 2918
rect 443422 2682 443658 2918
rect 443742 2682 443978 2918
rect 444062 2682 444298 2918
rect 444382 2682 444618 2918
rect 440862 2362 441098 2598
rect 441182 2362 441418 2598
rect 441502 2362 441738 2598
rect 441822 2362 442058 2598
rect 442142 2362 442378 2598
rect 442462 2362 442698 2598
rect 442782 2362 443018 2598
rect 443102 2362 443338 2598
rect 443422 2362 443658 2598
rect 443742 2362 443978 2598
rect 444062 2362 444298 2598
rect 444382 2362 444618 2598
rect 440862 2042 441098 2278
rect 441182 2042 441418 2278
rect 441502 2042 441738 2278
rect 441822 2042 442058 2278
rect 442142 2042 442378 2278
rect 442462 2042 442698 2278
rect 442782 2042 443018 2278
rect 443102 2042 443338 2278
rect 443422 2042 443658 2278
rect 443742 2042 443978 2278
rect 444062 2042 444298 2278
rect 444382 2042 444618 2278
rect 440862 1722 441098 1958
rect 441182 1722 441418 1958
rect 441502 1722 441738 1958
rect 441822 1722 442058 1958
rect 442142 1722 442378 1958
rect 442462 1722 442698 1958
rect 442782 1722 443018 1958
rect 443102 1722 443338 1958
rect 443422 1722 443658 1958
rect 443742 1722 443978 1958
rect 444062 1722 444298 1958
rect 444382 1722 444618 1958
rect 440862 1402 441098 1638
rect 441182 1402 441418 1638
rect 441502 1402 441738 1638
rect 441822 1402 442058 1638
rect 442142 1402 442378 1638
rect 442462 1402 442698 1638
rect 442782 1402 443018 1638
rect 443102 1402 443338 1638
rect 443422 1402 443658 1638
rect 443742 1402 443978 1638
rect 444062 1402 444298 1638
rect 444382 1402 444618 1638
rect 440862 1082 441098 1318
rect 441182 1082 441418 1318
rect 441502 1082 441738 1318
rect 441822 1082 442058 1318
rect 442142 1082 442378 1318
rect 442462 1082 442698 1318
rect 442782 1082 443018 1318
rect 443102 1082 443338 1318
rect 443422 1082 443658 1318
rect 443742 1082 443978 1318
rect 444062 1082 444298 1318
rect 444382 1082 444618 1318
rect 440862 762 441098 998
rect 441182 762 441418 998
rect 441502 762 441738 998
rect 441822 762 442058 998
rect 442142 762 442378 998
rect 442462 762 442698 998
rect 442782 762 443018 998
rect 443102 762 443338 998
rect 443422 762 443658 998
rect 443742 762 443978 998
rect 444062 762 444298 998
rect 444382 762 444618 998
rect 440862 442 441098 678
rect 441182 442 441418 678
rect 441502 442 441738 678
rect 441822 442 442058 678
rect 442142 442 442378 678
rect 442462 442 442698 678
rect 442782 442 443018 678
rect 443102 442 443338 678
rect 443422 442 443658 678
rect 443742 442 443978 678
rect 444062 442 444298 678
rect 444382 442 444618 678
rect 440862 122 441098 358
rect 441182 122 441418 358
rect 441502 122 441738 358
rect 441822 122 442058 358
rect 442142 122 442378 358
rect 442462 122 442698 358
rect 442782 122 443018 358
rect 443102 122 443338 358
rect 443422 122 443658 358
rect 443742 122 443978 358
rect 444062 122 444298 358
rect 444382 122 444618 358
<< metal5 >>
rect 0 405398 444740 405520
rect 0 405162 122 405398
rect 358 405162 442 405398
rect 678 405162 762 405398
rect 998 405162 1082 405398
rect 1318 405162 1402 405398
rect 1638 405162 1722 405398
rect 1958 405162 2042 405398
rect 2278 405162 2362 405398
rect 2598 405162 2682 405398
rect 2918 405162 3002 405398
rect 3238 405162 3322 405398
rect 3558 405162 3642 405398
rect 3878 405162 440862 405398
rect 441098 405162 441182 405398
rect 441418 405162 441502 405398
rect 441738 405162 441822 405398
rect 442058 405162 442142 405398
rect 442378 405162 442462 405398
rect 442698 405162 442782 405398
rect 443018 405162 443102 405398
rect 443338 405162 443422 405398
rect 443658 405162 443742 405398
rect 443978 405162 444062 405398
rect 444298 405162 444382 405398
rect 444618 405162 444740 405398
rect 0 405078 444740 405162
rect 0 404842 122 405078
rect 358 404842 442 405078
rect 678 404842 762 405078
rect 998 404842 1082 405078
rect 1318 404842 1402 405078
rect 1638 404842 1722 405078
rect 1958 404842 2042 405078
rect 2278 404842 2362 405078
rect 2598 404842 2682 405078
rect 2918 404842 3002 405078
rect 3238 404842 3322 405078
rect 3558 404842 3642 405078
rect 3878 404842 440862 405078
rect 441098 404842 441182 405078
rect 441418 404842 441502 405078
rect 441738 404842 441822 405078
rect 442058 404842 442142 405078
rect 442378 404842 442462 405078
rect 442698 404842 442782 405078
rect 443018 404842 443102 405078
rect 443338 404842 443422 405078
rect 443658 404842 443742 405078
rect 443978 404842 444062 405078
rect 444298 404842 444382 405078
rect 444618 404842 444740 405078
rect 0 404758 444740 404842
rect 0 404522 122 404758
rect 358 404522 442 404758
rect 678 404522 762 404758
rect 998 404522 1082 404758
rect 1318 404522 1402 404758
rect 1638 404522 1722 404758
rect 1958 404522 2042 404758
rect 2278 404522 2362 404758
rect 2598 404522 2682 404758
rect 2918 404522 3002 404758
rect 3238 404522 3322 404758
rect 3558 404522 3642 404758
rect 3878 404522 440862 404758
rect 441098 404522 441182 404758
rect 441418 404522 441502 404758
rect 441738 404522 441822 404758
rect 442058 404522 442142 404758
rect 442378 404522 442462 404758
rect 442698 404522 442782 404758
rect 443018 404522 443102 404758
rect 443338 404522 443422 404758
rect 443658 404522 443742 404758
rect 443978 404522 444062 404758
rect 444298 404522 444382 404758
rect 444618 404522 444740 404758
rect 0 404438 444740 404522
rect 0 404202 122 404438
rect 358 404202 442 404438
rect 678 404202 762 404438
rect 998 404202 1082 404438
rect 1318 404202 1402 404438
rect 1638 404202 1722 404438
rect 1958 404202 2042 404438
rect 2278 404202 2362 404438
rect 2598 404202 2682 404438
rect 2918 404202 3002 404438
rect 3238 404202 3322 404438
rect 3558 404202 3642 404438
rect 3878 404202 440862 404438
rect 441098 404202 441182 404438
rect 441418 404202 441502 404438
rect 441738 404202 441822 404438
rect 442058 404202 442142 404438
rect 442378 404202 442462 404438
rect 442698 404202 442782 404438
rect 443018 404202 443102 404438
rect 443338 404202 443422 404438
rect 443658 404202 443742 404438
rect 443978 404202 444062 404438
rect 444298 404202 444382 404438
rect 444618 404202 444740 404438
rect 0 404118 444740 404202
rect 0 403882 122 404118
rect 358 403882 442 404118
rect 678 403882 762 404118
rect 998 403882 1082 404118
rect 1318 403882 1402 404118
rect 1638 403882 1722 404118
rect 1958 403882 2042 404118
rect 2278 403882 2362 404118
rect 2598 403882 2682 404118
rect 2918 403882 3002 404118
rect 3238 403882 3322 404118
rect 3558 403882 3642 404118
rect 3878 403882 440862 404118
rect 441098 403882 441182 404118
rect 441418 403882 441502 404118
rect 441738 403882 441822 404118
rect 442058 403882 442142 404118
rect 442378 403882 442462 404118
rect 442698 403882 442782 404118
rect 443018 403882 443102 404118
rect 443338 403882 443422 404118
rect 443658 403882 443742 404118
rect 443978 403882 444062 404118
rect 444298 403882 444382 404118
rect 444618 403882 444740 404118
rect 0 403798 444740 403882
rect 0 403562 122 403798
rect 358 403562 442 403798
rect 678 403562 762 403798
rect 998 403562 1082 403798
rect 1318 403562 1402 403798
rect 1638 403562 1722 403798
rect 1958 403562 2042 403798
rect 2278 403562 2362 403798
rect 2598 403562 2682 403798
rect 2918 403562 3002 403798
rect 3238 403562 3322 403798
rect 3558 403562 3642 403798
rect 3878 403562 440862 403798
rect 441098 403562 441182 403798
rect 441418 403562 441502 403798
rect 441738 403562 441822 403798
rect 442058 403562 442142 403798
rect 442378 403562 442462 403798
rect 442698 403562 442782 403798
rect 443018 403562 443102 403798
rect 443338 403562 443422 403798
rect 443658 403562 443742 403798
rect 443978 403562 444062 403798
rect 444298 403562 444382 403798
rect 444618 403562 444740 403798
rect 0 403478 444740 403562
rect 0 403242 122 403478
rect 358 403242 442 403478
rect 678 403242 762 403478
rect 998 403242 1082 403478
rect 1318 403242 1402 403478
rect 1638 403242 1722 403478
rect 1958 403242 2042 403478
rect 2278 403242 2362 403478
rect 2598 403242 2682 403478
rect 2918 403242 3002 403478
rect 3238 403242 3322 403478
rect 3558 403242 3642 403478
rect 3878 403242 440862 403478
rect 441098 403242 441182 403478
rect 441418 403242 441502 403478
rect 441738 403242 441822 403478
rect 442058 403242 442142 403478
rect 442378 403242 442462 403478
rect 442698 403242 442782 403478
rect 443018 403242 443102 403478
rect 443338 403242 443422 403478
rect 443658 403242 443742 403478
rect 443978 403242 444062 403478
rect 444298 403242 444382 403478
rect 444618 403242 444740 403478
rect 0 403158 444740 403242
rect 0 402922 122 403158
rect 358 402922 442 403158
rect 678 402922 762 403158
rect 998 402922 1082 403158
rect 1318 402922 1402 403158
rect 1638 402922 1722 403158
rect 1958 402922 2042 403158
rect 2278 402922 2362 403158
rect 2598 402922 2682 403158
rect 2918 402922 3002 403158
rect 3238 402922 3322 403158
rect 3558 402922 3642 403158
rect 3878 402922 440862 403158
rect 441098 402922 441182 403158
rect 441418 402922 441502 403158
rect 441738 402922 441822 403158
rect 442058 402922 442142 403158
rect 442378 402922 442462 403158
rect 442698 402922 442782 403158
rect 443018 402922 443102 403158
rect 443338 402922 443422 403158
rect 443658 402922 443742 403158
rect 443978 402922 444062 403158
rect 444298 402922 444382 403158
rect 444618 402922 444740 403158
rect 0 402838 444740 402922
rect 0 402602 122 402838
rect 358 402602 442 402838
rect 678 402602 762 402838
rect 998 402602 1082 402838
rect 1318 402602 1402 402838
rect 1638 402602 1722 402838
rect 1958 402602 2042 402838
rect 2278 402602 2362 402838
rect 2598 402602 2682 402838
rect 2918 402602 3002 402838
rect 3238 402602 3322 402838
rect 3558 402602 3642 402838
rect 3878 402602 440862 402838
rect 441098 402602 441182 402838
rect 441418 402602 441502 402838
rect 441738 402602 441822 402838
rect 442058 402602 442142 402838
rect 442378 402602 442462 402838
rect 442698 402602 442782 402838
rect 443018 402602 443102 402838
rect 443338 402602 443422 402838
rect 443658 402602 443742 402838
rect 443978 402602 444062 402838
rect 444298 402602 444382 402838
rect 444618 402602 444740 402838
rect 0 402518 444740 402602
rect 0 402282 122 402518
rect 358 402282 442 402518
rect 678 402282 762 402518
rect 998 402282 1082 402518
rect 1318 402282 1402 402518
rect 1638 402282 1722 402518
rect 1958 402282 2042 402518
rect 2278 402282 2362 402518
rect 2598 402282 2682 402518
rect 2918 402282 3002 402518
rect 3238 402282 3322 402518
rect 3558 402282 3642 402518
rect 3878 402282 440862 402518
rect 441098 402282 441182 402518
rect 441418 402282 441502 402518
rect 441738 402282 441822 402518
rect 442058 402282 442142 402518
rect 442378 402282 442462 402518
rect 442698 402282 442782 402518
rect 443018 402282 443102 402518
rect 443338 402282 443422 402518
rect 443658 402282 443742 402518
rect 443978 402282 444062 402518
rect 444298 402282 444382 402518
rect 444618 402282 444740 402518
rect 0 402198 444740 402282
rect 0 401962 122 402198
rect 358 401962 442 402198
rect 678 401962 762 402198
rect 998 401962 1082 402198
rect 1318 401962 1402 402198
rect 1638 401962 1722 402198
rect 1958 401962 2042 402198
rect 2278 401962 2362 402198
rect 2598 401962 2682 402198
rect 2918 401962 3002 402198
rect 3238 401962 3322 402198
rect 3558 401962 3642 402198
rect 3878 401962 440862 402198
rect 441098 401962 441182 402198
rect 441418 401962 441502 402198
rect 441738 401962 441822 402198
rect 442058 401962 442142 402198
rect 442378 401962 442462 402198
rect 442698 401962 442782 402198
rect 443018 401962 443102 402198
rect 443338 401962 443422 402198
rect 443658 401962 443742 402198
rect 443978 401962 444062 402198
rect 444298 401962 444382 402198
rect 444618 401962 444740 402198
rect 0 401878 444740 401962
rect 0 401642 122 401878
rect 358 401642 442 401878
rect 678 401642 762 401878
rect 998 401642 1082 401878
rect 1318 401642 1402 401878
rect 1638 401642 1722 401878
rect 1958 401642 2042 401878
rect 2278 401642 2362 401878
rect 2598 401642 2682 401878
rect 2918 401642 3002 401878
rect 3238 401642 3322 401878
rect 3558 401642 3642 401878
rect 3878 401642 440862 401878
rect 441098 401642 441182 401878
rect 441418 401642 441502 401878
rect 441738 401642 441822 401878
rect 442058 401642 442142 401878
rect 442378 401642 442462 401878
rect 442698 401642 442782 401878
rect 443018 401642 443102 401878
rect 443338 401642 443422 401878
rect 443658 401642 443742 401878
rect 443978 401642 444062 401878
rect 444298 401642 444382 401878
rect 444618 401642 444740 401878
rect 0 401520 444740 401642
rect 5000 400398 439740 400520
rect 5000 400162 5122 400398
rect 5358 400162 5442 400398
rect 5678 400162 5762 400398
rect 5998 400162 6082 400398
rect 6318 400162 6402 400398
rect 6638 400162 6722 400398
rect 6958 400162 7042 400398
rect 7278 400162 7362 400398
rect 7598 400162 7682 400398
rect 7918 400162 8002 400398
rect 8238 400162 8322 400398
rect 8558 400162 8642 400398
rect 8878 400162 435862 400398
rect 436098 400162 436182 400398
rect 436418 400162 436502 400398
rect 436738 400162 436822 400398
rect 437058 400162 437142 400398
rect 437378 400162 437462 400398
rect 437698 400162 437782 400398
rect 438018 400162 438102 400398
rect 438338 400162 438422 400398
rect 438658 400162 438742 400398
rect 438978 400162 439062 400398
rect 439298 400162 439382 400398
rect 439618 400162 439740 400398
rect 5000 400078 439740 400162
rect 5000 399842 5122 400078
rect 5358 399842 5442 400078
rect 5678 399842 5762 400078
rect 5998 399842 6082 400078
rect 6318 399842 6402 400078
rect 6638 399842 6722 400078
rect 6958 399842 7042 400078
rect 7278 399842 7362 400078
rect 7598 399842 7682 400078
rect 7918 399842 8002 400078
rect 8238 399842 8322 400078
rect 8558 399842 8642 400078
rect 8878 399842 435862 400078
rect 436098 399842 436182 400078
rect 436418 399842 436502 400078
rect 436738 399842 436822 400078
rect 437058 399842 437142 400078
rect 437378 399842 437462 400078
rect 437698 399842 437782 400078
rect 438018 399842 438102 400078
rect 438338 399842 438422 400078
rect 438658 399842 438742 400078
rect 438978 399842 439062 400078
rect 439298 399842 439382 400078
rect 439618 399842 439740 400078
rect 5000 399758 439740 399842
rect 5000 399522 5122 399758
rect 5358 399522 5442 399758
rect 5678 399522 5762 399758
rect 5998 399522 6082 399758
rect 6318 399522 6402 399758
rect 6638 399522 6722 399758
rect 6958 399522 7042 399758
rect 7278 399522 7362 399758
rect 7598 399522 7682 399758
rect 7918 399522 8002 399758
rect 8238 399522 8322 399758
rect 8558 399522 8642 399758
rect 8878 399522 435862 399758
rect 436098 399522 436182 399758
rect 436418 399522 436502 399758
rect 436738 399522 436822 399758
rect 437058 399522 437142 399758
rect 437378 399522 437462 399758
rect 437698 399522 437782 399758
rect 438018 399522 438102 399758
rect 438338 399522 438422 399758
rect 438658 399522 438742 399758
rect 438978 399522 439062 399758
rect 439298 399522 439382 399758
rect 439618 399522 439740 399758
rect 5000 399438 439740 399522
rect 5000 399202 5122 399438
rect 5358 399202 5442 399438
rect 5678 399202 5762 399438
rect 5998 399202 6082 399438
rect 6318 399202 6402 399438
rect 6638 399202 6722 399438
rect 6958 399202 7042 399438
rect 7278 399202 7362 399438
rect 7598 399202 7682 399438
rect 7918 399202 8002 399438
rect 8238 399202 8322 399438
rect 8558 399202 8642 399438
rect 8878 399202 435862 399438
rect 436098 399202 436182 399438
rect 436418 399202 436502 399438
rect 436738 399202 436822 399438
rect 437058 399202 437142 399438
rect 437378 399202 437462 399438
rect 437698 399202 437782 399438
rect 438018 399202 438102 399438
rect 438338 399202 438422 399438
rect 438658 399202 438742 399438
rect 438978 399202 439062 399438
rect 439298 399202 439382 399438
rect 439618 399202 439740 399438
rect 5000 399118 439740 399202
rect 5000 398882 5122 399118
rect 5358 398882 5442 399118
rect 5678 398882 5762 399118
rect 5998 398882 6082 399118
rect 6318 398882 6402 399118
rect 6638 398882 6722 399118
rect 6958 398882 7042 399118
rect 7278 398882 7362 399118
rect 7598 398882 7682 399118
rect 7918 398882 8002 399118
rect 8238 398882 8322 399118
rect 8558 398882 8642 399118
rect 8878 398882 435862 399118
rect 436098 398882 436182 399118
rect 436418 398882 436502 399118
rect 436738 398882 436822 399118
rect 437058 398882 437142 399118
rect 437378 398882 437462 399118
rect 437698 398882 437782 399118
rect 438018 398882 438102 399118
rect 438338 398882 438422 399118
rect 438658 398882 438742 399118
rect 438978 398882 439062 399118
rect 439298 398882 439382 399118
rect 439618 398882 439740 399118
rect 5000 398798 439740 398882
rect 5000 398562 5122 398798
rect 5358 398562 5442 398798
rect 5678 398562 5762 398798
rect 5998 398562 6082 398798
rect 6318 398562 6402 398798
rect 6638 398562 6722 398798
rect 6958 398562 7042 398798
rect 7278 398562 7362 398798
rect 7598 398562 7682 398798
rect 7918 398562 8002 398798
rect 8238 398562 8322 398798
rect 8558 398562 8642 398798
rect 8878 398562 435862 398798
rect 436098 398562 436182 398798
rect 436418 398562 436502 398798
rect 436738 398562 436822 398798
rect 437058 398562 437142 398798
rect 437378 398562 437462 398798
rect 437698 398562 437782 398798
rect 438018 398562 438102 398798
rect 438338 398562 438422 398798
rect 438658 398562 438742 398798
rect 438978 398562 439062 398798
rect 439298 398562 439382 398798
rect 439618 398562 439740 398798
rect 5000 398478 439740 398562
rect 5000 398242 5122 398478
rect 5358 398242 5442 398478
rect 5678 398242 5762 398478
rect 5998 398242 6082 398478
rect 6318 398242 6402 398478
rect 6638 398242 6722 398478
rect 6958 398242 7042 398478
rect 7278 398242 7362 398478
rect 7598 398242 7682 398478
rect 7918 398242 8002 398478
rect 8238 398242 8322 398478
rect 8558 398242 8642 398478
rect 8878 398242 435862 398478
rect 436098 398242 436182 398478
rect 436418 398242 436502 398478
rect 436738 398242 436822 398478
rect 437058 398242 437142 398478
rect 437378 398242 437462 398478
rect 437698 398242 437782 398478
rect 438018 398242 438102 398478
rect 438338 398242 438422 398478
rect 438658 398242 438742 398478
rect 438978 398242 439062 398478
rect 439298 398242 439382 398478
rect 439618 398242 439740 398478
rect 5000 398158 439740 398242
rect 5000 397922 5122 398158
rect 5358 397922 5442 398158
rect 5678 397922 5762 398158
rect 5998 397922 6082 398158
rect 6318 397922 6402 398158
rect 6638 397922 6722 398158
rect 6958 397922 7042 398158
rect 7278 397922 7362 398158
rect 7598 397922 7682 398158
rect 7918 397922 8002 398158
rect 8238 397922 8322 398158
rect 8558 397922 8642 398158
rect 8878 397922 435862 398158
rect 436098 397922 436182 398158
rect 436418 397922 436502 398158
rect 436738 397922 436822 398158
rect 437058 397922 437142 398158
rect 437378 397922 437462 398158
rect 437698 397922 437782 398158
rect 438018 397922 438102 398158
rect 438338 397922 438422 398158
rect 438658 397922 438742 398158
rect 438978 397922 439062 398158
rect 439298 397922 439382 398158
rect 439618 397922 439740 398158
rect 5000 397838 439740 397922
rect 5000 397602 5122 397838
rect 5358 397602 5442 397838
rect 5678 397602 5762 397838
rect 5998 397602 6082 397838
rect 6318 397602 6402 397838
rect 6638 397602 6722 397838
rect 6958 397602 7042 397838
rect 7278 397602 7362 397838
rect 7598 397602 7682 397838
rect 7918 397602 8002 397838
rect 8238 397602 8322 397838
rect 8558 397602 8642 397838
rect 8878 397602 435862 397838
rect 436098 397602 436182 397838
rect 436418 397602 436502 397838
rect 436738 397602 436822 397838
rect 437058 397602 437142 397838
rect 437378 397602 437462 397838
rect 437698 397602 437782 397838
rect 438018 397602 438102 397838
rect 438338 397602 438422 397838
rect 438658 397602 438742 397838
rect 438978 397602 439062 397838
rect 439298 397602 439382 397838
rect 439618 397602 439740 397838
rect 5000 397518 439740 397602
rect 5000 397282 5122 397518
rect 5358 397282 5442 397518
rect 5678 397282 5762 397518
rect 5998 397282 6082 397518
rect 6318 397282 6402 397518
rect 6638 397282 6722 397518
rect 6958 397282 7042 397518
rect 7278 397282 7362 397518
rect 7598 397282 7682 397518
rect 7918 397282 8002 397518
rect 8238 397282 8322 397518
rect 8558 397282 8642 397518
rect 8878 397282 435862 397518
rect 436098 397282 436182 397518
rect 436418 397282 436502 397518
rect 436738 397282 436822 397518
rect 437058 397282 437142 397518
rect 437378 397282 437462 397518
rect 437698 397282 437782 397518
rect 438018 397282 438102 397518
rect 438338 397282 438422 397518
rect 438658 397282 438742 397518
rect 438978 397282 439062 397518
rect 439298 397282 439382 397518
rect 439618 397282 439740 397518
rect 5000 397198 439740 397282
rect 5000 396962 5122 397198
rect 5358 396962 5442 397198
rect 5678 396962 5762 397198
rect 5998 396962 6082 397198
rect 6318 396962 6402 397198
rect 6638 396962 6722 397198
rect 6958 396962 7042 397198
rect 7278 396962 7362 397198
rect 7598 396962 7682 397198
rect 7918 396962 8002 397198
rect 8238 396962 8322 397198
rect 8558 396962 8642 397198
rect 8878 396962 435862 397198
rect 436098 396962 436182 397198
rect 436418 396962 436502 397198
rect 436738 396962 436822 397198
rect 437058 396962 437142 397198
rect 437378 396962 437462 397198
rect 437698 396962 437782 397198
rect 438018 396962 438102 397198
rect 438338 396962 438422 397198
rect 438658 396962 438742 397198
rect 438978 396962 439062 397198
rect 439298 396962 439382 397198
rect 439618 396962 439740 397198
rect 5000 396878 439740 396962
rect 5000 396642 5122 396878
rect 5358 396642 5442 396878
rect 5678 396642 5762 396878
rect 5998 396642 6082 396878
rect 6318 396642 6402 396878
rect 6638 396642 6722 396878
rect 6958 396642 7042 396878
rect 7278 396642 7362 396878
rect 7598 396642 7682 396878
rect 7918 396642 8002 396878
rect 8238 396642 8322 396878
rect 8558 396642 8642 396878
rect 8878 396642 435862 396878
rect 436098 396642 436182 396878
rect 436418 396642 436502 396878
rect 436738 396642 436822 396878
rect 437058 396642 437142 396878
rect 437378 396642 437462 396878
rect 437698 396642 437782 396878
rect 438018 396642 438102 396878
rect 438338 396642 438422 396878
rect 438658 396642 438742 396878
rect 438978 396642 439062 396878
rect 439298 396642 439382 396878
rect 439618 396642 439740 396878
rect 5000 396520 439740 396642
rect 0 391750 444740 391792
rect 0 391514 5122 391750
rect 5358 391514 5442 391750
rect 5678 391514 5762 391750
rect 5998 391514 6082 391750
rect 6318 391514 6402 391750
rect 6638 391514 6722 391750
rect 6958 391514 7042 391750
rect 7278 391514 7362 391750
rect 7598 391514 7682 391750
rect 7918 391514 8002 391750
rect 8238 391514 8322 391750
rect 8558 391514 8642 391750
rect 8878 391514 435862 391750
rect 436098 391514 436182 391750
rect 436418 391514 436502 391750
rect 436738 391514 436822 391750
rect 437058 391514 437142 391750
rect 437378 391514 437462 391750
rect 437698 391514 437782 391750
rect 438018 391514 438102 391750
rect 438338 391514 438422 391750
rect 438658 391514 438742 391750
rect 438978 391514 439062 391750
rect 439298 391514 439382 391750
rect 439618 391514 444740 391750
rect 0 391472 444740 391514
rect 0 376432 444740 376474
rect 0 376196 122 376432
rect 358 376196 442 376432
rect 678 376196 762 376432
rect 998 376196 1082 376432
rect 1318 376196 1402 376432
rect 1638 376196 1722 376432
rect 1958 376196 2042 376432
rect 2278 376196 2362 376432
rect 2598 376196 2682 376432
rect 2918 376196 3002 376432
rect 3238 376196 3322 376432
rect 3558 376196 3642 376432
rect 3878 376196 440862 376432
rect 441098 376196 441182 376432
rect 441418 376196 441502 376432
rect 441738 376196 441822 376432
rect 442058 376196 442142 376432
rect 442378 376196 442462 376432
rect 442698 376196 442782 376432
rect 443018 376196 443102 376432
rect 443338 376196 443422 376432
rect 443658 376196 443742 376432
rect 443978 376196 444062 376432
rect 444298 376196 444382 376432
rect 444618 376196 444740 376432
rect 0 376154 444740 376196
rect 0 361114 444740 361156
rect 0 360878 5122 361114
rect 5358 360878 5442 361114
rect 5678 360878 5762 361114
rect 5998 360878 6082 361114
rect 6318 360878 6402 361114
rect 6638 360878 6722 361114
rect 6958 360878 7042 361114
rect 7278 360878 7362 361114
rect 7598 360878 7682 361114
rect 7918 360878 8002 361114
rect 8238 360878 8322 361114
rect 8558 360878 8642 361114
rect 8878 360878 435862 361114
rect 436098 360878 436182 361114
rect 436418 360878 436502 361114
rect 436738 360878 436822 361114
rect 437058 360878 437142 361114
rect 437378 360878 437462 361114
rect 437698 360878 437782 361114
rect 438018 360878 438102 361114
rect 438338 360878 438422 361114
rect 438658 360878 438742 361114
rect 438978 360878 439062 361114
rect 439298 360878 439382 361114
rect 439618 360878 444740 361114
rect 0 360836 444740 360878
rect 0 345796 444740 345838
rect 0 345560 122 345796
rect 358 345560 442 345796
rect 678 345560 762 345796
rect 998 345560 1082 345796
rect 1318 345560 1402 345796
rect 1638 345560 1722 345796
rect 1958 345560 2042 345796
rect 2278 345560 2362 345796
rect 2598 345560 2682 345796
rect 2918 345560 3002 345796
rect 3238 345560 3322 345796
rect 3558 345560 3642 345796
rect 3878 345560 440862 345796
rect 441098 345560 441182 345796
rect 441418 345560 441502 345796
rect 441738 345560 441822 345796
rect 442058 345560 442142 345796
rect 442378 345560 442462 345796
rect 442698 345560 442782 345796
rect 443018 345560 443102 345796
rect 443338 345560 443422 345796
rect 443658 345560 443742 345796
rect 443978 345560 444062 345796
rect 444298 345560 444382 345796
rect 444618 345560 444740 345796
rect 0 345518 444740 345560
rect 231732 333642 306388 333684
rect 231732 333406 231774 333642
rect 232010 333406 262318 333642
rect 262554 333406 306110 333642
rect 306346 333406 306388 333642
rect 231732 333364 306388 333406
rect 137156 332282 198932 332324
rect 137156 332046 137198 332282
rect 137434 332046 168478 332282
rect 168714 332046 198654 332282
rect 198890 332046 198932 332282
rect 137156 332004 198932 332046
rect 231732 332282 296268 332324
rect 231732 332046 231774 332282
rect 232010 332046 295990 332282
rect 296226 332046 296268 332282
rect 231732 332004 296268 332046
rect 137156 331602 204636 331644
rect 137156 331366 137198 331602
rect 137434 331366 159462 331602
rect 159698 331366 204358 331602
rect 204594 331366 204636 331602
rect 137156 331324 204636 331366
rect 231732 331602 251740 331644
rect 231732 331366 231774 331602
rect 232010 331366 251462 331602
rect 251698 331366 251740 331602
rect 231732 331324 251740 331366
rect 252156 331602 252476 332004
rect 252156 331366 252198 331602
rect 252434 331366 252476 331602
rect 252156 331324 252476 331366
rect 252892 331602 294244 331644
rect 252892 331366 252934 331602
rect 253170 331366 293966 331602
rect 294202 331366 294244 331602
rect 252892 331324 294244 331366
rect 0 330478 444740 330520
rect 0 330242 5122 330478
rect 5358 330242 5442 330478
rect 5678 330242 5762 330478
rect 5998 330242 6082 330478
rect 6318 330242 6402 330478
rect 6638 330242 6722 330478
rect 6958 330242 7042 330478
rect 7278 330242 7362 330478
rect 7598 330242 7682 330478
rect 7918 330242 8002 330478
rect 8238 330242 8322 330478
rect 8558 330242 8642 330478
rect 8878 330242 435862 330478
rect 436098 330242 436182 330478
rect 436418 330242 436502 330478
rect 436738 330242 436822 330478
rect 437058 330242 437142 330478
rect 437378 330242 437462 330478
rect 437698 330242 437782 330478
rect 438018 330242 438102 330478
rect 438338 330242 438422 330478
rect 438658 330242 438742 330478
rect 438978 330242 439062 330478
rect 439298 330242 439382 330478
rect 439618 330242 444740 330478
rect 0 330200 444740 330242
rect 161628 329562 212364 329604
rect 161628 329326 161670 329562
rect 161906 329326 212086 329562
rect 212322 329326 212364 329562
rect 161628 329284 212364 329326
rect 104588 320042 105092 320084
rect 104588 319806 104814 320042
rect 105050 319806 105092 320042
rect 104588 319764 105092 319806
rect 104588 315962 104908 319764
rect 104588 315726 104630 315962
rect 104866 315726 104908 315962
rect 104588 315684 104908 315726
rect 0 315160 444740 315202
rect 0 314924 122 315160
rect 358 314924 442 315160
rect 678 314924 762 315160
rect 998 314924 1082 315160
rect 1318 314924 1402 315160
rect 1638 314924 1722 315160
rect 1958 314924 2042 315160
rect 2278 314924 2362 315160
rect 2598 314924 2682 315160
rect 2918 314924 3002 315160
rect 3238 314924 3322 315160
rect 3558 314924 3642 315160
rect 3878 314924 104506 315160
rect 104742 314924 198506 315160
rect 198742 314924 292506 315160
rect 292742 314924 440862 315160
rect 441098 314924 441182 315160
rect 441418 314924 441502 315160
rect 441738 314924 441822 315160
rect 442058 314924 442142 315160
rect 442378 314924 442462 315160
rect 442698 314924 442782 315160
rect 443018 314924 443102 315160
rect 443338 314924 443422 315160
rect 443658 314924 443742 315160
rect 443978 314924 444062 315160
rect 444298 314924 444382 315160
rect 444618 314924 444740 315160
rect 0 314882 444740 314924
rect 104588 314602 104908 314644
rect 104588 314366 104630 314602
rect 104866 314366 104908 314602
rect 104588 306484 104908 314366
rect 103852 306164 104908 306484
rect 103852 301044 104172 306164
rect 103852 301002 104908 301044
rect 103852 300766 104630 301002
rect 104866 300766 104908 301002
rect 103852 300724 104908 300766
rect 0 299842 444740 299884
rect 0 299606 5122 299842
rect 5358 299606 5442 299842
rect 5678 299606 5762 299842
rect 5998 299606 6082 299842
rect 6318 299606 6402 299842
rect 6638 299606 6722 299842
rect 6958 299606 7042 299842
rect 7278 299606 7362 299842
rect 7598 299606 7682 299842
rect 7918 299606 8002 299842
rect 8238 299606 8322 299842
rect 8558 299606 8642 299842
rect 8878 299606 89146 299842
rect 89382 299642 183146 299842
rect 89382 299606 104446 299642
rect 0 299564 104446 299606
rect 104404 299406 104446 299564
rect 104682 299606 183146 299642
rect 183382 299606 277146 299842
rect 277382 299606 435862 299842
rect 436098 299606 436182 299842
rect 436418 299606 436502 299842
rect 436738 299606 436822 299842
rect 437058 299606 437142 299842
rect 437378 299606 437462 299842
rect 437698 299606 437782 299842
rect 438018 299606 438102 299842
rect 438338 299606 438422 299842
rect 438658 299606 438742 299842
rect 438978 299606 439062 299842
rect 439298 299606 439382 299842
rect 439618 299606 444740 299842
rect 104682 299564 444740 299606
rect 104682 299406 104724 299564
rect 104404 296964 104724 299406
rect 118756 298282 134900 298324
rect 118756 298046 134622 298282
rect 134858 298046 134900 298282
rect 118756 298004 134900 298046
rect 118756 296964 119076 298004
rect 104404 296644 119076 296964
rect 104404 296284 104724 296644
rect 104404 295964 105828 296284
rect 105508 291524 105828 295964
rect 231732 295562 323684 295604
rect 231732 295326 231774 295562
rect 232010 295326 323406 295562
rect 323642 295326 323684 295562
rect 231732 295284 323684 295326
rect 136788 294882 228924 294924
rect 136788 294646 136830 294882
rect 137066 294646 228646 294882
rect 228882 294646 228924 294882
rect 136788 294604 228924 294646
rect 280492 293924 289828 294244
rect 280492 292204 280812 293924
rect 136788 292162 280812 292204
rect 136788 291926 136830 292162
rect 137066 291926 230670 292162
rect 230906 291926 280812 292162
rect 136788 291884 280812 291926
rect 289508 292204 289828 293924
rect 299812 293924 309148 294244
rect 299812 292204 300132 293924
rect 289508 291884 300132 292204
rect 308828 292204 309148 293924
rect 308828 292162 322948 292204
rect 308828 291926 322670 292162
rect 322906 291926 322948 292162
rect 308828 291884 322948 291926
rect 104404 291204 105828 291524
rect 98884 286444 100308 286764
rect 98884 286084 99204 286444
rect 92628 285764 99204 286084
rect 99988 286084 100308 286444
rect 104404 286322 104724 291204
rect 215356 290524 225428 290844
rect 215356 289484 215676 290524
rect 137892 289442 215676 289484
rect 137892 289206 137934 289442
rect 138170 289206 215676 289442
rect 137892 289164 215676 289206
rect 225108 289484 225428 290524
rect 234308 290524 241988 290844
rect 234308 289484 234628 290524
rect 241668 290164 241988 290524
rect 253812 290802 261308 290844
rect 253812 290566 261030 290802
rect 261266 290566 261308 290802
rect 253812 290524 261308 290566
rect 273132 290524 289828 290844
rect 241668 289844 251372 290164
rect 225108 289442 234628 289484
rect 225108 289206 228646 289442
rect 228882 289206 234628 289442
rect 225108 289164 234628 289206
rect 251052 289484 251372 289844
rect 253812 289484 254132 290524
rect 273132 289484 273452 290524
rect 251052 289164 254132 289484
rect 270372 289442 273452 289484
rect 270372 289206 270414 289442
rect 270650 289206 273452 289442
rect 270372 289164 273452 289206
rect 289508 289484 289828 290524
rect 292452 290524 309148 290844
rect 292452 289484 292772 290524
rect 289508 289164 292772 289484
rect 308828 289484 309148 290524
rect 311772 290524 319268 290844
rect 311772 289484 312092 290524
rect 308828 289164 312092 289484
rect 318948 289484 319268 290524
rect 318948 289442 323316 289484
rect 318948 289206 323038 289442
rect 323274 289206 323316 289442
rect 318948 289164 323316 289206
rect 104404 286086 104446 286322
rect 104682 286086 104724 286322
rect 99988 285764 101228 286084
rect 104404 286044 104724 286086
rect 106060 286444 113372 286764
rect 92628 285404 92948 285764
rect 84532 285362 92948 285404
rect 84532 285126 84574 285362
rect 84810 285126 92948 285362
rect 84532 285084 92948 285126
rect 100908 285404 101228 285764
rect 106060 285404 106380 286444
rect 100908 285084 106380 285404
rect 113052 285404 113372 286444
rect 113052 285362 135084 285404
rect 113052 285126 134806 285362
rect 135042 285126 135084 285362
rect 113052 285084 135084 285126
rect 351700 285362 353860 285404
rect 351700 285126 351742 285362
rect 351978 285126 353582 285362
rect 353818 285126 353860 285362
rect 351700 285084 353860 285126
rect 0 284524 444740 284566
rect 0 284288 122 284524
rect 358 284288 442 284524
rect 678 284288 762 284524
rect 998 284288 1082 284524
rect 1318 284288 1402 284524
rect 1638 284288 1722 284524
rect 1958 284288 2042 284524
rect 2278 284288 2362 284524
rect 2598 284288 2682 284524
rect 2918 284288 3002 284524
rect 3238 284288 3322 284524
rect 3558 284288 3642 284524
rect 3878 284288 104506 284524
rect 104742 284288 198506 284524
rect 198742 284288 292506 284524
rect 292742 284288 440862 284524
rect 441098 284288 441182 284524
rect 441418 284288 441502 284524
rect 441738 284288 441822 284524
rect 442058 284288 442142 284524
rect 442378 284288 442462 284524
rect 442698 284288 442782 284524
rect 443018 284288 443102 284524
rect 443338 284288 443422 284524
rect 443658 284288 443742 284524
rect 443978 284288 444062 284524
rect 444298 284288 444382 284524
rect 444618 284288 444740 284524
rect 0 284246 444740 284288
rect 104404 283562 104724 283604
rect 104404 283326 104446 283562
rect 104682 283326 104724 283562
rect 104404 282684 104724 283326
rect 84348 282642 104724 282684
rect 84348 282406 84390 282642
rect 84626 282406 104724 282642
rect 84348 282364 104724 282406
rect 0 269206 444740 269248
rect 0 268970 5122 269206
rect 5358 268970 5442 269206
rect 5678 268970 5762 269206
rect 5998 268970 6082 269206
rect 6318 268970 6402 269206
rect 6638 268970 6722 269206
rect 6958 268970 7042 269206
rect 7278 268970 7362 269206
rect 7598 268970 7682 269206
rect 7918 268970 8002 269206
rect 8238 268970 8322 269206
rect 8558 268970 8642 269206
rect 8878 268970 435862 269206
rect 436098 268970 436182 269206
rect 436418 268970 436502 269206
rect 436738 268970 436822 269206
rect 437058 268970 437142 269206
rect 437378 268970 437462 269206
rect 437698 268970 437782 269206
rect 438018 268970 438102 269206
rect 438338 268970 438422 269206
rect 438658 268970 438742 269206
rect 438978 268970 439062 269206
rect 439298 268970 439382 269206
rect 439618 268970 444740 269206
rect 0 268928 444740 268970
rect 229708 264004 232236 264324
rect 229708 263644 230028 264004
rect 224740 263602 230028 263644
rect 224740 263366 224782 263602
rect 225018 263366 230028 263602
rect 224740 263324 230028 263366
rect 231916 263644 232236 264004
rect 234676 264004 241804 264324
rect 234676 263644 234996 264004
rect 231916 263324 234996 263644
rect 241484 263644 241804 264004
rect 241484 263602 245300 263644
rect 241484 263366 245022 263602
rect 245258 263366 245300 263602
rect 241484 263324 245300 263366
rect 154452 262922 161948 262964
rect 154452 262686 154494 262922
rect 154730 262686 161948 262922
rect 154452 262644 161948 262686
rect 148932 262242 149252 262284
rect 148932 262006 148974 262242
rect 149210 262006 149252 262242
rect 48836 259522 75284 259564
rect 48836 259286 48878 259522
rect 49114 259286 75006 259522
rect 75242 259286 75284 259522
rect 48836 259244 75284 259286
rect 63556 258162 76204 258204
rect 63556 257926 75926 258162
rect 76162 257926 76204 258162
rect 63556 257884 76204 257926
rect 63556 256164 63876 257884
rect 148932 256844 149252 262006
rect 161628 260924 161948 262644
rect 259516 262644 269404 262964
rect 167700 262242 184028 262284
rect 167700 262006 183750 262242
rect 183986 262006 184028 262242
rect 167700 261964 184028 262006
rect 212412 262242 215492 262284
rect 212412 262006 212454 262242
rect 212690 262006 215492 262242
rect 212412 261964 215492 262006
rect 167700 261604 168020 261964
rect 164388 261284 168020 261604
rect 164388 260924 164708 261284
rect 215172 260924 215492 261964
rect 241300 262242 241620 262284
rect 241300 262006 241342 262242
rect 241578 262006 241620 262242
rect 161628 260604 164708 260924
rect 193092 260882 203348 260924
rect 193092 260646 193134 260882
rect 193370 260646 203070 260882
rect 203306 260646 203348 260882
rect 193092 260604 203348 260646
rect 215172 260882 225060 260924
rect 215172 260646 224782 260882
rect 225018 260646 225060 260882
rect 215172 260604 225060 260646
rect 241300 259564 241620 262006
rect 247188 262242 248060 262284
rect 247188 262006 247782 262242
rect 248018 262006 248060 262242
rect 247188 261964 248060 262006
rect 251052 262242 251372 262284
rect 251052 262006 251094 262242
rect 251330 262006 251372 262242
rect 247188 259564 247508 261964
rect 251052 261604 251372 262006
rect 251052 261284 254316 261604
rect 251052 260604 251556 261284
rect 253996 260924 254316 261284
rect 259516 260924 259836 262644
rect 269084 261604 269404 262644
rect 269084 261562 279156 261604
rect 269084 261326 278878 261562
rect 279114 261326 279156 261562
rect 269084 261284 279156 261326
rect 288404 261562 298476 261604
rect 288404 261326 288446 261562
rect 288682 261326 298198 261562
rect 298434 261326 298476 261562
rect 288404 261284 298476 261326
rect 307724 261562 317796 261604
rect 307724 261326 307766 261562
rect 308002 261326 317518 261562
rect 317754 261326 317796 261562
rect 307724 261284 317796 261326
rect 327044 261562 337116 261604
rect 327044 261326 327086 261562
rect 327322 261326 337116 261562
rect 327044 261284 337116 261326
rect 253996 260604 259836 260924
rect 336796 260244 337116 261284
rect 346364 261562 356436 261604
rect 346364 261326 356158 261562
rect 356394 261326 356436 261562
rect 346364 261284 356436 261326
rect 346364 260244 346684 261284
rect 336796 259924 346684 260244
rect 237988 259522 241620 259564
rect 237988 259286 238030 259522
rect 238266 259286 241620 259522
rect 237988 259244 241620 259286
rect 242220 259244 247508 259564
rect 143964 256802 149252 256844
rect 143964 256566 144006 256802
rect 144242 256566 149252 256802
rect 143964 256524 149252 256566
rect 48836 256122 63876 256164
rect 48836 255886 48878 256122
rect 49114 255886 63876 256122
rect 48836 255844 63876 255886
rect 242220 255484 242540 259244
rect 237620 255442 242540 255484
rect 237620 255206 237662 255442
rect 237898 255206 242540 255442
rect 237620 255164 242540 255206
rect 74044 254762 75652 254804
rect 74044 254526 74086 254762
rect 74322 254526 75374 254762
rect 75610 254526 75652 254762
rect 74044 254484 75652 254526
rect 0 253888 444740 253930
rect 0 253652 122 253888
rect 358 253652 442 253888
rect 678 253652 762 253888
rect 998 253652 1082 253888
rect 1318 253652 1402 253888
rect 1638 253652 1722 253888
rect 1958 253652 2042 253888
rect 2278 253652 2362 253888
rect 2598 253652 2682 253888
rect 2918 253652 3002 253888
rect 3238 253652 3322 253888
rect 3558 253652 3642 253888
rect 3878 253652 440862 253888
rect 441098 253652 441182 253888
rect 441418 253652 441502 253888
rect 441738 253652 441822 253888
rect 442058 253652 442142 253888
rect 442378 253652 442462 253888
rect 442698 253652 442782 253888
rect 443018 253652 443102 253888
rect 443338 253652 443422 253888
rect 443658 253652 443742 253888
rect 443978 253652 444062 253888
rect 444298 253652 444382 253888
rect 444618 253652 444740 253888
rect 0 253610 444740 253652
rect 74044 252042 75652 252084
rect 74044 251806 75374 252042
rect 75610 251806 75652 252042
rect 74044 251764 75652 251806
rect 74044 251404 74364 251764
rect 73860 251084 74364 251404
rect 73860 250044 74180 251084
rect 63556 249724 74180 250044
rect 63556 249364 63876 249724
rect 48836 249322 63876 249364
rect 48836 249086 48878 249322
rect 49114 249086 63876 249322
rect 48836 249044 63876 249086
rect 237620 248642 247692 248684
rect 237620 248406 237662 248642
rect 237898 248406 247692 248642
rect 237620 248364 247692 248406
rect 143964 247962 149252 248004
rect 143964 247726 144006 247962
rect 144242 247726 149252 247962
rect 143964 247684 149252 247726
rect 148932 245964 149252 247684
rect 237988 246602 242908 246644
rect 237988 246366 238030 246602
rect 238266 246366 242908 246602
rect 237988 246324 242908 246366
rect 242588 245964 242908 246324
rect 74228 245922 74548 245964
rect 74228 245686 74270 245922
rect 74506 245686 74548 245922
rect 74228 244604 74548 245686
rect 142860 245922 149252 245964
rect 142860 245686 142902 245922
rect 143138 245686 149252 245922
rect 142860 245644 149252 245686
rect 237988 245922 242908 245964
rect 237988 245686 238030 245922
rect 238266 245686 242908 245922
rect 237988 245644 242908 245686
rect 74044 244562 74548 244604
rect 74044 244326 74086 244562
rect 74322 244326 74548 244562
rect 74044 244284 74548 244326
rect 141020 244562 153484 244604
rect 141020 244326 141062 244562
rect 141298 244326 153484 244562
rect 141020 244284 153484 244326
rect 58772 243604 65164 243924
rect 58772 243244 59092 243604
rect 53252 242924 59092 243244
rect 53252 242564 53572 242924
rect 46812 242522 53572 242564
rect 46812 242286 46854 242522
rect 47090 242286 53572 242522
rect 46812 242244 53572 242286
rect 63372 242244 63876 243604
rect 64844 242564 65164 243604
rect 71836 243882 77124 243924
rect 71836 243646 76846 243882
rect 77082 243646 77124 243882
rect 71836 243604 77124 243646
rect 71836 242564 72156 243604
rect 64844 242244 72156 242564
rect 72940 242522 76756 242564
rect 72940 242286 76478 242522
rect 76714 242286 76756 242522
rect 72940 242244 76756 242286
rect 72940 241884 73260 242244
rect 53988 241564 62588 241884
rect 53988 241204 54308 241564
rect 49020 241162 54308 241204
rect 49020 240926 49062 241162
rect 49298 240926 54308 241162
rect 49020 240884 54308 240926
rect 62268 240524 62588 241564
rect 63556 241564 71972 241884
rect 63556 240524 63876 241564
rect 62268 240204 63876 240524
rect 71652 240524 71972 241564
rect 72572 241564 73260 241884
rect 95204 241564 96260 241884
rect 72572 241204 72892 241564
rect 95204 241204 95524 241564
rect 72388 240884 72892 241204
rect 76436 241162 84668 241204
rect 76436 240926 76478 241162
rect 76714 240926 84390 241162
rect 84626 240926 84668 241162
rect 76436 240884 84668 240926
rect 93732 241162 95524 241204
rect 93732 240926 93774 241162
rect 94010 240926 95524 241162
rect 93732 240884 95524 240926
rect 95940 241162 96260 241564
rect 95940 240926 95982 241162
rect 96218 240926 96260 241162
rect 95940 240884 96260 240926
rect 128508 241842 137108 241884
rect 128508 241606 136830 241842
rect 137066 241606 137108 241842
rect 128508 241564 137108 241606
rect 72388 240524 72708 240884
rect 128508 240524 128828 241564
rect 71652 240204 72708 240524
rect 73492 240482 76204 240524
rect 73492 240246 75926 240482
rect 76162 240246 76204 240482
rect 73492 240204 76204 240246
rect 104772 240482 128828 240524
rect 104772 240246 104814 240482
rect 105050 240246 128828 240482
rect 104772 240204 128828 240246
rect 153164 240524 153484 244284
rect 158500 242244 161764 242564
rect 158500 240524 158820 242244
rect 153164 240204 158820 240524
rect 73492 239844 73812 240204
rect 161444 239844 161764 242244
rect 168068 240482 196356 240524
rect 168068 240246 168110 240482
rect 168346 240246 196078 240482
rect 196314 240246 196356 240482
rect 168068 240204 196356 240246
rect 247372 239844 247692 248364
rect 261908 240482 305284 240524
rect 261908 240246 261950 240482
rect 262186 240246 305006 240482
rect 305242 240246 305284 240482
rect 261908 240204 305284 240246
rect 49020 239802 73812 239844
rect 49020 239566 49062 239802
rect 49298 239566 73812 239802
rect 49020 239524 73812 239566
rect 76804 239802 141340 239844
rect 76804 239566 76846 239802
rect 77082 239566 95062 239802
rect 95298 239566 138302 239802
rect 138538 239566 141062 239802
rect 141298 239566 141340 239802
rect 76804 239524 141340 239566
rect 161444 239802 188076 239844
rect 161444 239566 187798 239802
rect 188034 239566 188076 239802
rect 161444 239524 188076 239566
rect 237620 239802 247692 239844
rect 237620 239566 237662 239802
rect 237898 239566 247692 239802
rect 237620 239524 247692 239566
rect 295396 239802 324788 239844
rect 295396 239566 295438 239802
rect 295674 239566 324510 239802
rect 324746 239566 324788 239802
rect 295396 239524 324788 239566
rect 0 238570 444740 238612
rect 0 238334 5122 238570
rect 5358 238334 5442 238570
rect 5678 238334 5762 238570
rect 5998 238334 6082 238570
rect 6318 238334 6402 238570
rect 6638 238334 6722 238570
rect 6958 238334 7042 238570
rect 7278 238334 7362 238570
rect 7598 238334 7682 238570
rect 7918 238334 8002 238570
rect 8238 238334 8322 238570
rect 8558 238334 8642 238570
rect 8878 238334 435862 238570
rect 436098 238334 436182 238570
rect 436418 238334 436502 238570
rect 436738 238334 436822 238570
rect 437058 238334 437142 238570
rect 437378 238334 437462 238570
rect 437698 238334 437782 238570
rect 438018 238334 438102 238570
rect 438338 238334 438422 238570
rect 438658 238334 438742 238570
rect 438978 238334 439062 238570
rect 439298 238334 439382 238570
rect 439618 238334 444740 238570
rect 0 238292 444740 238334
rect 99988 237762 109508 237804
rect 99988 237526 100030 237762
rect 100266 237526 109508 237762
rect 99988 237484 109508 237526
rect 81220 237082 90188 237124
rect 81220 236846 81262 237082
rect 81498 236846 89910 237082
rect 90146 236846 90188 237082
rect 81220 236804 90188 236846
rect 109188 236444 109508 237484
rect 135500 237762 147964 237804
rect 135500 237526 147686 237762
rect 147922 237526 147964 237762
rect 135500 237484 147964 237526
rect 237620 237762 247324 237804
rect 237620 237526 237662 237762
rect 237898 237526 247046 237762
rect 247282 237526 247324 237762
rect 237620 237484 247324 237526
rect 261540 237762 264988 237804
rect 261540 237526 261582 237762
rect 261818 237526 264710 237762
rect 264946 237526 264988 237762
rect 261540 237484 264988 237526
rect 135500 236444 135820 237484
rect 142860 237082 145388 237124
rect 142860 236846 142902 237082
rect 143138 236846 145110 237082
rect 145346 236846 145388 237082
rect 142860 236804 145388 236846
rect 145804 237082 148884 237124
rect 145804 236846 145846 237082
rect 146082 236846 148606 237082
rect 148842 236846 148884 237082
rect 145804 236804 148884 236846
rect 176900 237082 186788 237124
rect 176900 236846 176942 237082
rect 177178 236846 186510 237082
rect 186746 236846 186788 237082
rect 176900 236804 186788 236846
rect 231732 237082 241988 237124
rect 231732 236846 231774 237082
rect 232010 236846 238030 237082
rect 238266 236846 241988 237082
rect 231732 236804 241988 236846
rect 273684 237082 290196 237124
rect 273684 236846 273726 237082
rect 273962 236846 289918 237082
rect 290154 236846 290196 237082
rect 273684 236804 290196 236846
rect 241668 236444 241988 236804
rect 74780 236402 105276 236444
rect 74780 236166 104998 236402
rect 105234 236166 105276 236402
rect 74780 236124 105276 236166
rect 109188 236124 118892 236444
rect 133844 236402 136556 236444
rect 133844 236166 133886 236402
rect 134122 236166 136278 236402
rect 136514 236166 136556 236402
rect 133844 236124 136556 236166
rect 156660 236402 203348 236444
rect 156660 236166 156702 236402
rect 156938 236166 168846 236402
rect 169082 236166 203070 236402
rect 203306 236166 203348 236402
rect 156660 236124 203348 236166
rect 241668 236402 244748 236444
rect 241668 236166 244102 236402
rect 244338 236308 244748 236402
rect 247004 236402 287068 236444
rect 244338 236166 245300 236308
rect 241668 236124 245300 236166
rect 247004 236166 247046 236402
rect 247282 236166 286790 236402
rect 287026 236166 287068 236402
rect 247004 236124 287068 236166
rect 74780 235722 75100 236124
rect 118572 235764 118892 236124
rect 244428 235988 245300 236124
rect 244980 235764 245300 235988
rect 74780 235486 74822 235722
rect 75058 235486 75100 235722
rect 74780 235444 75100 235486
rect 76252 235722 116316 235764
rect 76252 235486 76294 235722
rect 76530 235486 116038 235722
rect 116274 235486 116316 235722
rect 76252 235444 116316 235486
rect 118572 235722 124596 235764
rect 118572 235486 124318 235722
rect 124554 235486 124596 235722
rect 118572 235444 124596 235486
rect 148932 235722 192308 235764
rect 148932 235486 192030 235722
rect 192266 235486 192308 235722
rect 148932 235444 192308 235486
rect 244980 235722 295716 235764
rect 244980 235486 295438 235722
rect 295674 235486 295716 235722
rect 244980 235444 295716 235486
rect 148932 235084 149252 235444
rect 137156 235042 149252 235084
rect 137156 234806 137198 235042
rect 137434 234806 148054 235042
rect 148290 234806 149252 235042
rect 137156 234764 149252 234806
rect 158684 235042 207396 235084
rect 158684 234806 158726 235042
rect 158962 234806 168478 235042
rect 168714 234806 207118 235042
rect 207354 234806 207396 235042
rect 158684 234764 207396 234806
rect 231180 235042 245668 235084
rect 231180 234806 231222 235042
rect 231458 234806 245390 235042
rect 245626 234806 245668 235042
rect 231180 234764 245668 234806
rect 246084 235042 301236 235084
rect 246084 234806 246126 235042
rect 246362 234806 262318 235042
rect 262554 234806 300958 235042
rect 301194 234806 301236 235042
rect 246084 234764 301236 234806
rect 137524 234362 137844 234404
rect 137524 234126 137566 234362
rect 137802 234126 137844 234362
rect 137524 233724 137844 234126
rect 148564 234362 152196 234404
rect 148564 234126 151918 234362
rect 152154 234126 152196 234362
rect 148564 234084 152196 234126
rect 230628 234362 245668 234404
rect 230628 234126 230670 234362
rect 230906 234126 245390 234362
rect 245626 234126 245668 234362
rect 230628 234084 245668 234126
rect 249764 234362 283388 234404
rect 249764 234126 249806 234362
rect 250042 234126 283110 234362
rect 283346 234126 283388 234362
rect 249764 234084 283388 234126
rect 148564 233724 148884 234084
rect 137524 233404 148884 233724
rect 0 223252 444740 223294
rect 0 223016 122 223252
rect 358 223016 442 223252
rect 678 223016 762 223252
rect 998 223016 1082 223252
rect 1318 223016 1402 223252
rect 1638 223016 1722 223252
rect 1958 223016 2042 223252
rect 2278 223016 2362 223252
rect 2598 223016 2682 223252
rect 2918 223016 3002 223252
rect 3238 223016 3322 223252
rect 3558 223016 3642 223252
rect 3878 223016 104506 223252
rect 104742 223016 198506 223252
rect 198742 223016 292506 223252
rect 292742 223016 380882 223252
rect 381118 223016 440862 223252
rect 441098 223016 441182 223252
rect 441418 223016 441502 223252
rect 441738 223016 441822 223252
rect 442058 223016 442142 223252
rect 442378 223016 442462 223252
rect 442698 223016 442782 223252
rect 443018 223016 443102 223252
rect 443338 223016 443422 223252
rect 443658 223016 443742 223252
rect 443978 223016 444062 223252
rect 444298 223016 444382 223252
rect 444618 223016 444740 223252
rect 0 222974 444740 223016
rect 292452 217404 292956 218084
rect 283068 217084 292956 217404
rect 283068 216724 283388 217084
rect 242588 216682 259100 216724
rect 242588 216446 242630 216682
rect 242866 216446 258822 216682
rect 259058 216446 259100 216682
rect 242588 216404 259100 216446
rect 272580 216682 283388 216724
rect 272580 216446 272622 216682
rect 272858 216446 283388 216682
rect 272580 216404 283388 216446
rect 292636 216724 292956 217084
rect 311956 218042 322948 218084
rect 311956 217806 322670 218042
rect 322906 217806 322948 218042
rect 311956 217764 322948 217806
rect 311956 216724 312276 217764
rect 292636 216404 312276 216724
rect 336612 216682 352940 216724
rect 336612 216446 336654 216682
rect 336890 216446 352662 216682
rect 352898 216446 352940 216682
rect 336612 216404 352940 216446
rect 357404 216002 406116 216044
rect 357404 215766 357446 216002
rect 357682 215766 405838 216002
rect 406074 215766 406116 216002
rect 357404 215724 406116 215766
rect 178556 214642 182924 214684
rect 178556 214406 178598 214642
rect 178834 214406 182924 214642
rect 178556 214364 182924 214406
rect 182604 211284 182924 214364
rect 178556 211242 182924 211284
rect 178556 211006 178598 211242
rect 178834 211006 182924 211242
rect 178556 210964 182924 211006
rect 0 207934 444740 207976
rect 0 207698 5122 207934
rect 5358 207698 5442 207934
rect 5678 207698 5762 207934
rect 5998 207698 6082 207934
rect 6318 207698 6402 207934
rect 6638 207698 6722 207934
rect 6958 207698 7042 207934
rect 7278 207698 7362 207934
rect 7598 207698 7682 207934
rect 7918 207698 8002 207934
rect 8238 207698 8322 207934
rect 8558 207698 8642 207934
rect 8878 207698 89146 207934
rect 89382 207698 183146 207934
rect 183382 207698 277146 207934
rect 277382 207698 435862 207934
rect 436098 207698 436182 207934
rect 436418 207698 436502 207934
rect 436738 207698 436822 207934
rect 437058 207698 437142 207934
rect 437378 207698 437462 207934
rect 437698 207698 437782 207934
rect 438018 207698 438102 207934
rect 438338 207698 438422 207934
rect 438658 207698 438742 207934
rect 438978 207698 439062 207934
rect 439298 207698 439382 207934
rect 439618 207698 444740 207934
rect 0 207656 444740 207698
rect 93916 206204 109140 206524
rect 93916 204484 94236 206204
rect 108820 205164 109140 206204
rect 115996 206204 119076 206524
rect 115996 205844 116316 206204
rect 115444 205524 116316 205844
rect 118756 205844 119076 206204
rect 120780 206204 128644 206524
rect 120780 205844 121100 206204
rect 118756 205524 121100 205844
rect 115444 205164 115764 205524
rect 108820 204844 115764 205164
rect 128324 205164 128644 206204
rect 128324 205122 134900 205164
rect 128324 204886 134622 205122
rect 134858 204886 134900 205122
rect 128324 204844 134900 204886
rect 84532 204442 94236 204484
rect 84532 204206 84574 204442
rect 84810 204206 94236 204442
rect 84532 204164 94236 204206
rect 239460 204442 322948 204484
rect 239460 204206 239502 204442
rect 239738 204206 322670 204442
rect 322906 204206 322948 204442
rect 239460 204164 322948 204206
rect 136788 201042 322948 201084
rect 136788 200806 136830 201042
rect 137066 200806 228646 201042
rect 228882 200806 322670 201042
rect 322906 200806 322948 201042
rect 136788 200764 322948 200806
rect 136788 199002 138396 199044
rect 136788 198766 136830 199002
rect 137066 198766 138396 199002
rect 136788 198724 138396 198766
rect 138076 197684 138396 198724
rect 154452 198724 157532 199044
rect 154452 198364 154772 198724
rect 145068 198044 154772 198364
rect 145068 197684 145388 198044
rect 138076 197364 145388 197684
rect 157212 197684 157532 198724
rect 212412 198724 215492 199044
rect 212412 198364 212732 198724
rect 176532 198322 176852 198364
rect 176532 198086 176574 198322
rect 176810 198086 176852 198322
rect 176532 197684 176852 198086
rect 193092 198044 195988 198364
rect 157212 197642 164708 197684
rect 157212 197406 164430 197642
rect 164666 197406 164708 197642
rect 157212 197364 164708 197406
rect 176532 197364 184028 197684
rect 183708 196324 184028 197364
rect 193092 196324 193412 198044
rect 195668 197684 195988 198044
rect 203028 198044 212732 198364
rect 203028 197684 203348 198044
rect 195668 197364 203348 197684
rect 215172 197684 215492 198724
rect 222348 199002 234812 199044
rect 222348 198766 230670 199002
rect 230906 198766 234812 199002
rect 222348 198724 234812 198766
rect 222348 197684 222668 198724
rect 215172 197364 222668 197684
rect 234492 197684 234812 198724
rect 251052 198724 254132 199044
rect 251052 197684 251372 198724
rect 234492 197364 251372 197684
rect 253812 197684 254132 198724
rect 289692 198724 292772 199044
rect 270372 198322 273452 198364
rect 270372 198086 270414 198322
rect 270650 198086 273452 198322
rect 270372 198044 273452 198086
rect 273132 197684 273452 198044
rect 253812 197642 261308 197684
rect 253812 197406 261030 197642
rect 261266 197406 261308 197642
rect 253812 197364 261308 197406
rect 273132 197364 280628 197684
rect 183708 196004 193412 196324
rect 280308 196324 280628 197364
rect 289692 196324 290012 198724
rect 292452 197684 292772 198724
rect 309012 198724 312092 199044
rect 292452 197364 299948 197684
rect 280308 196004 290012 196324
rect 299628 196324 299948 197364
rect 309012 196324 309332 198724
rect 311772 197684 312092 198724
rect 318948 199002 322948 199044
rect 318948 198766 322670 199002
rect 322906 198766 322948 199002
rect 318948 198724 322948 198766
rect 318948 197684 319268 198724
rect 311772 197364 319268 197684
rect 299628 196004 309332 196324
rect 178556 195602 183476 195644
rect 178556 195366 178598 195602
rect 178834 195366 183476 195602
rect 178556 195324 183476 195366
rect 183156 194964 183476 195324
rect 178556 194922 183476 194964
rect 178556 194686 178598 194922
rect 178834 194686 183476 194922
rect 178556 194644 183476 194686
rect 137892 194242 322948 194284
rect 137892 194006 137934 194242
rect 138170 194006 230670 194242
rect 230906 194006 322670 194242
rect 322906 194006 322948 194242
rect 137892 193964 322948 194006
rect 0 192616 444740 192658
rect 0 192380 122 192616
rect 358 192380 442 192616
rect 678 192380 762 192616
rect 998 192380 1082 192616
rect 1318 192380 1402 192616
rect 1638 192380 1722 192616
rect 1958 192380 2042 192616
rect 2278 192380 2362 192616
rect 2598 192380 2682 192616
rect 2918 192380 3002 192616
rect 3238 192380 3322 192616
rect 3558 192380 3642 192616
rect 3878 192380 104506 192616
rect 104742 192380 198506 192616
rect 198742 192380 292506 192616
rect 292742 192380 440862 192616
rect 441098 192380 441182 192616
rect 441418 192380 441502 192616
rect 441738 192380 441822 192616
rect 442058 192380 442142 192616
rect 442378 192380 442462 192616
rect 442698 192380 442782 192616
rect 443018 192380 443102 192616
rect 443338 192380 443422 192616
rect 443658 192380 443742 192616
rect 443978 192380 444062 192616
rect 444298 192380 444382 192616
rect 444618 192380 444740 192616
rect 0 192338 444740 192380
rect 178556 186082 183476 186124
rect 178556 185846 178598 186082
rect 178834 185846 183476 186082
rect 178556 185804 183476 185846
rect 183156 185444 183476 185804
rect 182972 185124 183476 185444
rect 182972 182724 183292 185124
rect 302204 183404 302708 184084
rect 178188 182682 183292 182724
rect 178188 182446 178230 182682
rect 178466 182446 183292 182682
rect 178188 182404 183292 182446
rect 195852 182044 196356 183404
rect 288404 183084 302708 183404
rect 271292 182682 280444 182724
rect 271292 182446 271334 182682
rect 271570 182446 280444 182682
rect 271292 182404 280444 182446
rect 280124 182044 280444 182404
rect 186468 181724 219724 182044
rect 280124 181724 287068 182044
rect 186468 181364 186788 181724
rect 183524 181044 186788 181364
rect 219404 181364 219724 181724
rect 219404 181322 229108 181364
rect 219404 181086 228830 181322
rect 229066 181086 229108 181322
rect 219404 181044 229108 181086
rect 280124 181044 283204 181364
rect 183524 180004 183844 181044
rect 280124 180004 280444 181044
rect 282884 180684 283204 181044
rect 282884 180364 286332 180684
rect 174692 179962 183844 180004
rect 174692 179726 174734 179962
rect 174970 179726 183844 179962
rect 174692 179684 183844 179726
rect 271292 179962 280444 180004
rect 271292 179726 271334 179962
rect 271570 179726 280444 179962
rect 271292 179684 280444 179726
rect 286012 179282 286332 180364
rect 286748 180004 287068 181724
rect 286748 179684 287620 180004
rect 286012 179046 286054 179282
rect 286290 179046 286332 179282
rect 286012 179004 286332 179046
rect 287300 179282 287620 179684
rect 287300 179046 287342 179282
rect 287578 179046 287620 179282
rect 287300 179004 287620 179046
rect 288404 179282 288724 183084
rect 302388 182724 302708 183084
rect 316188 183362 323132 183404
rect 316188 183126 322854 183362
rect 323090 183126 323132 183362
rect 316188 183084 323132 183126
rect 302388 182404 311356 182724
rect 311036 180004 311356 182404
rect 316188 182044 316508 183084
rect 288404 179046 288446 179282
rect 288682 179046 288724 179282
rect 288404 179004 288724 179046
rect 289324 179684 310068 180004
rect 289324 179282 289644 179684
rect 289324 179046 289366 179282
rect 289602 179046 289644 179282
rect 289324 179004 289644 179046
rect 309748 179282 310068 179684
rect 309748 179046 309790 179282
rect 310026 179046 310068 179282
rect 309748 179004 310068 179046
rect 310852 179684 311356 180004
rect 311772 181724 316508 182044
rect 316924 182002 323132 182044
rect 316924 181766 322854 182002
rect 323090 181766 323132 182002
rect 316924 181724 323132 181766
rect 310852 179282 311172 179684
rect 310852 179046 310894 179282
rect 311130 179046 311172 179282
rect 310852 179004 311172 179046
rect 311772 179282 312092 181724
rect 311772 179046 311814 179282
rect 312050 179046 312092 179282
rect 311772 179004 312092 179046
rect 316924 179282 317244 181724
rect 316924 179046 316966 179282
rect 317202 179046 317244 179282
rect 316924 179004 317244 179046
rect 0 177298 444740 177340
rect 0 177062 5122 177298
rect 5358 177062 5442 177298
rect 5678 177062 5762 177298
rect 5998 177062 6082 177298
rect 6318 177062 6402 177298
rect 6638 177062 6722 177298
rect 6958 177062 7042 177298
rect 7278 177062 7362 177298
rect 7598 177062 7682 177298
rect 7918 177062 8002 177298
rect 8238 177062 8322 177298
rect 8558 177062 8642 177298
rect 8878 177062 435862 177298
rect 436098 177062 436182 177298
rect 436418 177062 436502 177298
rect 436738 177062 436822 177298
rect 437058 177062 437142 177298
rect 437378 177062 437462 177298
rect 437698 177062 437782 177298
rect 438018 177062 438102 177298
rect 438338 177062 438422 177298
rect 438658 177062 438742 177298
rect 438978 177062 439062 177298
rect 439298 177062 439382 177298
rect 439618 177062 444740 177298
rect 0 177020 444740 177062
rect 241668 169082 244196 169124
rect 241668 168846 241710 169082
rect 241946 168846 244196 169082
rect 241668 168804 244196 168846
rect 241852 168402 242540 168444
rect 241852 168166 242262 168402
rect 242498 168166 242540 168402
rect 241852 168124 242540 168166
rect 243140 168402 243460 168444
rect 243140 168166 243182 168402
rect 243418 168166 243460 168402
rect 241852 165724 242172 168124
rect 237988 165682 242172 165724
rect 237988 165446 238030 165682
rect 238266 165446 242172 165682
rect 237988 165404 242172 165446
rect 243140 165044 243460 168166
rect 75332 165002 76940 165044
rect 75332 164766 75374 165002
rect 75610 164766 76662 165002
rect 76898 164766 76940 165002
rect 75332 164724 76940 164766
rect 237620 165002 243460 165044
rect 237620 164766 237662 165002
rect 237898 164766 243460 165002
rect 237620 164724 243460 164766
rect 243876 164364 244196 168804
rect 237252 164322 244196 164364
rect 237252 164086 237294 164322
rect 237530 164086 244196 164322
rect 237252 164044 244196 164086
rect 48836 162962 76940 163004
rect 48836 162726 48878 162962
rect 49114 162726 76662 162962
rect 76898 162726 76940 162962
rect 48836 162684 76940 162726
rect 0 161980 444740 162022
rect 0 161744 122 161980
rect 358 161744 442 161980
rect 678 161744 762 161980
rect 998 161744 1082 161980
rect 1318 161744 1402 161980
rect 1638 161744 1722 161980
rect 1958 161744 2042 161980
rect 2278 161744 2362 161980
rect 2598 161744 2682 161980
rect 2918 161744 3002 161980
rect 3238 161744 3322 161980
rect 3558 161744 3642 161980
rect 3878 161744 440862 161980
rect 441098 161744 441182 161980
rect 441418 161744 441502 161980
rect 441738 161744 441822 161980
rect 442058 161744 442142 161980
rect 442378 161744 442462 161980
rect 442698 161744 442782 161980
rect 443018 161744 443102 161980
rect 443338 161744 443422 161980
rect 443658 161744 443742 161980
rect 443978 161744 444062 161980
rect 444298 161744 444382 161980
rect 444618 161744 444740 161980
rect 0 161702 444740 161744
rect 143964 160922 148700 160964
rect 143964 160686 144006 160922
rect 144242 160686 148700 160922
rect 143964 160644 148700 160686
rect 237252 160922 247324 160964
rect 237252 160686 237294 160922
rect 237530 160686 247324 160922
rect 237252 160644 247324 160686
rect 75332 160242 76940 160284
rect 75332 160006 75374 160242
rect 75610 160006 76662 160242
rect 76898 160006 76940 160242
rect 75332 159964 76940 160006
rect 49020 158202 72892 158244
rect 49020 157966 49062 158202
rect 49298 157966 72892 158202
rect 49020 157924 72892 157966
rect 72572 157564 72892 157924
rect 75148 158202 75468 158244
rect 75148 157966 75190 158202
rect 75426 157966 75468 158202
rect 75148 157564 75468 157966
rect 72572 157244 76572 157564
rect 74044 156842 75652 156884
rect 74044 156606 74086 156842
rect 74322 156606 75374 156842
rect 75610 156606 75652 156842
rect 74044 156564 75652 156606
rect 76252 156842 76572 157244
rect 76252 156606 76294 156842
rect 76530 156606 76572 156842
rect 76252 156564 76572 156606
rect 49020 155482 76204 155524
rect 49020 155246 49062 155482
rect 49298 155246 76204 155482
rect 49020 155204 76204 155246
rect 75700 154844 76204 155204
rect 75700 154802 76940 154844
rect 75700 154566 76662 154802
rect 76898 154566 76940 154802
rect 75700 154524 76940 154566
rect 75700 153484 76020 154524
rect 75700 153442 77308 153484
rect 75700 153206 77030 153442
rect 77266 153206 77308 153442
rect 75700 153164 77308 153206
rect 49020 152762 74548 152804
rect 49020 152526 49062 152762
rect 49298 152526 74270 152762
rect 74506 152526 74548 152762
rect 49020 152484 74548 152526
rect 148380 151444 148700 160644
rect 237988 157522 242540 157564
rect 237988 157286 238030 157522
rect 238266 157286 242540 157522
rect 237988 157244 242540 157286
rect 237620 156842 241804 156884
rect 237620 156606 237662 156842
rect 237898 156606 241804 156842
rect 237620 156564 241804 156606
rect 241484 153484 241804 156564
rect 236700 153442 241804 153484
rect 236700 153206 236742 153442
rect 236978 153206 241804 153442
rect 236700 153164 241804 153206
rect 147828 151124 148700 151444
rect 147828 150764 148148 151124
rect 143964 150722 148148 150764
rect 143964 150486 144006 150722
rect 144242 150486 148148 150722
rect 143964 150444 148148 150486
rect 242220 148724 242540 157244
rect 49020 148682 74916 148724
rect 49020 148446 49062 148682
rect 49298 148446 74638 148682
rect 74874 148446 74916 148682
rect 49020 148404 74916 148446
rect 237252 148682 242540 148724
rect 237252 148446 237294 148682
rect 237530 148446 242540 148682
rect 237252 148404 242540 148446
rect 247004 147364 247324 160644
rect 237436 147322 247324 147364
rect 237436 147086 237478 147322
rect 237714 147086 247324 147322
rect 237436 147044 247324 147086
rect 0 146662 444740 146704
rect 0 146426 5122 146662
rect 5358 146426 5442 146662
rect 5678 146426 5762 146662
rect 5998 146426 6082 146662
rect 6318 146426 6402 146662
rect 6638 146426 6722 146662
rect 6958 146426 7042 146662
rect 7278 146426 7362 146662
rect 7598 146426 7682 146662
rect 7918 146426 8002 146662
rect 8238 146426 8322 146662
rect 8558 146426 8642 146662
rect 8878 146426 435862 146662
rect 436098 146426 436182 146662
rect 436418 146426 436502 146662
rect 436738 146426 436822 146662
rect 437058 146426 437142 146662
rect 437378 146426 437462 146662
rect 437698 146426 437782 146662
rect 438018 146426 438102 146662
rect 438338 146426 438422 146662
rect 438658 146426 438742 146662
rect 438978 146426 439062 146662
rect 439298 146426 439382 146662
rect 439618 146426 444740 146662
rect 0 146384 444740 146426
rect 49020 145962 76756 146004
rect 49020 145726 49062 145962
rect 49298 145726 74454 145962
rect 74690 145726 76478 145962
rect 76714 145726 76756 145962
rect 49020 145684 76756 145726
rect 74780 145282 77308 145324
rect 74780 145046 74822 145282
rect 75058 145046 77030 145282
rect 77266 145046 77308 145282
rect 74780 145004 77308 145046
rect 153348 145004 163052 145324
rect 169356 145282 176484 145324
rect 169356 145046 169398 145282
rect 169634 145046 176206 145282
rect 176442 145046 176484 145282
rect 169356 145004 176484 145046
rect 138076 144602 142628 144644
rect 138076 144366 142350 144602
rect 142586 144366 142628 144602
rect 138076 144324 142628 144366
rect 74780 143922 98468 143964
rect 74780 143686 74822 143922
rect 75058 143686 98190 143922
rect 98426 143686 98468 143922
rect 74780 143644 98468 143686
rect 138076 143284 138396 144324
rect 153348 143964 153668 145004
rect 75884 143242 110612 143284
rect 75884 143006 75926 143242
rect 76162 143006 110334 143242
rect 110570 143006 110612 143242
rect 75884 142964 110612 143006
rect 136788 143242 138396 143284
rect 136788 143006 136830 143242
rect 137066 143006 138396 143242
rect 136788 142964 138396 143006
rect 151692 143644 153668 143964
rect 151692 143242 152012 143644
rect 151692 143006 151734 143242
rect 151970 143006 152012 143242
rect 151692 142964 152012 143006
rect 162732 143284 163052 145004
rect 187020 144602 196356 144644
rect 187020 144366 187062 144602
rect 187298 144366 196078 144602
rect 196314 144366 196356 144602
rect 187020 144324 196356 144366
rect 162732 143242 169676 143284
rect 162732 143006 169398 143242
rect 169634 143006 169676 143242
rect 162732 142964 169676 143006
rect 170092 143242 210340 143284
rect 170092 143006 170134 143242
rect 170370 143006 210062 143242
rect 210298 143006 210340 143242
rect 170092 142964 210340 143006
rect 262828 143242 294428 143284
rect 262828 143006 262870 143242
rect 263106 143006 294150 143242
rect 294386 143006 294428 143242
rect 262828 142964 294428 143006
rect 78092 141882 105276 141924
rect 78092 141646 78134 141882
rect 78370 141646 104998 141882
rect 105234 141646 105276 141882
rect 78092 141604 105276 141646
rect 148932 141882 168572 141924
rect 148932 141646 168294 141882
rect 168530 141646 168572 141882
rect 148932 141604 168572 141646
rect 235964 141882 237940 141924
rect 235964 141646 236006 141882
rect 236242 141646 237662 141882
rect 237898 141646 237940 141882
rect 235964 141604 237940 141646
rect 256572 141882 290196 141924
rect 256572 141646 256614 141882
rect 256850 141646 289918 141882
rect 290154 141646 290196 141882
rect 256572 141604 290196 141646
rect 148932 141244 149252 141604
rect 137340 141202 149252 141244
rect 137340 140966 137382 141202
rect 137618 140966 148974 141202
rect 149210 140966 149252 141202
rect 137340 140924 149252 140966
rect 151876 141202 207396 141244
rect 151876 140966 168478 141202
rect 168714 140966 207118 141202
rect 207354 140966 207396 141202
rect 151876 140924 207396 140966
rect 258228 141202 273084 141244
rect 258228 140966 262318 141202
rect 262554 140966 273084 141202
rect 258228 140924 273084 140966
rect 151876 140564 152196 140924
rect 258228 140564 258548 140924
rect 137156 140522 152196 140564
rect 137156 140286 137198 140522
rect 137434 140286 151918 140522
rect 152154 140286 152196 140522
rect 137156 140244 152196 140286
rect 230628 140522 243276 140564
rect 230628 140286 230670 140522
rect 230906 140286 242998 140522
rect 243234 140286 243276 140522
rect 230628 140244 243276 140286
rect 251236 140522 258548 140564
rect 251236 140286 251278 140522
rect 251514 140286 258548 140522
rect 251236 140244 258548 140286
rect 272764 139884 273084 140924
rect 296684 141202 297188 141244
rect 296684 140966 296910 141202
rect 297146 140966 297188 141202
rect 296684 140924 297188 140966
rect 283068 140244 292772 140564
rect 283068 139884 283388 140244
rect 272764 139564 283388 139884
rect 292452 139884 292772 140244
rect 296684 139884 297004 140924
rect 292452 139564 297004 139884
rect 0 131344 444740 131386
rect 0 131108 122 131344
rect 358 131108 442 131344
rect 678 131108 762 131344
rect 998 131108 1082 131344
rect 1318 131108 1402 131344
rect 1638 131108 1722 131344
rect 1958 131108 2042 131344
rect 2278 131108 2362 131344
rect 2598 131108 2682 131344
rect 2918 131108 3002 131344
rect 3238 131108 3322 131344
rect 3558 131108 3642 131344
rect 3878 131108 440862 131344
rect 441098 131108 441182 131344
rect 441418 131108 441502 131344
rect 441738 131108 441822 131344
rect 442058 131108 442142 131344
rect 442378 131108 442462 131344
rect 442698 131108 442782 131344
rect 443018 131108 443102 131344
rect 443338 131108 443422 131344
rect 443658 131108 443742 131344
rect 443978 131108 444062 131344
rect 444298 131108 444382 131344
rect 444618 131108 444740 131344
rect 0 131066 444740 131108
rect 199164 131002 199484 131044
rect 199164 130766 199206 131002
rect 199442 130766 199484 131002
rect 178556 124882 181268 124924
rect 178556 124646 178598 124882
rect 178834 124646 181268 124882
rect 178556 124604 181268 124646
rect 180948 124244 181268 124604
rect 178556 124202 181268 124244
rect 178556 123966 178598 124202
rect 178834 123966 181268 124202
rect 178556 123924 181268 123966
rect 199164 122204 199484 130766
rect 249028 127602 249532 127644
rect 249028 127366 249070 127602
rect 249306 127366 249532 127602
rect 249028 127324 249532 127366
rect 248476 126922 248796 126964
rect 248476 126686 248518 126922
rect 248754 126686 248796 126922
rect 248476 124244 248796 126686
rect 245716 124202 248796 124244
rect 245716 123966 245758 124202
rect 245994 123966 248796 124202
rect 245716 123924 248796 123966
rect 249212 123564 249532 127324
rect 245348 123522 249532 123564
rect 245348 123286 245390 123522
rect 245626 123286 249532 123522
rect 245348 123244 249532 123286
rect 198612 121884 199484 122204
rect 198612 121524 198932 121884
rect 198428 121204 198932 121524
rect 198428 120844 198748 121204
rect 198244 120524 198748 120844
rect 198244 118124 198564 120524
rect 231732 119442 242356 119484
rect 231732 119206 231774 119442
rect 232010 119206 242078 119442
rect 242314 119206 242356 119442
rect 231732 119164 242356 119206
rect 142124 117804 145388 118124
rect 142124 116764 142444 117804
rect 145068 117444 145388 117804
rect 161628 118082 171332 118124
rect 161628 117846 163694 118082
rect 163930 117846 171332 118082
rect 161628 117804 171332 117846
rect 145068 117402 148884 117444
rect 145068 117166 148422 117402
rect 148658 117166 148884 117402
rect 145068 117124 148884 117166
rect 136788 116722 142444 116764
rect 136788 116486 136830 116722
rect 137066 116486 142444 116722
rect 136788 116444 142444 116486
rect 148564 116764 148884 117124
rect 161628 116764 161948 117804
rect 148564 116444 161948 116764
rect 171012 116764 171332 117804
rect 180948 117804 200404 118124
rect 180948 116764 181268 117804
rect 171012 116444 181268 116764
rect 190332 116444 190836 117804
rect 200084 116764 200404 117804
rect 219404 118082 229476 118124
rect 219404 117846 229198 118082
rect 229434 117846 229476 118082
rect 219404 117804 229476 117846
rect 219404 117444 219724 117804
rect 209836 117124 219724 117444
rect 209836 116764 210156 117124
rect 200084 116444 210156 116764
rect 238724 116722 245668 116764
rect 238724 116486 238766 116722
rect 239002 116486 245390 116722
rect 245626 116486 245668 116722
rect 238724 116444 245668 116486
rect 0 116026 444740 116068
rect 0 115790 5122 116026
rect 5358 115790 5442 116026
rect 5678 115790 5762 116026
rect 5998 115790 6082 116026
rect 6318 115790 6402 116026
rect 6638 115790 6722 116026
rect 6958 115790 7042 116026
rect 7278 115790 7362 116026
rect 7598 115790 7682 116026
rect 7918 115790 8002 116026
rect 8238 115790 8322 116026
rect 8558 115790 8642 116026
rect 8878 115790 89146 116026
rect 89382 115790 183146 116026
rect 183382 115790 277146 116026
rect 277382 115790 435862 116026
rect 436098 115790 436182 116026
rect 436418 115790 436502 116026
rect 436738 115790 436822 116026
rect 437058 115790 437142 116026
rect 437378 115790 437462 116026
rect 437698 115790 437782 116026
rect 438018 115790 438102 116026
rect 438338 115790 438422 116026
rect 438658 115790 438742 116026
rect 438978 115790 439062 116026
rect 439298 115790 439382 116026
rect 439618 115790 444740 116026
rect 0 115748 444740 115790
rect 157212 115362 163972 115404
rect 157212 115126 163694 115362
rect 163930 115126 163972 115362
rect 157212 115084 163972 115126
rect 157212 114724 157532 115084
rect 157212 114682 163972 114724
rect 157212 114446 163694 114682
rect 163930 114446 163972 114682
rect 157212 114404 163972 114446
rect 151508 114002 156612 114044
rect 151508 113766 152102 114002
rect 152338 113766 156612 114002
rect 151508 113724 156612 113766
rect 151508 113364 151828 113724
rect 146540 113322 151828 113364
rect 146540 113086 146582 113322
rect 146818 113086 151828 113322
rect 146540 113044 151828 113086
rect 156292 111324 156612 113724
rect 238908 114002 246036 114044
rect 238908 113766 245758 114002
rect 245994 113766 246036 114002
rect 238908 113724 246036 113766
rect 238908 112684 239228 113724
rect 164204 112642 239228 112684
rect 164204 112406 230670 112642
rect 230906 112406 239228 112642
rect 164204 112364 239228 112406
rect 164204 111324 164524 112364
rect 156292 111004 164524 111324
rect 84532 109922 87612 109964
rect 84532 109686 84574 109922
rect 84810 109686 87612 109922
rect 84532 109644 87612 109686
rect 87292 109284 87612 109644
rect 99436 109644 109508 109964
rect 99436 109284 99756 109644
rect 87292 108964 99756 109284
rect 109188 109284 109508 109644
rect 118756 109922 134900 109964
rect 118756 109686 134622 109922
rect 134858 109686 134900 109922
rect 118756 109644 134900 109686
rect 240012 109922 322948 109964
rect 240012 109686 240054 109922
rect 240290 109686 322670 109922
rect 322906 109686 322948 109922
rect 240012 109644 322948 109686
rect 118756 109284 119076 109644
rect 109188 108964 119076 109284
rect 99252 108284 99756 108964
rect 118572 108284 119076 108964
rect 178556 108562 183292 108604
rect 178556 108326 178598 108562
rect 178834 108326 183292 108562
rect 178556 108284 183292 108326
rect 182972 107244 183292 108284
rect 177820 107202 183292 107244
rect 177820 106966 177862 107202
rect 178098 106966 183292 107202
rect 177820 106924 183292 106966
rect 244796 106244 249716 106564
rect 244796 105884 245116 106244
rect 249396 105884 249716 106244
rect 156292 105842 163972 105884
rect 156292 105606 163694 105842
rect 163930 105606 163972 105842
rect 156292 105564 163972 105606
rect 244612 105564 245116 105884
rect 245532 105564 248796 105884
rect 249396 105564 250084 105884
rect 156292 105204 156612 105564
rect 156292 105162 163972 105204
rect 156292 104926 163694 105162
rect 163930 104926 163972 105162
rect 156292 104884 163972 104926
rect 244612 104524 244932 105564
rect 245532 105204 245852 105564
rect 245348 105162 245852 105204
rect 245348 104926 245390 105162
rect 245626 104926 245852 105162
rect 245348 104884 245852 104926
rect 248476 105204 248796 105564
rect 248476 104884 249164 105204
rect 137892 104482 165076 104524
rect 137892 104246 137934 104482
rect 138170 104246 164798 104482
rect 165034 104246 165076 104482
rect 137892 104204 165076 104246
rect 231732 104482 244932 104524
rect 231732 104246 231774 104482
rect 232010 104246 244932 104482
rect 231732 104204 244932 104246
rect 248844 104524 249164 104884
rect 248844 104204 249348 104524
rect 249028 103844 249348 104204
rect 178556 103802 188996 103844
rect 178556 103566 178598 103802
rect 178834 103566 188996 103802
rect 178556 103524 188996 103566
rect 245348 103802 249348 103844
rect 245348 103566 245390 103802
rect 245626 103566 249348 103802
rect 245348 103524 249348 103566
rect 249764 103844 250084 105564
rect 249764 103802 258916 103844
rect 249764 103566 258638 103802
rect 258874 103566 258916 103802
rect 249764 103524 258916 103566
rect 188676 103164 188996 103524
rect 176900 103122 180348 103164
rect 176900 102886 176942 103122
rect 177178 102886 180348 103122
rect 176900 102844 180348 102886
rect 188676 102844 193412 103164
rect 180028 101804 180348 102844
rect 193092 102484 193412 102844
rect 249028 102844 251188 103164
rect 193092 102442 229292 102484
rect 193092 102206 229014 102442
rect 229250 102206 229292 102442
rect 193092 102164 229292 102206
rect 249028 101804 249348 102844
rect 250868 102484 251188 102844
rect 253812 103122 261308 103164
rect 253812 102886 261030 103122
rect 261266 102886 261308 103122
rect 253812 102844 261308 102886
rect 253812 102484 254132 102844
rect 250868 102164 254132 102484
rect 272580 102442 323316 102484
rect 272580 102206 272622 102442
rect 272858 102206 323038 102442
rect 323274 102206 323316 102442
rect 272580 102164 323316 102206
rect 137340 101762 171516 101804
rect 137340 101526 137382 101762
rect 137618 101526 171238 101762
rect 171474 101526 171516 101762
rect 137340 101484 171516 101526
rect 180028 101762 249348 101804
rect 180028 101526 230670 101762
rect 230906 101526 249348 101762
rect 180028 101484 249348 101526
rect 270372 101762 324788 101804
rect 270372 101526 270414 101762
rect 270650 101526 324510 101762
rect 324746 101526 324788 101762
rect 270372 101484 324788 101526
rect 0 100708 444740 100750
rect 0 100472 122 100708
rect 358 100472 442 100708
rect 678 100472 762 100708
rect 998 100472 1082 100708
rect 1318 100472 1402 100708
rect 1638 100472 1722 100708
rect 1958 100472 2042 100708
rect 2278 100472 2362 100708
rect 2598 100472 2682 100708
rect 2918 100472 3002 100708
rect 3238 100472 3322 100708
rect 3558 100472 3642 100708
rect 3878 100472 104506 100708
rect 104742 100472 198506 100708
rect 198742 100472 292506 100708
rect 292742 100472 440862 100708
rect 441098 100472 441182 100708
rect 441418 100472 441502 100708
rect 441738 100472 441822 100708
rect 442058 100472 442142 100708
rect 442378 100472 442462 100708
rect 442698 100472 442782 100708
rect 443018 100472 443102 100708
rect 443338 100472 443422 100708
rect 443658 100472 443742 100708
rect 443978 100472 444062 100708
rect 444298 100472 444382 100708
rect 444618 100472 444740 100708
rect 0 100430 444740 100472
rect 145620 99722 161948 99764
rect 145620 99486 145662 99722
rect 145898 99486 161948 99722
rect 145620 99444 161948 99486
rect 161628 98404 161948 99444
rect 184444 99444 200588 99764
rect 178556 99042 181268 99084
rect 178556 98806 178598 99042
rect 178834 98806 181268 99042
rect 178556 98764 181268 98806
rect 161628 98362 165076 98404
rect 161628 98126 164798 98362
rect 165034 98126 165076 98362
rect 161628 98084 165076 98126
rect 180948 97724 181268 98764
rect 184444 97724 184764 99444
rect 200268 98404 200588 99444
rect 209652 99444 219908 99764
rect 242588 99722 258916 99764
rect 242588 99486 242630 99722
rect 242866 99486 258638 99722
rect 258874 99486 258916 99722
rect 242588 99444 258916 99486
rect 272580 99722 297188 99764
rect 272580 99486 272622 99722
rect 272858 99486 297188 99722
rect 272580 99444 297188 99486
rect 209652 98404 209972 99444
rect 200268 98084 209972 98404
rect 219588 98404 219908 99444
rect 296868 98404 297188 99444
rect 306252 99444 316508 99764
rect 306252 98404 306572 99444
rect 219588 98362 228924 98404
rect 219588 98126 228646 98362
rect 228882 98126 228924 98362
rect 219588 98084 228924 98126
rect 296868 98084 306572 98404
rect 316188 98404 316508 99444
rect 316188 98362 322948 98404
rect 316188 98126 322670 98362
rect 322906 98126 322948 98362
rect 316188 98084 322948 98126
rect 180948 97404 184764 97724
rect 177820 96322 183108 96364
rect 177820 96086 177862 96322
rect 178098 96086 183108 96322
rect 177820 96044 183108 96086
rect 245348 96322 249716 96364
rect 245348 96086 245390 96322
rect 245626 96086 249716 96322
rect 245348 96044 249716 96086
rect 155188 94282 163972 94324
rect 155188 94046 163694 94282
rect 163930 94046 163972 94282
rect 155188 94004 163972 94046
rect 74412 93602 84852 93644
rect 74412 93366 74454 93602
rect 74690 93366 84574 93602
rect 84810 93366 84852 93602
rect 74412 93324 84852 93366
rect 155188 90882 155508 94004
rect 182788 92964 183108 96044
rect 182788 92644 183660 92964
rect 155188 90646 155230 90882
rect 155466 90646 155508 90882
rect 155188 90604 155508 90646
rect 183340 88884 183660 92644
rect 249396 90202 249716 96044
rect 249396 89966 249438 90202
rect 249674 89966 249716 90202
rect 249396 89924 249716 89966
rect 178556 88842 183660 88884
rect 178556 88606 178598 88842
rect 178834 88606 183660 88842
rect 178556 88564 183660 88606
rect 249396 88842 264068 88884
rect 249396 88606 249438 88842
rect 249674 88606 263790 88842
rect 264026 88606 264068 88842
rect 249396 88564 264068 88606
rect 251604 88162 261860 88204
rect 251604 87926 251646 88162
rect 251882 87926 259558 88162
rect 259794 87926 261582 88162
rect 261818 87926 261860 88162
rect 251604 87884 261860 87926
rect 0 85390 444740 85432
rect 0 85154 5122 85390
rect 5358 85154 5442 85390
rect 5678 85154 5762 85390
rect 5998 85154 6082 85390
rect 6318 85154 6402 85390
rect 6638 85154 6722 85390
rect 6958 85154 7042 85390
rect 7278 85154 7362 85390
rect 7598 85154 7682 85390
rect 7918 85154 8002 85390
rect 8238 85154 8322 85390
rect 8558 85154 8642 85390
rect 8878 85154 435862 85390
rect 436098 85154 436182 85390
rect 436418 85154 436502 85390
rect 436738 85154 436822 85390
rect 437058 85154 437142 85390
rect 437378 85154 437462 85390
rect 437698 85154 437782 85390
rect 438018 85154 438102 85390
rect 438338 85154 438422 85390
rect 438658 85154 438742 85390
rect 438978 85154 439062 85390
rect 439298 85154 439382 85390
rect 439618 85154 444740 85390
rect 0 85112 444740 85154
rect 148380 73882 148700 73924
rect 148380 73646 148422 73882
rect 148658 73646 148700 73882
rect 148380 73244 148700 73646
rect 155924 73882 170228 73924
rect 155924 73646 155966 73882
rect 156202 73646 169950 73882
rect 170186 73646 170228 73882
rect 155924 73604 170228 73646
rect 249764 73882 264436 73924
rect 249764 73646 249806 73882
rect 250042 73646 264158 73882
rect 264394 73646 264436 73882
rect 249764 73604 264436 73646
rect 144516 73202 148700 73244
rect 144516 72966 144558 73202
rect 144794 72966 148700 73202
rect 144516 72924 148700 72966
rect 0 70072 444740 70114
rect 0 69836 122 70072
rect 358 69836 442 70072
rect 678 69836 762 70072
rect 998 69836 1082 70072
rect 1318 69836 1402 70072
rect 1638 69836 1722 70072
rect 1958 69836 2042 70072
rect 2278 69836 2362 70072
rect 2598 69836 2682 70072
rect 2918 69836 3002 70072
rect 3238 69836 3322 70072
rect 3558 69836 3642 70072
rect 3878 69836 440862 70072
rect 441098 69836 441182 70072
rect 441418 69836 441502 70072
rect 441738 69836 441822 70072
rect 442058 69836 442142 70072
rect 442378 69836 442462 70072
rect 442698 69836 442782 70072
rect 443018 69836 443102 70072
rect 443338 69836 443422 70072
rect 443658 69836 443742 70072
rect 443978 69836 444062 70072
rect 444298 69836 444382 70072
rect 444618 69836 444740 70072
rect 0 69794 444740 69836
rect 144516 64362 148148 64404
rect 144516 64126 144558 64362
rect 144794 64126 148148 64362
rect 144516 64084 148148 64126
rect 147828 63724 148148 64084
rect 144700 63682 148148 63724
rect 144700 63446 144742 63682
rect 144978 63446 148148 63682
rect 144700 63404 148148 63446
rect 238540 60282 242908 60324
rect 238540 60046 238582 60282
rect 238818 60046 242908 60282
rect 238540 60004 242908 60046
rect 242588 59644 242908 60004
rect 237252 59602 242908 59644
rect 237252 59366 237294 59602
rect 237530 59366 242908 59602
rect 237252 59324 242908 59366
rect 0 54754 444740 54796
rect 0 54518 5122 54754
rect 5358 54518 5442 54754
rect 5678 54518 5762 54754
rect 5998 54518 6082 54754
rect 6318 54518 6402 54754
rect 6638 54518 6722 54754
rect 6958 54518 7042 54754
rect 7278 54518 7362 54754
rect 7598 54518 7682 54754
rect 7918 54518 8002 54754
rect 8238 54518 8322 54754
rect 8558 54518 8642 54754
rect 8878 54518 435862 54754
rect 436098 54518 436182 54754
rect 436418 54518 436502 54754
rect 436738 54518 436822 54754
rect 437058 54518 437142 54754
rect 437378 54518 437462 54754
rect 437698 54518 437782 54754
rect 438018 54518 438102 54754
rect 438338 54518 438422 54754
rect 438658 54518 438742 54754
rect 438978 54518 439062 54754
rect 439298 54518 439382 54754
rect 439618 54518 444740 54754
rect 0 54476 444740 54518
rect 269084 52122 270876 52164
rect 269084 51886 270598 52122
rect 270834 51886 270876 52122
rect 269084 51844 270876 51886
rect 102380 51442 142628 51484
rect 102380 51206 102422 51442
rect 102658 51206 142350 51442
rect 142586 51206 142628 51442
rect 102380 51164 142628 51206
rect 238540 51442 248796 51484
rect 238540 51206 238582 51442
rect 238818 51206 248796 51442
rect 238540 51164 248796 51206
rect 93548 50762 187340 50804
rect 93548 50526 93590 50762
rect 93826 50526 187062 50762
rect 187298 50526 187340 50762
rect 93548 50484 187340 50526
rect 237620 50762 242908 50804
rect 237620 50526 237662 50762
rect 237898 50526 242908 50762
rect 237620 50484 242908 50526
rect 74412 49402 88532 49444
rect 74412 49166 74454 49402
rect 74690 49166 88254 49402
rect 88490 49166 88532 49402
rect 74412 49124 88532 49166
rect 105140 49402 145756 49444
rect 105140 49166 105182 49402
rect 105418 49166 145478 49402
rect 145714 49166 145756 49402
rect 105140 49124 145756 49166
rect 147828 49402 148148 50484
rect 147828 49166 147870 49402
rect 148106 49166 148148 49402
rect 147828 49124 148148 49166
rect 167884 49402 182188 49444
rect 167884 49166 167926 49402
rect 168162 49166 181910 49402
rect 182146 49166 182188 49402
rect 167884 49124 182188 49166
rect 67788 48722 88348 48764
rect 67788 48486 67830 48722
rect 68066 48486 73166 48722
rect 73402 48486 88070 48722
rect 88306 48486 88348 48722
rect 67788 48444 88348 48486
rect 154636 48722 191572 48764
rect 154636 48486 154678 48722
rect 154914 48486 167558 48722
rect 167794 48486 191294 48722
rect 191530 48486 191572 48722
rect 154636 48444 191572 48486
rect 242588 48084 242908 50484
rect 248476 50124 248796 51164
rect 251236 51164 260020 51484
rect 251236 50124 251556 51164
rect 248476 49804 251556 50124
rect 259700 50124 260020 51164
rect 269084 50124 269404 51844
rect 259700 49804 269404 50124
rect 248844 48722 264436 48764
rect 248844 48486 248886 48722
rect 249122 48486 264158 48722
rect 264394 48486 264436 48722
rect 248844 48444 264436 48486
rect 159972 48042 182004 48084
rect 159972 47806 160014 48042
rect 160250 47806 169030 48042
rect 169266 47806 181726 48042
rect 181962 47806 182004 48042
rect 159972 47764 182004 47806
rect 242588 48042 250636 48084
rect 242588 47806 250358 48042
rect 250594 47806 250636 48042
rect 242588 47764 250636 47806
rect 260988 48042 276212 48084
rect 260988 47806 261030 48042
rect 261266 47806 275934 48042
rect 276170 47806 276212 48042
rect 260988 47764 276212 47806
rect 110292 47362 159188 47404
rect 110292 47126 110334 47362
rect 110570 47126 158910 47362
rect 159146 47126 159188 47362
rect 110292 47084 159188 47126
rect 248476 47362 264068 47404
rect 248476 47126 248518 47362
rect 248754 47126 263790 47362
rect 264026 47126 264068 47362
rect 248476 47084 264068 47126
rect 107348 46682 157716 46724
rect 107348 46446 107390 46682
rect 107626 46446 157438 46682
rect 157674 46446 157716 46682
rect 107348 46404 157716 46446
rect 162732 46682 182004 46724
rect 162732 46446 162774 46682
rect 163010 46446 181726 46682
rect 181962 46446 182004 46682
rect 162732 46404 182004 46446
rect 204132 46682 253028 46724
rect 204132 46446 204174 46682
rect 204410 46446 252750 46682
rect 252986 46446 253028 46682
rect 204132 46404 253028 46446
rect 261724 46682 276028 46724
rect 261724 46446 261766 46682
rect 262002 46446 275750 46682
rect 275986 46446 276028 46682
rect 261724 46404 276028 46446
rect 0 39436 444740 39478
rect 0 39200 122 39436
rect 358 39200 442 39436
rect 678 39200 762 39436
rect 998 39200 1082 39436
rect 1318 39200 1402 39436
rect 1638 39200 1722 39436
rect 1958 39200 2042 39436
rect 2278 39200 2362 39436
rect 2598 39200 2682 39436
rect 2918 39200 3002 39436
rect 3238 39200 3322 39436
rect 3558 39200 3642 39436
rect 3878 39200 440862 39436
rect 441098 39200 441182 39436
rect 441418 39200 441502 39436
rect 441738 39200 441822 39436
rect 442058 39200 442142 39436
rect 442378 39200 442462 39436
rect 442698 39200 442782 39436
rect 443018 39200 443102 39436
rect 443338 39200 443422 39436
rect 443658 39200 443742 39436
rect 443978 39200 444062 39436
rect 444298 39200 444382 39436
rect 444618 39200 444740 39436
rect 0 39158 444740 39200
rect 0 24118 444740 24160
rect 0 23882 5122 24118
rect 5358 23882 5442 24118
rect 5678 23882 5762 24118
rect 5998 23882 6082 24118
rect 6318 23882 6402 24118
rect 6638 23882 6722 24118
rect 6958 23882 7042 24118
rect 7278 23882 7362 24118
rect 7598 23882 7682 24118
rect 7918 23882 8002 24118
rect 8238 23882 8322 24118
rect 8558 23882 8642 24118
rect 8878 23882 435862 24118
rect 436098 23882 436182 24118
rect 436418 23882 436502 24118
rect 436738 23882 436822 24118
rect 437058 23882 437142 24118
rect 437378 23882 437462 24118
rect 437698 23882 437782 24118
rect 438018 23882 438102 24118
rect 438338 23882 438422 24118
rect 438658 23882 438742 24118
rect 438978 23882 439062 24118
rect 439298 23882 439382 24118
rect 439618 23882 444740 24118
rect 0 23840 444740 23882
rect 5000 8878 439740 9000
rect 5000 8642 5122 8878
rect 5358 8642 5442 8878
rect 5678 8642 5762 8878
rect 5998 8642 6082 8878
rect 6318 8642 6402 8878
rect 6638 8642 6722 8878
rect 6958 8642 7042 8878
rect 7278 8642 7362 8878
rect 7598 8642 7682 8878
rect 7918 8642 8002 8878
rect 8238 8642 8322 8878
rect 8558 8642 8642 8878
rect 8878 8642 435862 8878
rect 436098 8642 436182 8878
rect 436418 8642 436502 8878
rect 436738 8642 436822 8878
rect 437058 8642 437142 8878
rect 437378 8642 437462 8878
rect 437698 8642 437782 8878
rect 438018 8642 438102 8878
rect 438338 8642 438422 8878
rect 438658 8642 438742 8878
rect 438978 8642 439062 8878
rect 439298 8642 439382 8878
rect 439618 8642 439740 8878
rect 5000 8558 439740 8642
rect 5000 8322 5122 8558
rect 5358 8322 5442 8558
rect 5678 8322 5762 8558
rect 5998 8322 6082 8558
rect 6318 8322 6402 8558
rect 6638 8322 6722 8558
rect 6958 8322 7042 8558
rect 7278 8322 7362 8558
rect 7598 8322 7682 8558
rect 7918 8322 8002 8558
rect 8238 8322 8322 8558
rect 8558 8322 8642 8558
rect 8878 8322 435862 8558
rect 436098 8322 436182 8558
rect 436418 8322 436502 8558
rect 436738 8322 436822 8558
rect 437058 8322 437142 8558
rect 437378 8322 437462 8558
rect 437698 8322 437782 8558
rect 438018 8322 438102 8558
rect 438338 8322 438422 8558
rect 438658 8322 438742 8558
rect 438978 8322 439062 8558
rect 439298 8322 439382 8558
rect 439618 8322 439740 8558
rect 5000 8238 439740 8322
rect 5000 8002 5122 8238
rect 5358 8002 5442 8238
rect 5678 8002 5762 8238
rect 5998 8002 6082 8238
rect 6318 8002 6402 8238
rect 6638 8002 6722 8238
rect 6958 8002 7042 8238
rect 7278 8002 7362 8238
rect 7598 8002 7682 8238
rect 7918 8002 8002 8238
rect 8238 8002 8322 8238
rect 8558 8002 8642 8238
rect 8878 8002 435862 8238
rect 436098 8002 436182 8238
rect 436418 8002 436502 8238
rect 436738 8002 436822 8238
rect 437058 8002 437142 8238
rect 437378 8002 437462 8238
rect 437698 8002 437782 8238
rect 438018 8002 438102 8238
rect 438338 8002 438422 8238
rect 438658 8002 438742 8238
rect 438978 8002 439062 8238
rect 439298 8002 439382 8238
rect 439618 8002 439740 8238
rect 5000 7918 439740 8002
rect 5000 7682 5122 7918
rect 5358 7682 5442 7918
rect 5678 7682 5762 7918
rect 5998 7682 6082 7918
rect 6318 7682 6402 7918
rect 6638 7682 6722 7918
rect 6958 7682 7042 7918
rect 7278 7682 7362 7918
rect 7598 7682 7682 7918
rect 7918 7682 8002 7918
rect 8238 7682 8322 7918
rect 8558 7682 8642 7918
rect 8878 7682 435862 7918
rect 436098 7682 436182 7918
rect 436418 7682 436502 7918
rect 436738 7682 436822 7918
rect 437058 7682 437142 7918
rect 437378 7682 437462 7918
rect 437698 7682 437782 7918
rect 438018 7682 438102 7918
rect 438338 7682 438422 7918
rect 438658 7682 438742 7918
rect 438978 7682 439062 7918
rect 439298 7682 439382 7918
rect 439618 7682 439740 7918
rect 5000 7598 439740 7682
rect 5000 7362 5122 7598
rect 5358 7362 5442 7598
rect 5678 7362 5762 7598
rect 5998 7362 6082 7598
rect 6318 7362 6402 7598
rect 6638 7362 6722 7598
rect 6958 7362 7042 7598
rect 7278 7362 7362 7598
rect 7598 7362 7682 7598
rect 7918 7362 8002 7598
rect 8238 7362 8322 7598
rect 8558 7362 8642 7598
rect 8878 7362 435862 7598
rect 436098 7362 436182 7598
rect 436418 7362 436502 7598
rect 436738 7362 436822 7598
rect 437058 7362 437142 7598
rect 437378 7362 437462 7598
rect 437698 7362 437782 7598
rect 438018 7362 438102 7598
rect 438338 7362 438422 7598
rect 438658 7362 438742 7598
rect 438978 7362 439062 7598
rect 439298 7362 439382 7598
rect 439618 7362 439740 7598
rect 5000 7278 439740 7362
rect 5000 7042 5122 7278
rect 5358 7042 5442 7278
rect 5678 7042 5762 7278
rect 5998 7042 6082 7278
rect 6318 7042 6402 7278
rect 6638 7042 6722 7278
rect 6958 7042 7042 7278
rect 7278 7042 7362 7278
rect 7598 7042 7682 7278
rect 7918 7042 8002 7278
rect 8238 7042 8322 7278
rect 8558 7042 8642 7278
rect 8878 7042 435862 7278
rect 436098 7042 436182 7278
rect 436418 7042 436502 7278
rect 436738 7042 436822 7278
rect 437058 7042 437142 7278
rect 437378 7042 437462 7278
rect 437698 7042 437782 7278
rect 438018 7042 438102 7278
rect 438338 7042 438422 7278
rect 438658 7042 438742 7278
rect 438978 7042 439062 7278
rect 439298 7042 439382 7278
rect 439618 7042 439740 7278
rect 5000 6958 439740 7042
rect 5000 6722 5122 6958
rect 5358 6722 5442 6958
rect 5678 6722 5762 6958
rect 5998 6722 6082 6958
rect 6318 6722 6402 6958
rect 6638 6722 6722 6958
rect 6958 6722 7042 6958
rect 7278 6722 7362 6958
rect 7598 6722 7682 6958
rect 7918 6722 8002 6958
rect 8238 6722 8322 6958
rect 8558 6722 8642 6958
rect 8878 6722 435862 6958
rect 436098 6722 436182 6958
rect 436418 6722 436502 6958
rect 436738 6722 436822 6958
rect 437058 6722 437142 6958
rect 437378 6722 437462 6958
rect 437698 6722 437782 6958
rect 438018 6722 438102 6958
rect 438338 6722 438422 6958
rect 438658 6722 438742 6958
rect 438978 6722 439062 6958
rect 439298 6722 439382 6958
rect 439618 6722 439740 6958
rect 5000 6638 439740 6722
rect 5000 6402 5122 6638
rect 5358 6402 5442 6638
rect 5678 6402 5762 6638
rect 5998 6402 6082 6638
rect 6318 6402 6402 6638
rect 6638 6402 6722 6638
rect 6958 6402 7042 6638
rect 7278 6402 7362 6638
rect 7598 6402 7682 6638
rect 7918 6402 8002 6638
rect 8238 6402 8322 6638
rect 8558 6402 8642 6638
rect 8878 6402 435862 6638
rect 436098 6402 436182 6638
rect 436418 6402 436502 6638
rect 436738 6402 436822 6638
rect 437058 6402 437142 6638
rect 437378 6402 437462 6638
rect 437698 6402 437782 6638
rect 438018 6402 438102 6638
rect 438338 6402 438422 6638
rect 438658 6402 438742 6638
rect 438978 6402 439062 6638
rect 439298 6402 439382 6638
rect 439618 6402 439740 6638
rect 5000 6318 439740 6402
rect 5000 6082 5122 6318
rect 5358 6082 5442 6318
rect 5678 6082 5762 6318
rect 5998 6082 6082 6318
rect 6318 6082 6402 6318
rect 6638 6082 6722 6318
rect 6958 6082 7042 6318
rect 7278 6082 7362 6318
rect 7598 6082 7682 6318
rect 7918 6082 8002 6318
rect 8238 6082 8322 6318
rect 8558 6082 8642 6318
rect 8878 6082 435862 6318
rect 436098 6082 436182 6318
rect 436418 6082 436502 6318
rect 436738 6082 436822 6318
rect 437058 6082 437142 6318
rect 437378 6082 437462 6318
rect 437698 6082 437782 6318
rect 438018 6082 438102 6318
rect 438338 6082 438422 6318
rect 438658 6082 438742 6318
rect 438978 6082 439062 6318
rect 439298 6082 439382 6318
rect 439618 6082 439740 6318
rect 5000 5998 439740 6082
rect 5000 5762 5122 5998
rect 5358 5762 5442 5998
rect 5678 5762 5762 5998
rect 5998 5762 6082 5998
rect 6318 5762 6402 5998
rect 6638 5762 6722 5998
rect 6958 5762 7042 5998
rect 7278 5762 7362 5998
rect 7598 5762 7682 5998
rect 7918 5762 8002 5998
rect 8238 5762 8322 5998
rect 8558 5762 8642 5998
rect 8878 5762 435862 5998
rect 436098 5762 436182 5998
rect 436418 5762 436502 5998
rect 436738 5762 436822 5998
rect 437058 5762 437142 5998
rect 437378 5762 437462 5998
rect 437698 5762 437782 5998
rect 438018 5762 438102 5998
rect 438338 5762 438422 5998
rect 438658 5762 438742 5998
rect 438978 5762 439062 5998
rect 439298 5762 439382 5998
rect 439618 5762 439740 5998
rect 5000 5678 439740 5762
rect 5000 5442 5122 5678
rect 5358 5442 5442 5678
rect 5678 5442 5762 5678
rect 5998 5442 6082 5678
rect 6318 5442 6402 5678
rect 6638 5442 6722 5678
rect 6958 5442 7042 5678
rect 7278 5442 7362 5678
rect 7598 5442 7682 5678
rect 7918 5442 8002 5678
rect 8238 5442 8322 5678
rect 8558 5442 8642 5678
rect 8878 5442 435862 5678
rect 436098 5442 436182 5678
rect 436418 5442 436502 5678
rect 436738 5442 436822 5678
rect 437058 5442 437142 5678
rect 437378 5442 437462 5678
rect 437698 5442 437782 5678
rect 438018 5442 438102 5678
rect 438338 5442 438422 5678
rect 438658 5442 438742 5678
rect 438978 5442 439062 5678
rect 439298 5442 439382 5678
rect 439618 5442 439740 5678
rect 5000 5358 439740 5442
rect 5000 5122 5122 5358
rect 5358 5122 5442 5358
rect 5678 5122 5762 5358
rect 5998 5122 6082 5358
rect 6318 5122 6402 5358
rect 6638 5122 6722 5358
rect 6958 5122 7042 5358
rect 7278 5122 7362 5358
rect 7598 5122 7682 5358
rect 7918 5122 8002 5358
rect 8238 5122 8322 5358
rect 8558 5122 8642 5358
rect 8878 5122 435862 5358
rect 436098 5122 436182 5358
rect 436418 5122 436502 5358
rect 436738 5122 436822 5358
rect 437058 5122 437142 5358
rect 437378 5122 437462 5358
rect 437698 5122 437782 5358
rect 438018 5122 438102 5358
rect 438338 5122 438422 5358
rect 438658 5122 438742 5358
rect 438978 5122 439062 5358
rect 439298 5122 439382 5358
rect 439618 5122 439740 5358
rect 5000 5000 439740 5122
rect 0 3878 444740 4000
rect 0 3642 122 3878
rect 358 3642 442 3878
rect 678 3642 762 3878
rect 998 3642 1082 3878
rect 1318 3642 1402 3878
rect 1638 3642 1722 3878
rect 1958 3642 2042 3878
rect 2278 3642 2362 3878
rect 2598 3642 2682 3878
rect 2918 3642 3002 3878
rect 3238 3642 3322 3878
rect 3558 3642 3642 3878
rect 3878 3642 440862 3878
rect 441098 3642 441182 3878
rect 441418 3642 441502 3878
rect 441738 3642 441822 3878
rect 442058 3642 442142 3878
rect 442378 3642 442462 3878
rect 442698 3642 442782 3878
rect 443018 3642 443102 3878
rect 443338 3642 443422 3878
rect 443658 3642 443742 3878
rect 443978 3642 444062 3878
rect 444298 3642 444382 3878
rect 444618 3642 444740 3878
rect 0 3558 444740 3642
rect 0 3322 122 3558
rect 358 3322 442 3558
rect 678 3322 762 3558
rect 998 3322 1082 3558
rect 1318 3322 1402 3558
rect 1638 3322 1722 3558
rect 1958 3322 2042 3558
rect 2278 3322 2362 3558
rect 2598 3322 2682 3558
rect 2918 3322 3002 3558
rect 3238 3322 3322 3558
rect 3558 3322 3642 3558
rect 3878 3322 440862 3558
rect 441098 3322 441182 3558
rect 441418 3322 441502 3558
rect 441738 3322 441822 3558
rect 442058 3322 442142 3558
rect 442378 3322 442462 3558
rect 442698 3322 442782 3558
rect 443018 3322 443102 3558
rect 443338 3322 443422 3558
rect 443658 3322 443742 3558
rect 443978 3322 444062 3558
rect 444298 3322 444382 3558
rect 444618 3322 444740 3558
rect 0 3238 444740 3322
rect 0 3002 122 3238
rect 358 3002 442 3238
rect 678 3002 762 3238
rect 998 3002 1082 3238
rect 1318 3002 1402 3238
rect 1638 3002 1722 3238
rect 1958 3002 2042 3238
rect 2278 3002 2362 3238
rect 2598 3002 2682 3238
rect 2918 3002 3002 3238
rect 3238 3002 3322 3238
rect 3558 3002 3642 3238
rect 3878 3002 440862 3238
rect 441098 3002 441182 3238
rect 441418 3002 441502 3238
rect 441738 3002 441822 3238
rect 442058 3002 442142 3238
rect 442378 3002 442462 3238
rect 442698 3002 442782 3238
rect 443018 3002 443102 3238
rect 443338 3002 443422 3238
rect 443658 3002 443742 3238
rect 443978 3002 444062 3238
rect 444298 3002 444382 3238
rect 444618 3002 444740 3238
rect 0 2918 444740 3002
rect 0 2682 122 2918
rect 358 2682 442 2918
rect 678 2682 762 2918
rect 998 2682 1082 2918
rect 1318 2682 1402 2918
rect 1638 2682 1722 2918
rect 1958 2682 2042 2918
rect 2278 2682 2362 2918
rect 2598 2682 2682 2918
rect 2918 2682 3002 2918
rect 3238 2682 3322 2918
rect 3558 2682 3642 2918
rect 3878 2682 440862 2918
rect 441098 2682 441182 2918
rect 441418 2682 441502 2918
rect 441738 2682 441822 2918
rect 442058 2682 442142 2918
rect 442378 2682 442462 2918
rect 442698 2682 442782 2918
rect 443018 2682 443102 2918
rect 443338 2682 443422 2918
rect 443658 2682 443742 2918
rect 443978 2682 444062 2918
rect 444298 2682 444382 2918
rect 444618 2682 444740 2918
rect 0 2598 444740 2682
rect 0 2362 122 2598
rect 358 2362 442 2598
rect 678 2362 762 2598
rect 998 2362 1082 2598
rect 1318 2362 1402 2598
rect 1638 2362 1722 2598
rect 1958 2362 2042 2598
rect 2278 2362 2362 2598
rect 2598 2362 2682 2598
rect 2918 2362 3002 2598
rect 3238 2362 3322 2598
rect 3558 2362 3642 2598
rect 3878 2362 440862 2598
rect 441098 2362 441182 2598
rect 441418 2362 441502 2598
rect 441738 2362 441822 2598
rect 442058 2362 442142 2598
rect 442378 2362 442462 2598
rect 442698 2362 442782 2598
rect 443018 2362 443102 2598
rect 443338 2362 443422 2598
rect 443658 2362 443742 2598
rect 443978 2362 444062 2598
rect 444298 2362 444382 2598
rect 444618 2362 444740 2598
rect 0 2278 444740 2362
rect 0 2042 122 2278
rect 358 2042 442 2278
rect 678 2042 762 2278
rect 998 2042 1082 2278
rect 1318 2042 1402 2278
rect 1638 2042 1722 2278
rect 1958 2042 2042 2278
rect 2278 2042 2362 2278
rect 2598 2042 2682 2278
rect 2918 2042 3002 2278
rect 3238 2042 3322 2278
rect 3558 2042 3642 2278
rect 3878 2042 440862 2278
rect 441098 2042 441182 2278
rect 441418 2042 441502 2278
rect 441738 2042 441822 2278
rect 442058 2042 442142 2278
rect 442378 2042 442462 2278
rect 442698 2042 442782 2278
rect 443018 2042 443102 2278
rect 443338 2042 443422 2278
rect 443658 2042 443742 2278
rect 443978 2042 444062 2278
rect 444298 2042 444382 2278
rect 444618 2042 444740 2278
rect 0 1958 444740 2042
rect 0 1722 122 1958
rect 358 1722 442 1958
rect 678 1722 762 1958
rect 998 1722 1082 1958
rect 1318 1722 1402 1958
rect 1638 1722 1722 1958
rect 1958 1722 2042 1958
rect 2278 1722 2362 1958
rect 2598 1722 2682 1958
rect 2918 1722 3002 1958
rect 3238 1722 3322 1958
rect 3558 1722 3642 1958
rect 3878 1722 440862 1958
rect 441098 1722 441182 1958
rect 441418 1722 441502 1958
rect 441738 1722 441822 1958
rect 442058 1722 442142 1958
rect 442378 1722 442462 1958
rect 442698 1722 442782 1958
rect 443018 1722 443102 1958
rect 443338 1722 443422 1958
rect 443658 1722 443742 1958
rect 443978 1722 444062 1958
rect 444298 1722 444382 1958
rect 444618 1722 444740 1958
rect 0 1638 444740 1722
rect 0 1402 122 1638
rect 358 1402 442 1638
rect 678 1402 762 1638
rect 998 1402 1082 1638
rect 1318 1402 1402 1638
rect 1638 1402 1722 1638
rect 1958 1402 2042 1638
rect 2278 1402 2362 1638
rect 2598 1402 2682 1638
rect 2918 1402 3002 1638
rect 3238 1402 3322 1638
rect 3558 1402 3642 1638
rect 3878 1402 440862 1638
rect 441098 1402 441182 1638
rect 441418 1402 441502 1638
rect 441738 1402 441822 1638
rect 442058 1402 442142 1638
rect 442378 1402 442462 1638
rect 442698 1402 442782 1638
rect 443018 1402 443102 1638
rect 443338 1402 443422 1638
rect 443658 1402 443742 1638
rect 443978 1402 444062 1638
rect 444298 1402 444382 1638
rect 444618 1402 444740 1638
rect 0 1318 444740 1402
rect 0 1082 122 1318
rect 358 1082 442 1318
rect 678 1082 762 1318
rect 998 1082 1082 1318
rect 1318 1082 1402 1318
rect 1638 1082 1722 1318
rect 1958 1082 2042 1318
rect 2278 1082 2362 1318
rect 2598 1082 2682 1318
rect 2918 1082 3002 1318
rect 3238 1082 3322 1318
rect 3558 1082 3642 1318
rect 3878 1082 440862 1318
rect 441098 1082 441182 1318
rect 441418 1082 441502 1318
rect 441738 1082 441822 1318
rect 442058 1082 442142 1318
rect 442378 1082 442462 1318
rect 442698 1082 442782 1318
rect 443018 1082 443102 1318
rect 443338 1082 443422 1318
rect 443658 1082 443742 1318
rect 443978 1082 444062 1318
rect 444298 1082 444382 1318
rect 444618 1082 444740 1318
rect 0 998 444740 1082
rect 0 762 122 998
rect 358 762 442 998
rect 678 762 762 998
rect 998 762 1082 998
rect 1318 762 1402 998
rect 1638 762 1722 998
rect 1958 762 2042 998
rect 2278 762 2362 998
rect 2598 762 2682 998
rect 2918 762 3002 998
rect 3238 762 3322 998
rect 3558 762 3642 998
rect 3878 762 440862 998
rect 441098 762 441182 998
rect 441418 762 441502 998
rect 441738 762 441822 998
rect 442058 762 442142 998
rect 442378 762 442462 998
rect 442698 762 442782 998
rect 443018 762 443102 998
rect 443338 762 443422 998
rect 443658 762 443742 998
rect 443978 762 444062 998
rect 444298 762 444382 998
rect 444618 762 444740 998
rect 0 678 444740 762
rect 0 442 122 678
rect 358 442 442 678
rect 678 442 762 678
rect 998 442 1082 678
rect 1318 442 1402 678
rect 1638 442 1722 678
rect 1958 442 2042 678
rect 2278 442 2362 678
rect 2598 442 2682 678
rect 2918 442 3002 678
rect 3238 442 3322 678
rect 3558 442 3642 678
rect 3878 442 440862 678
rect 441098 442 441182 678
rect 441418 442 441502 678
rect 441738 442 441822 678
rect 442058 442 442142 678
rect 442378 442 442462 678
rect 442698 442 442782 678
rect 443018 442 443102 678
rect 443338 442 443422 678
rect 443658 442 443742 678
rect 443978 442 444062 678
rect 444298 442 444382 678
rect 444618 442 444740 678
rect 0 358 444740 442
rect 0 122 122 358
rect 358 122 442 358
rect 678 122 762 358
rect 998 122 1082 358
rect 1318 122 1402 358
rect 1638 122 1722 358
rect 1958 122 2042 358
rect 2278 122 2362 358
rect 2598 122 2682 358
rect 2918 122 3002 358
rect 3238 122 3322 358
rect 3558 122 3642 358
rect 3878 122 440862 358
rect 441098 122 441182 358
rect 441418 122 441502 358
rect 441738 122 441822 358
rect 442058 122 442142 358
rect 442378 122 442462 358
rect 442698 122 442782 358
rect 443018 122 443102 358
rect 443338 122 443422 358
rect 443658 122 443742 358
rect 443978 122 444062 358
rect 444298 122 444382 358
rect 444618 122 444740 358
rect 0 0 444740 122
use sb_0__0_  sb_0__0_
timestamp 1603810449
transform 1 0 48895 0 1 47824
box 1 0 27528 28000
use grid_io_bottom  grid_io_bottom_1__0_
timestamp 1603810449
transform 1 0 89896 0 1 18824
box 0 0 38862 16000
use cbx_1__0_  cbx_1__0_
timestamp 1603810449
transform 1 0 89896 0 1 53824
box 0 0 40000 16000
use sb_1__0_  sb_1__0_
timestamp 1603810449
transform 1 0 142896 0 1 47824
box 0 0 28000 28000
use grid_io_bottom  grid_io_bottom_2__0_
timestamp 1603810449
transform 1 0 183896 0 1 18824
box 0 0 38862 16000
use cbx_1__0_  cbx_2__0_
timestamp 1603810449
transform 1 0 183896 0 1 53824
box 0 0 40000 16000
use sb_1__0_  sb_2__0_
timestamp 1603810449
transform 1 0 236896 0 1 47824
box 0 0 28000 28000
use grid_io_bottom  grid_io_bottom_3__0_
timestamp 1603810449
transform 1 0 277896 0 1 18824
box 0 0 38862 16000
use cbx_1__0_  cbx_3__0_
timestamp 1603810449
transform 1 0 277896 0 1 53824
box 0 0 40000 16000
use sb_3__0_  sb_3__0_
timestamp 1603810449
transform 1 0 330896 0 1 47824
box 0 0 27403 28000
use grid_io_left  grid_io_left_0__1_
timestamp 1603810449
transform 1 0 19896 0 1 88824
box 0 0 16000 38752
use cby_0__1_  cby_0__1_
timestamp 1603810449
transform 1 0 54896 0 1 88824
box 0 0 16000 40000
use grid_clb  grid_clb_1__1_
timestamp 1603810449
transform 1 0 84896 0 1 83824
box 0 0 50000 50000
use cby_1__1_  cby_1__1_
timestamp 1603810449
transform 1 0 148896 0 1 88824
box 0 0 16000 40000
use grid_clb  grid_clb_2__1_
timestamp 1603810449
transform 1 0 178896 0 1 83824
box 0 0 50000 50000
use cby_1__1_  cby_2__1_
timestamp 1603810449
transform 1 0 242896 0 1 88824
box 0 0 16000 40000
use grid_clb  grid_clb_3__1_
timestamp 1603810449
transform 1 0 272896 0 1 83824
box 0 0 50000 50000
use cby_3__1_  cby_3__1_
timestamp 1603810449
transform 1 0 336896 0 1 88824
box 0 0 16000 40000
use grid_io_right  grid_io_right_4__1_
timestamp 1603810449
transform 1 0 408896 0 1 88824
box 0 0 16000 38752
use grid_io_left  grid_io_left_0__2_
timestamp 1603810449
transform 1 0 19896 0 1 182824
box 0 0 16000 38752
use sb_0__1_  sb_0__1_
timestamp 1603810449
transform 1 0 48896 0 1 141824
box 0 0 28000 28000
use cby_0__1_  cby_0__2_
timestamp 1603810449
transform 1 0 54896 0 1 182824
box 0 0 16000 40000
use grid_clb  grid_clb_1__2_
timestamp 1603810449
transform 1 0 84896 0 1 177824
box 0 0 50000 50000
use cbx_1__1_  cbx_1__1_
timestamp 1603810449
transform 1 0 89896 0 1 147824
box 0 0 40000 16000
use sb_1__1_  sb_1__1_
timestamp 1603810449
transform 1 0 142896 0 1 141824
box 0 0 28000 28000
use cby_1__1_  cby_1__2_
timestamp 1603810449
transform 1 0 148896 0 1 182824
box 0 0 16000 40000
use grid_clb  grid_clb_2__2_
timestamp 1603810449
transform 1 0 178896 0 1 177824
box 0 0 50000 50000
use cbx_1__1_  cbx_2__1_
timestamp 1603810449
transform 1 0 183896 0 1 147824
box 0 0 40000 16000
use sb_1__1_  sb_2__1_
timestamp 1603810449
transform 1 0 236896 0 1 141824
box 0 0 28000 28000
use cby_1__1_  cby_2__2_
timestamp 1603810449
transform 1 0 242896 0 1 182824
box 0 0 16000 40000
use grid_clb  grid_clb_3__2_
timestamp 1603810449
transform 1 0 272896 0 1 177824
box 0 0 50000 50000
use cbx_1__1_  cbx_3__1_
timestamp 1603810449
transform 1 0 277896 0 1 147824
box 0 0 40000 16000
use sb_3__1_  sb_3__1_
timestamp 1603810449
transform 1 0 330896 0 1 141824
box 0 0 28000 28000
use cby_3__1_  cby_3__2_
timestamp 1603810449
transform 1 0 336896 0 1 182824
box 0 0 16000 40000
use grid_io_right  grid_io_right_4__2_
timestamp 1603810449
transform 1 0 408896 0 1 182824
box 0 0 16000 38752
use sb_0__1_  sb_0__2_
timestamp 1603810449
transform 1 0 48896 0 1 235824
box 0 0 28000 28000
use cbx_1__1_  cbx_1__2_
timestamp 1603810449
transform 1 0 89896 0 1 241824
box 0 0 40000 16000
use sb_1__1_  sb_1__2_
timestamp 1603810449
transform 1 0 142896 0 1 235824
box 0 0 28000 28000
use cbx_1__1_  cbx_2__2_
timestamp 1603810449
transform 1 0 183896 0 1 241824
box 0 0 40000 16000
use sb_1__1_  sb_2__2_
timestamp 1603810449
transform 1 0 236896 0 1 235824
box 0 0 28000 28000
use cbx_1__1_  cbx_3__2_
timestamp 1603810449
transform 1 0 277896 0 1 241824
box 0 0 40000 16000
use sb_3__1_  sb_3__2_
timestamp 1603810449
transform 1 0 330896 0 1 235824
box 0 0 28000 28000
use decoder6to61  decoder6to61_0_
timestamp 1603810449
transform 1 0 371896 0 1 212824
box 0 0 22854 24000
use grid_io_left  grid_io_left_0__3_
timestamp 1603810449
transform 1 0 19896 0 1 276824
box 0 0 16000 38752
use cby_0__1_  cby_0__3_
timestamp 1603810449
transform 1 0 54896 0 1 276824
box 0 0 16000 40000
use grid_clb  grid_clb_1__3_
timestamp 1603810449
transform 1 0 84896 0 1 271824
box 0 0 50000 50000
use cby_1__1_  cby_1__3_
timestamp 1603810449
transform 1 0 148896 0 1 276824
box 0 0 16000 40000
use grid_clb  grid_clb_2__3_
timestamp 1603810449
transform 1 0 178896 0 1 271824
box 0 0 50000 50000
use cby_1__1_  cby_2__3_
timestamp 1603810449
transform 1 0 242896 0 1 276824
box 0 0 16000 40000
use grid_clb  grid_clb_3__3_
timestamp 1603810449
transform 1 0 272896 0 1 271824
box 0 0 50000 50000
use cby_3__1_  cby_3__3_
timestamp 1603810449
transform 1 0 336896 0 1 276824
box 0 0 16000 40000
use grid_io_right  grid_io_right_4__3_
timestamp 1603810449
transform 1 0 408896 0 1 276824
box 0 0 16000 38752
use sb_0__3_  sb_0__3_
timestamp 1603810449
transform 1 0 48895 0 1 329824
box 1 0 27528 28000
use grid_io_top  grid_io_top_1__4_
timestamp 1603810449
transform 1 0 89896 0 1 370824
box 0 0 38934 16000
use cbx_1__3_  cbx_1__3_
timestamp 1603810449
transform 1 0 89896 0 1 335824
box 0 0 40000 16000
use sb_1__3_  sb_1__3_
timestamp 1603810449
transform 1 0 142896 0 1 329824
box 0 0 28000 27464
use grid_io_top  grid_io_top_2__4_
timestamp 1603810449
transform 1 0 183896 0 1 370824
box 0 0 38934 16000
use cbx_1__3_  cbx_2__3_
timestamp 1603810449
transform 1 0 183896 0 1 335824
box 0 0 40000 16000
use sb_1__3_  sb_2__3_
timestamp 1603810449
transform 1 0 236896 0 1 329824
box 0 0 28000 27464
use grid_io_top  grid_io_top_3__4_
timestamp 1603810449
transform 1 0 277896 0 1 370824
box 0 0 38934 16000
use cbx_1__3_  cbx_3__3_
timestamp 1603810449
transform 1 0 277896 0 1 335824
box 0 0 40000 16000
use sb_3__3_  sb_3__3_
timestamp 1603810449
transform 1 0 330896 0 1 329824
box 0 0 27587 27464
<< labels >>
rlabel metal2 s 231266 396344 231322 396824 6 address[0]
port 0 nsew default input
rlabel metal2 s 337526 396344 337582 396824 6 address[10]
port 1 nsew default input
rlabel metal2 s 355190 396344 355246 396824 6 address[11]
port 2 nsew default input
rlabel metal3 s 9896 336592 10376 336712 6 address[12]
port 3 nsew default input
rlabel metal2 s 351234 8824 351290 9304 6 address[13]
port 4 nsew default input
rlabel metal2 s 364114 8824 364170 9304 6 address[14]
port 5 nsew default input
rlabel metal3 s 434416 340400 434896 340520 6 address[15]
port 6 nsew default input
rlabel metal3 s 434416 315376 434896 315496 6 address[1]
port 7 nsew default input
rlabel metal2 s 325474 8824 325530 9304 6 address[2]
port 8 nsew default input
rlabel metal2 s 248930 396344 248986 396824 6 address[3]
port 9 nsew default input
rlabel metal2 s 338354 8824 338410 9304 6 address[4]
port 10 nsew default input
rlabel metal2 s 266686 396344 266742 396824 6 address[5]
port 11 nsew default input
rlabel metal2 s 284350 396344 284406 396824 6 address[6]
port 12 nsew default input
rlabel metal2 s 302106 396344 302162 396824 6 address[7]
port 13 nsew default input
rlabel metal3 s 434416 327888 434896 328008 6 address[8]
port 14 nsew default input
rlabel metal2 s 319770 396344 319826 396824 6 address[9]
port 15 nsew default input
rlabel metal3 s 434416 352912 434896 353032 6 clk
port 16 nsew default input
rlabel metal2 s 376994 8824 377050 9304 6 data_in
port 17 nsew default input
rlabel metal2 s 389874 8824 389930 9304 6 enable
port 18 nsew default input
rlabel metal2 s 18746 396344 18802 396824 6 gfpga_pad_GPIO_PAD[0]
port 19 nsew default bidirectional
rlabel metal2 s 89586 396344 89642 396824 6 gfpga_pad_GPIO_PAD[10]
port 20 nsew default bidirectional
rlabel metal2 s 107250 396344 107306 396824 6 gfpga_pad_GPIO_PAD[11]
port 21 nsew default bidirectional
rlabel metal2 s 125006 396344 125062 396824 6 gfpga_pad_GPIO_PAD[12]
port 22 nsew default bidirectional
rlabel metal2 s 142670 396344 142726 396824 6 gfpga_pad_GPIO_PAD[13]
port 23 nsew default bidirectional
rlabel metal2 s 402754 8824 402810 9304 6 gfpga_pad_GPIO_PAD[14]
port 24 nsew default bidirectional
rlabel metal2 s 415634 8824 415690 9304 6 gfpga_pad_GPIO_PAD[15]
port 25 nsew default bidirectional
rlabel metal3 s 434416 390448 434896 390568 6 gfpga_pad_GPIO_PAD[16]
port 26 nsew default bidirectional
rlabel metal3 s 9896 376712 10376 376832 6 gfpga_pad_GPIO_PAD[17]
port 27 nsew default bidirectional
rlabel metal2 s 408366 396344 408422 396824 6 gfpga_pad_GPIO_PAD[18]
port 28 nsew default bidirectional
rlabel metal2 s 426030 396344 426086 396824 6 gfpga_pad_GPIO_PAD[19]
port 29 nsew default bidirectional
rlabel metal2 s 36410 396344 36466 396824 6 gfpga_pad_GPIO_PAD[1]
port 30 nsew default bidirectional
rlabel metal2 s 160426 396344 160482 396824 6 gfpga_pad_GPIO_PAD[20]
port 31 nsew default bidirectional
rlabel metal2 s 178090 396344 178146 396824 6 gfpga_pad_GPIO_PAD[21]
port 32 nsew default bidirectional
rlabel metal2 s 195846 396344 195902 396824 6 gfpga_pad_GPIO_PAD[22]
port 33 nsew default bidirectional
rlabel metal2 s 213510 396344 213566 396824 6 gfpga_pad_GPIO_PAD[23]
port 34 nsew default bidirectional
rlabel metal3 s 434416 15088 434896 15208 6 gfpga_pad_GPIO_PAD[24]
port 35 nsew default bidirectional
rlabel metal3 s 434416 27600 434896 27720 6 gfpga_pad_GPIO_PAD[25]
port 36 nsew default bidirectional
rlabel metal3 s 434416 40112 434896 40232 6 gfpga_pad_GPIO_PAD[26]
port 37 nsew default bidirectional
rlabel metal3 s 434416 52624 434896 52744 6 gfpga_pad_GPIO_PAD[27]
port 38 nsew default bidirectional
rlabel metal3 s 434416 65136 434896 65256 6 gfpga_pad_GPIO_PAD[28]
port 39 nsew default bidirectional
rlabel metal3 s 434416 77648 434896 77768 6 gfpga_pad_GPIO_PAD[29]
port 40 nsew default bidirectional
rlabel metal2 s 54166 396344 54222 396824 6 gfpga_pad_GPIO_PAD[2]
port 41 nsew default bidirectional
rlabel metal3 s 434416 90160 434896 90280 6 gfpga_pad_GPIO_PAD[30]
port 42 nsew default bidirectional
rlabel metal3 s 434416 102672 434896 102792 6 gfpga_pad_GPIO_PAD[31]
port 43 nsew default bidirectional
rlabel metal3 s 434416 115184 434896 115304 6 gfpga_pad_GPIO_PAD[32]
port 44 nsew default bidirectional
rlabel metal3 s 434416 127696 434896 127816 6 gfpga_pad_GPIO_PAD[33]
port 45 nsew default bidirectional
rlabel metal3 s 434416 140208 434896 140328 6 gfpga_pad_GPIO_PAD[34]
port 46 nsew default bidirectional
rlabel metal3 s 434416 152720 434896 152840 6 gfpga_pad_GPIO_PAD[35]
port 47 nsew default bidirectional
rlabel metal3 s 434416 165232 434896 165352 6 gfpga_pad_GPIO_PAD[36]
port 48 nsew default bidirectional
rlabel metal3 s 434416 177744 434896 177864 6 gfpga_pad_GPIO_PAD[37]
port 49 nsew default bidirectional
rlabel metal3 s 434416 190256 434896 190376 6 gfpga_pad_GPIO_PAD[38]
port 50 nsew default bidirectional
rlabel metal3 s 434416 202768 434896 202888 6 gfpga_pad_GPIO_PAD[39]
port 51 nsew default bidirectional
rlabel metal2 s 71830 396344 71886 396824 6 gfpga_pad_GPIO_PAD[3]
port 52 nsew default bidirectional
rlabel metal3 s 434416 215280 434896 215400 6 gfpga_pad_GPIO_PAD[40]
port 53 nsew default bidirectional
rlabel metal3 s 434416 227792 434896 227912 6 gfpga_pad_GPIO_PAD[41]
port 54 nsew default bidirectional
rlabel metal3 s 434416 240304 434896 240424 6 gfpga_pad_GPIO_PAD[42]
port 55 nsew default bidirectional
rlabel metal3 s 434416 252816 434896 252936 6 gfpga_pad_GPIO_PAD[43]
port 56 nsew default bidirectional
rlabel metal3 s 434416 265328 434896 265448 6 gfpga_pad_GPIO_PAD[44]
port 57 nsew default bidirectional
rlabel metal3 s 434416 277840 434896 277960 6 gfpga_pad_GPIO_PAD[45]
port 58 nsew default bidirectional
rlabel metal3 s 434416 290352 434896 290472 6 gfpga_pad_GPIO_PAD[46]
port 59 nsew default bidirectional
rlabel metal3 s 434416 302864 434896 302984 6 gfpga_pad_GPIO_PAD[47]
port 60 nsew default bidirectional
rlabel metal2 s 16354 8824 16410 9304 6 gfpga_pad_GPIO_PAD[48]
port 61 nsew default bidirectional
rlabel metal2 s 29234 8824 29290 9304 6 gfpga_pad_GPIO_PAD[49]
port 62 nsew default bidirectional
rlabel metal2 s 372946 396344 373002 396824 6 gfpga_pad_GPIO_PAD[4]
port 63 nsew default bidirectional
rlabel metal2 s 42114 8824 42170 9304 6 gfpga_pad_GPIO_PAD[50]
port 64 nsew default bidirectional
rlabel metal2 s 54994 8824 55050 9304 6 gfpga_pad_GPIO_PAD[51]
port 65 nsew default bidirectional
rlabel metal2 s 67874 8824 67930 9304 6 gfpga_pad_GPIO_PAD[52]
port 66 nsew default bidirectional
rlabel metal2 s 80754 8824 80810 9304 6 gfpga_pad_GPIO_PAD[53]
port 67 nsew default bidirectional
rlabel metal2 s 93634 8824 93690 9304 6 gfpga_pad_GPIO_PAD[54]
port 68 nsew default bidirectional
rlabel metal2 s 106514 8824 106570 9304 6 gfpga_pad_GPIO_PAD[55]
port 69 nsew default bidirectional
rlabel metal2 s 119394 8824 119450 9304 6 gfpga_pad_GPIO_PAD[56]
port 70 nsew default bidirectional
rlabel metal2 s 132274 8824 132330 9304 6 gfpga_pad_GPIO_PAD[57]
port 71 nsew default bidirectional
rlabel metal2 s 145154 8824 145210 9304 6 gfpga_pad_GPIO_PAD[58]
port 72 nsew default bidirectional
rlabel metal2 s 158034 8824 158090 9304 6 gfpga_pad_GPIO_PAD[59]
port 73 nsew default bidirectional
rlabel metal3 s 9896 349920 10376 350040 6 gfpga_pad_GPIO_PAD[5]
port 74 nsew default bidirectional
rlabel metal2 s 170914 8824 170970 9304 6 gfpga_pad_GPIO_PAD[60]
port 75 nsew default bidirectional
rlabel metal2 s 183794 8824 183850 9304 6 gfpga_pad_GPIO_PAD[61]
port 76 nsew default bidirectional
rlabel metal2 s 196674 8824 196730 9304 6 gfpga_pad_GPIO_PAD[62]
port 77 nsew default bidirectional
rlabel metal2 s 209554 8824 209610 9304 6 gfpga_pad_GPIO_PAD[63]
port 78 nsew default bidirectional
rlabel metal2 s 222434 8824 222490 9304 6 gfpga_pad_GPIO_PAD[64]
port 79 nsew default bidirectional
rlabel metal2 s 235314 8824 235370 9304 6 gfpga_pad_GPIO_PAD[65]
port 80 nsew default bidirectional
rlabel metal2 s 248194 8824 248250 9304 6 gfpga_pad_GPIO_PAD[66]
port 81 nsew default bidirectional
rlabel metal2 s 261074 8824 261130 9304 6 gfpga_pad_GPIO_PAD[67]
port 82 nsew default bidirectional
rlabel metal2 s 273954 8824 274010 9304 6 gfpga_pad_GPIO_PAD[68]
port 83 nsew default bidirectional
rlabel metal2 s 286834 8824 286890 9304 6 gfpga_pad_GPIO_PAD[69]
port 84 nsew default bidirectional
rlabel metal3 s 434416 365424 434896 365544 6 gfpga_pad_GPIO_PAD[6]
port 85 nsew default bidirectional
rlabel metal2 s 299714 8824 299770 9304 6 gfpga_pad_GPIO_PAD[70]
port 86 nsew default bidirectional
rlabel metal2 s 312594 8824 312650 9304 6 gfpga_pad_GPIO_PAD[71]
port 87 nsew default bidirectional
rlabel metal3 s 9896 15496 10376 15616 6 gfpga_pad_GPIO_PAD[72]
port 88 nsew default bidirectional
rlabel metal3 s 9896 28824 10376 28944 6 gfpga_pad_GPIO_PAD[73]
port 89 nsew default bidirectional
rlabel metal3 s 9896 42152 10376 42272 6 gfpga_pad_GPIO_PAD[74]
port 90 nsew default bidirectional
rlabel metal3 s 9896 55616 10376 55736 6 gfpga_pad_GPIO_PAD[75]
port 91 nsew default bidirectional
rlabel metal3 s 9896 68944 10376 69064 6 gfpga_pad_GPIO_PAD[76]
port 92 nsew default bidirectional
rlabel metal3 s 9896 82272 10376 82392 6 gfpga_pad_GPIO_PAD[77]
port 93 nsew default bidirectional
rlabel metal3 s 9896 95736 10376 95856 6 gfpga_pad_GPIO_PAD[78]
port 94 nsew default bidirectional
rlabel metal3 s 9896 109064 10376 109184 6 gfpga_pad_GPIO_PAD[79]
port 95 nsew default bidirectional
rlabel metal2 s 390610 396344 390666 396824 6 gfpga_pad_GPIO_PAD[7]
port 96 nsew default bidirectional
rlabel metal3 s 9896 122528 10376 122648 6 gfpga_pad_GPIO_PAD[80]
port 97 nsew default bidirectional
rlabel metal3 s 9896 135856 10376 135976 6 gfpga_pad_GPIO_PAD[81]
port 98 nsew default bidirectional
rlabel metal3 s 9896 149184 10376 149304 6 gfpga_pad_GPIO_PAD[82]
port 99 nsew default bidirectional
rlabel metal3 s 9896 162648 10376 162768 6 gfpga_pad_GPIO_PAD[83]
port 100 nsew default bidirectional
rlabel metal3 s 9896 175976 10376 176096 6 gfpga_pad_GPIO_PAD[84]
port 101 nsew default bidirectional
rlabel metal3 s 9896 189304 10376 189424 6 gfpga_pad_GPIO_PAD[85]
port 102 nsew default bidirectional
rlabel metal3 s 9896 202768 10376 202888 6 gfpga_pad_GPIO_PAD[86]
port 103 nsew default bidirectional
rlabel metal3 s 9896 216096 10376 216216 6 gfpga_pad_GPIO_PAD[87]
port 104 nsew default bidirectional
rlabel metal3 s 9896 229560 10376 229680 6 gfpga_pad_GPIO_PAD[88]
port 105 nsew default bidirectional
rlabel metal3 s 9896 242888 10376 243008 6 gfpga_pad_GPIO_PAD[89]
port 106 nsew default bidirectional
rlabel metal3 s 434416 377936 434896 378056 6 gfpga_pad_GPIO_PAD[8]
port 107 nsew default bidirectional
rlabel metal3 s 9896 256216 10376 256336 6 gfpga_pad_GPIO_PAD[90]
port 108 nsew default bidirectional
rlabel metal3 s 9896 269680 10376 269800 6 gfpga_pad_GPIO_PAD[91]
port 109 nsew default bidirectional
rlabel metal3 s 9896 283008 10376 283128 6 gfpga_pad_GPIO_PAD[92]
port 110 nsew default bidirectional
rlabel metal3 s 9896 296336 10376 296456 6 gfpga_pad_GPIO_PAD[93]
port 111 nsew default bidirectional
rlabel metal3 s 9896 309800 10376 309920 6 gfpga_pad_GPIO_PAD[94]
port 112 nsew default bidirectional
rlabel metal3 s 9896 323128 10376 323248 6 gfpga_pad_GPIO_PAD[95]
port 113 nsew default bidirectional
rlabel metal3 s 9896 363248 10376 363368 6 gfpga_pad_GPIO_PAD[9]
port 114 nsew default bidirectional
rlabel metal3 s 9896 390040 10376 390160 6 reset
port 115 nsew default input
rlabel metal2 s 428514 8824 428570 9304 6 set
port 116 nsew default input
rlabel metal5 s 5000 5000 439740 9000 8 vpwr
port 117 nsew default input
rlabel metal5 s 0 0 444740 4000 8 vgnd
port 118 nsew default input
<< properties >>
string FIXED_BBOX 0 0 444740 405520
<< end >>
