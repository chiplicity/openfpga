* NGSPICE file created from sb_0__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

.subckt sb_0__1_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] bottom_left_grid_pin_11_ bottom_left_grid_pin_13_ bottom_left_grid_pin_15_
+ bottom_left_grid_pin_1_ bottom_left_grid_pin_3_ bottom_left_grid_pin_5_ bottom_left_grid_pin_7_
+ bottom_left_grid_pin_9_ bottom_right_grid_pin_11_ chanx_right_in[0] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chany_bottom_in[0] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_out[0] chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3]
+ chany_bottom_out[4] chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7]
+ chany_bottom_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ right_bottom_grid_pin_12_ right_top_grid_pin_10_ top_left_grid_pin_11_ top_left_grid_pin_13_
+ top_left_grid_pin_15_ top_left_grid_pin_1_ top_left_grid_pin_3_ top_left_grid_pin_5_
+ top_left_grid_pin_7_ top_left_grid_pin_9_ top_right_grid_pin_11_ vpwr vgnd
Xmem_right_track_12.LATCH_1_.latch data_in _181_/A _167_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_177 vgnd vpwr scs8hd_decap_8
XFILLER_22_111 vpwr vgnd scs8hd_fill_2
XFILLER_22_100 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_52 vgnd vpwr scs8hd_fill_1
XFILLER_13_100 vgnd vpwr scs8hd_decap_3
XFILLER_9_115 vpwr vgnd scs8hd_fill_2
XFILLER_13_166 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__113__B _109_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_3_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _181_/A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__214__A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_37_51 vgnd vpwr scs8hd_decap_8
XANTENNA__108__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _113_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _194_/HI _176_/Y mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_184 vpwr vgnd scs8hd_fill_2
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _188_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_4.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_200_ _200_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__209__A _209_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_206 vpwr vgnd scs8hd_fill_2
XFILLER_15_239 vgnd vpwr scs8hd_decap_3
X_131_ _110_/A _134_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_132 vpwr vgnd scs8hd_fill_2
XFILLER_0_68 vpwr vgnd scs8hd_fill_2
XFILLER_9_88 vpwr vgnd scs8hd_fill_2
XFILLER_14_250 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _139_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _213_/A vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_17.LATCH_2_.latch data_in mem_bottom_track_17.LATCH_2_.latch/Q _151_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_114_ address[4] _115_/B vgnd vpwr scs8hd_inv_8
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_7_ mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__121__B _118_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XANTENNA__222__A _222_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_74 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[6] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_23 vgnd vpwr scs8hd_decap_8
XANTENNA__132__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_67 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_1_.latch data_in _183_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_208 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XANTENNA__217__A _217_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_43 vgnd vpwr scs8hd_decap_6
XFILLER_31_97 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ _178_/A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_123 vpwr vgnd scs8hd_fill_2
XFILLER_31_101 vpwr vgnd scs8hd_fill_2
XANTENNA__127__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_131 vgnd vpwr scs8hd_decap_4
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_201 vpwr vgnd scs8hd_fill_2
XFILLER_39_245 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _188_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_167 vgnd vpwr scs8hd_fill_1
XFILLER_22_145 vgnd vpwr scs8hd_decap_3
Xmux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _191_/HI _182_/Y mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_105 vpwr vgnd scs8hd_fill_2
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_3_68 vpwr vgnd scs8hd_fill_2
XFILLER_3_57 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_259 vgnd vpwr scs8hd_decap_12
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _195_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_171 vgnd vpwr scs8hd_decap_8
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_27_259 vpwr vgnd scs8hd_fill_2
XFILLER_12_88 vgnd vpwr scs8hd_decap_4
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__124__B _118_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _109_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_1_ vgnd vpwr scs8hd_diode_2
XFILLER_17_270 vgnd vpwr scs8hd_decap_6
XFILLER_32_251 vgnd vpwr scs8hd_decap_4
X_130_ _109_/A _134_/B _130_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_15_229 vgnd vpwr scs8hd_decap_4
XANTENNA__225__A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_36 vpwr vgnd scs8hd_fill_2
XFILLER_0_47 vpwr vgnd scs8hd_fill_2
XFILLER_0_58 vgnd vpwr scs8hd_decap_4
XANTENNA__119__B _118_/X vgnd vpwr scs8hd_diode_2
XANTENNA__135__A _104_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_232 vgnd vpwr scs8hd_fill_1
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_214 vgnd vpwr scs8hd_decap_4
XFILLER_7_236 vpwr vgnd scs8hd_fill_2
XFILLER_11_232 vpwr vgnd scs8hd_fill_2
XFILLER_11_265 vpwr vgnd scs8hd_fill_2
X_113_ _113_/A _109_/B _113_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_15_7 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _186_/A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_88 vpwr vgnd scs8hd_fill_2
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_86 vgnd vpwr scs8hd_decap_6
XANTENNA__132__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_19_162 vpwr vgnd scs8hd_fill_2
XFILLER_19_140 vpwr vgnd scs8hd_fill_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XFILLER_34_143 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_187 vpwr vgnd scs8hd_fill_2
XFILLER_25_165 vpwr vgnd scs8hd_fill_2
XFILLER_15_66 vpwr vgnd scs8hd_fill_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_3
XFILLER_31_146 vpwr vgnd scs8hd_fill_2
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _167_/B vgnd vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_165 vpwr vgnd scs8hd_fill_2
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_235 vgnd vpwr scs8hd_decap_8
XFILLER_22_157 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.INVTX1_2_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _209_/A vgnd vpwr scs8hd_inv_1
XFILLER_3_36 vpwr vgnd scs8hd_fill_2
XFILLER_3_25 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A _137_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_194 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_105 vgnd vpwr scs8hd_decap_8
XFILLER_12_67 vpwr vgnd scs8hd_fill_2
XFILLER_5_6 vpwr vgnd scs8hd_fill_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_41_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__140__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_1_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_88 vpwr vgnd scs8hd_fill_2
XFILLER_23_77 vpwr vgnd scs8hd_fill_2
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_178 vpwr vgnd scs8hd_fill_2
XFILLER_2_167 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_35 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_12.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr
+ scs8hd_diode_2
XANTENNA__135__B _115_/B vgnd vpwr scs8hd_diode_2
X_189_ _189_/HI _189_/LO vgnd vpwr scs8hd_conb_1
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_211 vgnd vpwr scs8hd_decap_3
XFILLER_18_44 vgnd vpwr scs8hd_decap_8
XFILLER_34_32 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_88 vpwr vgnd scs8hd_fill_2
XFILLER_7_259 vgnd vpwr scs8hd_decap_4
X_112_ _123_/A _109_/B _112_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_211 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__146__A _160_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_80 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _173_/A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_20_67 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_207 vgnd vpwr scs8hd_fill_1
XFILLER_28_163 vgnd vpwr scs8hd_decap_3
XFILLER_3_262 vpwr vgnd scs8hd_fill_2
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_144 vpwr vgnd scs8hd_fill_2
XFILLER_0_265 vpwr vgnd scs8hd_fill_2
XFILLER_0_221 vpwr vgnd scs8hd_fill_2
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__C _170_/C vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_188 vpwr vgnd scs8hd_fill_2
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__143__B _139_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_214 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
Xmem_right_track_4.LATCH_1_.latch data_in _175_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_2.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
XFILLER_26_66 vgnd vpwr scs8hd_fill_1
XFILLER_26_44 vgnd vpwr scs8hd_decap_8
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_88 vpwr vgnd scs8hd_fill_2
XFILLER_13_114 vpwr vgnd scs8hd_fill_2
XFILLER_13_147 vpwr vgnd scs8hd_fill_2
Xmux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _177_/Y mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_4
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__154__A _117_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_14.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_128 vgnd vpwr scs8hd_decap_6
XFILLER_12_46 vgnd vpwr scs8hd_decap_8
XFILLER_18_206 vgnd vpwr scs8hd_decap_6
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_228 vgnd vpwr scs8hd_decap_4
XFILLER_41_275 vpwr vgnd scs8hd_fill_2
XFILLER_41_253 vpwr vgnd scs8hd_fill_2
XFILLER_5_121 vgnd vpwr scs8hd_fill_1
XFILLER_5_154 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _101_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A _109_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_3_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XFILLER_23_242 vpwr vgnd scs8hd_fill_2
XFILLER_23_56 vgnd vpwr scs8hd_decap_3
XFILLER_2_113 vpwr vgnd scs8hd_fill_2
XFILLER_2_102 vgnd vpwr scs8hd_decap_3
XFILLER_0_16 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_9_47 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__135__C _104_/C vgnd vpwr scs8hd_diode_2
X_188_ _188_/HI _188_/LO vgnd vpwr scs8hd_conb_1
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _179_/A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__151__B _149_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _193_/HI _174_/Y mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_67 vpwr vgnd scs8hd_fill_2
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
XFILLER_34_99 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_11_245 vpwr vgnd scs8hd_fill_2
X_111_ _122_/A _109_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__B _125_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _164_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_29_66 vpwr vgnd scs8hd_fill_2
XFILLER_28_131 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _196_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_15 vgnd vpwr scs8hd_decap_4
XFILLER_3_274 vgnd vpwr scs8hd_decap_3
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _159_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_197 vgnd vpwr scs8hd_decap_4
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_2_.latch data_in mem_bottom_track_1.LATCH_2_.latch/Q _132_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _192_/HI _185_/Y mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
XFILLER_15_57 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_112 vgnd vpwr scs8hd_decap_8
XFILLER_16_145 vgnd vpwr scs8hd_decap_6
XFILLER_31_159 vpwr vgnd scs8hd_fill_2
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_259 vpwr vgnd scs8hd_fill_2
XFILLER_39_226 vgnd vpwr scs8hd_fill_1
XFILLER_22_115 vpwr vgnd scs8hd_fill_2
XFILLER_22_104 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_80 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_119 vgnd vpwr scs8hd_decap_3
XFILLER_13_126 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ _176_/A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_181 vgnd vpwr scs8hd_decap_3
XANTENNA__170__A _160_/A vgnd vpwr scs8hd_diode_2
XANTENNA__080__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _190_/HI _180_/Y mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_188 vgnd vpwr scs8hd_decap_3
XANTENNA__149__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_251 vpwr vgnd scs8hd_fill_2
XFILLER_17_262 vpwr vgnd scs8hd_fill_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _164_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_210 vgnd vpwr scs8hd_decap_12
XANTENNA__075__A address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_0_.scs8hd_inv_1 chany_top_in[6] mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_136 vpwr vgnd scs8hd_fill_2
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_254 vgnd vpwr scs8hd_decap_4
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/HI _187_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_180 vgnd vpwr scs8hd_fill_1
XFILLER_20_224 vgnd vpwr scs8hd_decap_8
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _184_/Y mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
X_110_ _110_/A _109_/B _110_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__146__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _164_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_143 vpwr vgnd scs8hd_fill_2
XFILLER_3_242 vpwr vgnd scs8hd_fill_2
XFILLER_6_38 vgnd vpwr scs8hd_fill_1
XANTENNA__157__B _164_/B vgnd vpwr scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ _182_/A mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__083__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_127 vgnd vpwr scs8hd_decap_4
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_135 vgnd vpwr scs8hd_fill_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_205 vgnd vpwr scs8hd_decap_4
XFILLER_39_249 vgnd vpwr scs8hd_decap_6
XANTENNA__168__A _159_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_271 vgnd vpwr scs8hd_decap_4
XFILLER_26_79 vgnd vpwr scs8hd_decap_3
XANTENNA__078__A _077_/X vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_1_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_193 vpwr vgnd scs8hd_fill_2
XFILLER_21_171 vpwr vgnd scs8hd_fill_2
XFILLER_9_109 vgnd vpwr scs8hd_decap_4
XFILLER_16_90 vpwr vgnd scs8hd_fill_2
XANTENNA__170__B _165_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_5_123 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_1_.latch data_in mem_top_track_8.LATCH_1_.latch/Q _112_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_211 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__165__B _165_/B vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_71 vpwr vgnd scs8hd_fill_2
XFILLER_23_222 vgnd vpwr scs8hd_decap_12
XANTENNA__091__A _090_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_27 vgnd vpwr scs8hd_decap_8
XFILLER_14_233 vpwr vgnd scs8hd_fill_2
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_91 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_170 vgnd vpwr scs8hd_decap_4
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_258 vgnd vpwr scs8hd_decap_12
XFILLER_20_247 vgnd vpwr scs8hd_decap_8
XFILLER_20_236 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_5_ mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_7_218 vgnd vpwr scs8hd_fill_1
XFILLER_11_236 vpwr vgnd scs8hd_fill_2
XFILLER_11_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_3 vgnd vpwr scs8hd_decap_6
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__162__C _161_/C vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.INVTX1_0_.scs8hd_inv_1 chany_top_in[5] mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_169_ _160_/A _165_/B _170_/C _163_/D _169_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_114 vgnd vpwr scs8hd_decap_12
XFILLER_34_103 vpwr vgnd scs8hd_fill_2
XFILLER_19_144 vgnd vpwr scs8hd_decap_3
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XANTENNA__157__C _159_/C vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_3_.latch data_in mem_bottom_track_9.LATCH_3_.latch/Q _141_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_114 vpwr vgnd scs8hd_fill_2
XANTENNA__083__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_0_213 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_169 vgnd vpwr scs8hd_decap_4
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__168__B _167_/B vgnd vpwr scs8hd_diode_2
XFILLER_22_128 vpwr vgnd scs8hd_fill_2
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XFILLER_26_69 vgnd vpwr scs8hd_fill_1
XANTENNA__094__A _093_/X vgnd vpwr scs8hd_diode_2
XFILLER_21_161 vgnd vpwr scs8hd_fill_1
XFILLER_3_29 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_132 vpwr vgnd scs8hd_fill_2
XFILLER_8_154 vpwr vgnd scs8hd_fill_2
XFILLER_12_150 vgnd vpwr scs8hd_fill_1
XANTENNA__170__C _170_/C vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_253 vpwr vgnd scs8hd_fill_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.tap_buf4_0_.scs8hd_inv_1 mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ _202_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _149_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__089__A address[1] vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_245 vgnd vpwr scs8hd_decap_8
XFILLER_5_135 vpwr vgnd scs8hd_fill_2
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
XFILLER_17_231 vpwr vgnd scs8hd_fill_2
XANTENNA__165__C _159_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _175_/Y mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_50 vgnd vpwr scs8hd_decap_6
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XFILLER_23_234 vgnd vpwr scs8hd_decap_8
XFILLER_23_15 vgnd vpwr scs8hd_decap_12
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_14_212 vpwr vgnd scs8hd_fill_2
XFILLER_14_267 vgnd vpwr scs8hd_decap_8
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
Xmux_right_track_6.INVTX1_1_.scs8hd_inv_1 chany_top_in[8] mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_193 vpwr vgnd scs8hd_fill_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XANTENNA__086__B _086_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__162__D _164_/D vgnd vpwr scs8hd_diode_2
XFILLER_6_230 vpwr vgnd scs8hd_fill_2
X_168_ _159_/A _167_/B _161_/C _164_/D _168_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
X_099_ address[1] address[2] address[0] _099_/X vgnd vpwr scs8hd_or3_4
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
XFILLER_1_40 vpwr vgnd scs8hd_fill_2
XFILLER_1_62 vgnd vpwr scs8hd_decap_3
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_112 vgnd vpwr scs8hd_decap_6
XANTENNA__097__A _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_266 vgnd vpwr scs8hd_decap_8
XFILLER_10_93 vgnd vpwr scs8hd_decap_3
XFILLER_34_126 vgnd vpwr scs8hd_fill_1
XFILLER_19_112 vgnd vpwr scs8hd_decap_4
XFILLER_19_91 vpwr vgnd scs8hd_fill_2
XANTENNA__157__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_159 vgnd vpwr scs8hd_decap_4
XFILLER_15_49 vgnd vpwr scs8hd_fill_1
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XANTENNA__083__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
XFILLER_0_225 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_17.LATCH_3_.latch data_in mem_bottom_track_17.LATCH_3_.latch/Q _150_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_31_118 vpwr vgnd scs8hd_fill_2
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_81 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_218 vgnd vpwr scs8hd_decap_8
XFILLER_11_6 vpwr vgnd scs8hd_fill_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XANTENNA__168__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_251 vgnd vpwr scs8hd_decap_4
Xmux_right_track_6.tap_buf4_0_.scs8hd_inv_1 mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ _205_/A vgnd vpwr scs8hd_inv_1
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_118 vgnd vpwr scs8hd_decap_4
Xmux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _181_/Y mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_19 vgnd vpwr scs8hd_fill_1
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_122 vgnd vpwr scs8hd_decap_8
XFILLER_12_140 vpwr vgnd scs8hd_fill_2
XANTENNA__170__D _164_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_5_114 vgnd vpwr scs8hd_decap_4
XFILLER_5_158 vpwr vgnd scs8hd_fill_2
XFILLER_17_210 vgnd vpwr scs8hd_decap_4
XFILLER_27_80 vpwr vgnd scs8hd_fill_2
XANTENNA__165__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_17_243 vgnd vpwr scs8hd_fill_1
XFILLER_17_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_84 vgnd vpwr scs8hd_decap_4
Xmux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _174_/A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_0_.latch_SLEEPB _166_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_27 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_2_117 vpwr vgnd scs8hd_fill_2
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA__086__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_11_249 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_167_ _159_/A _167_/B _161_/C _163_/D _167_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_242 vgnd vpwr scs8hd_decap_4
X_098_ _095_/A _123_/A _098_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_260 vgnd vpwr scs8hd_decap_12
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
Xmux_right_track_4.INVTX1_1_.scs8hd_inv_1 chany_top_in[7] mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_168 vgnd vpwr scs8hd_decap_3
XFILLER_28_135 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ _178_/Y mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vpwr vgnd scs8hd_fill_2
XFILLER_3_234 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_19 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_138 vpwr vgnd scs8hd_fill_2
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
X_219_ chany_bottom_in[6] chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_33_182 vgnd vpwr scs8hd_fill_1
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_138 vpwr vgnd scs8hd_fill_2
XFILLER_24_193 vgnd vpwr scs8hd_decap_12
XFILLER_24_182 vpwr vgnd scs8hd_fill_2
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _198_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_130 vgnd vpwr scs8hd_decap_3
XPHY_2 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_182 vgnd vpwr scs8hd_fill_1
XANTENNA__168__D _164_/D vgnd vpwr scs8hd_diode_2
XFILLER_30_163 vgnd vpwr scs8hd_decap_12
XFILLER_30_152 vgnd vpwr scs8hd_fill_1
XFILLER_7_40 vpwr vgnd scs8hd_fill_2
XFILLER_7_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_82 vpwr vgnd scs8hd_fill_2
XFILLER_16_93 vpwr vgnd scs8hd_fill_2
Xmux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_0_.scs8hd_inv_1/Y
+ _180_/A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_8_112 vgnd vpwr scs8hd_fill_1
XFILLER_8_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_7_ vgnd vpwr scs8hd_diode_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_37_59 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_255 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_266 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XFILLER_23_39 vgnd vpwr scs8hd_decap_12
XFILLER_2_107 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_184 vgnd vpwr scs8hd_fill_1
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_240 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _186_/Y mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_217 vpwr vgnd scs8hd_fill_2
XFILLER_11_228 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_11_ mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_93 vgnd vpwr scs8hd_decap_3
XFILLER_24_82 vgnd vpwr scs8hd_decap_4
XFILLER_6_210 vgnd vpwr scs8hd_decap_4
X_166_ _164_/A _165_/B _159_/C _164_/D _166_/Y vgnd vpwr scs8hd_nor4_4
X_097_ _096_/X _123_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
XFILLER_10_272 vgnd vpwr scs8hd_decap_3
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XFILLER_1_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _140_/Y vgnd vpwr scs8hd_diode_2
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_28_147 vgnd vpwr scs8hd_decap_6
XFILLER_3_202 vpwr vgnd scs8hd_fill_2
XFILLER_19_60 vgnd vpwr scs8hd_fill_1
XFILLER_10_84 vpwr vgnd scs8hd_fill_2
XFILLER_35_92 vpwr vgnd scs8hd_fill_2
XFILLER_19_158 vpwr vgnd scs8hd_fill_2
X_218_ _218_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
X_149_ _109_/A _149_/B _149_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_191 vpwr vgnd scs8hd_fill_2
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XFILLER_0_249 vgnd vpwr scs8hd_decap_3
XFILLER_0_238 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_24_150 vgnd vpwr scs8hd_decap_3
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_39_209 vgnd vpwr scs8hd_fill_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_175 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _189_/HI mem_bottom_track_9.LATCH_2_.latch/Q
+ mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_197 vgnd vpwr scs8hd_decap_4
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XFILLER_21_153 vpwr vgnd scs8hd_fill_2
XFILLER_21_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_186 vgnd vpwr scs8hd_decap_3
XFILLER_35_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_27 vgnd vpwr scs8hd_decap_12
XFILLER_26_201 vgnd vpwr scs8hd_decap_12
XFILLER_41_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_93 vgnd vpwr scs8hd_decap_4
XFILLER_17_245 vgnd vpwr scs8hd_decap_3
XFILLER_32_259 vgnd vpwr scs8hd_decap_12
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _134_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_171 vgnd vpwr scs8hd_decap_8
XFILLER_4_193 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_215 vpwr vgnd scs8hd_fill_2
XFILLER_14_237 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_62 vgnd vpwr scs8hd_decap_3
XANTENNA__100__A _099_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_15_ mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ _173_/Y mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_165_ _164_/A _165_/B _159_/C _163_/D _165_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ address[1] address[2] _156_/A _096_/X vgnd vpwr scs8hd_or3_4
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
XFILLER_1_76 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _098_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_72 vpwr vgnd scs8hd_fill_2
XFILLER_34_107 vgnd vpwr scs8hd_decap_4
X_217_ _217_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
X_148_ _139_/A _149_/B _148_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
X_079_ address[5] _117_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_right_track_4.INVTX1_1_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_25_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_19 vgnd vpwr scs8hd_decap_12
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XFILLER_33_162 vgnd vpwr scs8hd_decap_12
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vpwr vgnd scs8hd_fill_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_187 vgnd vpwr scs8hd_decap_12
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_151 vgnd vpwr scs8hd_fill_1
XFILLER_15_195 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vgnd vpwr scs8hd_decap_3
XFILLER_7_97 vpwr vgnd scs8hd_fill_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_121 vgnd vpwr scs8hd_fill_1
XFILLER_21_110 vgnd vpwr scs8hd_fill_1
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XFILLER_12_154 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _152_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_158 vgnd vpwr scs8hd_decap_4
XANTENNA__103__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_14.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr
+ scs8hd_diode_2
XFILLER_37_39 vgnd vpwr scs8hd_decap_12
XFILLER_26_213 vgnd vpwr scs8hd_fill_1
XFILLER_5_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_3_.latch data_in mem_bottom_track_1.LATCH_3_.latch/Q _131_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_235 vpwr vgnd scs8hd_fill_2
XFILLER_40_271 vgnd vpwr scs8hd_decap_4
Xmux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ _179_/Y mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_22_271 vgnd vpwr scs8hd_decap_4
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_74 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
Xmem_right_track_14.LATCH_0_.latch data_in _186_/A _172_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XFILLER_1_153 vpwr vgnd scs8hd_fill_2
XFILLER_13_260 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
X_164_ _164_/A _164_/B _163_/C _164_/D _164_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_234 vgnd vpwr scs8hd_decap_4
XFILLER_10_230 vgnd vpwr scs8hd_decap_4
X_095_ _095_/A _122_/A _095_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__111__A _122_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_138 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_12.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_078_ _077_/X _139_/A vgnd vpwr scs8hd_buf_1
X_216_ chany_top_in[0] chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_147_ _146_/X _149_/B vgnd vpwr scs8hd_buf_1
XANTENNA__106__A _117_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_130 vpwr vgnd scs8hd_fill_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XFILLER_33_174 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_85 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
Xmux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_1_.scs8hd_inv_1/Y
+ _176_/Y mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_30_199 vgnd vpwr scs8hd_decap_12
XFILLER_30_122 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_163 vpwr vgnd scs8hd_fill_2
XFILLER_15_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_30 vgnd vpwr scs8hd_fill_1
XFILLER_16_52 vpwr vgnd scs8hd_fill_2
XFILLER_8_104 vpwr vgnd scs8hd_fill_2
XFILLER_12_100 vgnd vpwr scs8hd_decap_4
XFILLER_12_144 vgnd vpwr scs8hd_decap_6
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_118 vgnd vpwr scs8hd_fill_1
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_62 vgnd vpwr scs8hd_decap_3
XFILLER_17_214 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_6.LATCH_0_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_88 vgnd vpwr scs8hd_fill_1
XFILLER_4_140 vgnd vpwr scs8hd_decap_3
XFILLER_4_184 vgnd vpwr scs8hd_decap_3
XANTENNA__114__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_42 vgnd vpwr scs8hd_decap_6
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_13_97 vgnd vpwr scs8hd_fill_1
XFILLER_1_176 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_254 vpwr vgnd scs8hd_fill_2
XFILLER_9_265 vpwr vgnd scs8hd_fill_2
XFILLER_24_63 vgnd vpwr scs8hd_decap_6
XFILLER_24_52 vpwr vgnd scs8hd_fill_2
X_163_ _164_/A _164_/B _163_/C _163_/D _163_/Y vgnd vpwr scs8hd_nor4_4
X_094_ _093_/X _122_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_202 vpwr vgnd scs8hd_fill_2
XANTENNA__111__B _109_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _199_/HI vgnd vpwr
+ scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch data_in mem_top_track_8.LATCH_2_.latch/Q _111_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd
+ vpwr scs8hd_diode_2
Xmux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ _182_/Y mux_right_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_3_249 vpwr vgnd scs8hd_fill_2
XFILLER_3_238 vpwr vgnd scs8hd_fill_2
XANTENNA__212__A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_10_32 vpwr vgnd scs8hd_fill_2
XFILLER_10_65 vpwr vgnd scs8hd_fill_2
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_215_ chany_top_in[1] chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
X_077_ address[1] _086_/B _156_/A _077_/X vgnd vpwr scs8hd_or3_4
X_146_ _160_/A _125_/Y _161_/C _146_/X vgnd vpwr scs8hd_or3_4
XANTENNA__106__B _165_/B vgnd vpwr scs8hd_diode_2
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_161 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_186 vgnd vpwr scs8hd_decap_4
XFILLER_24_142 vgnd vpwr scs8hd_decap_6
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_30_145 vgnd vpwr scs8hd_decap_4
XANTENNA__117__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
X_129_ _139_/A _134_/B _129_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_21_123 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XFILLER_16_86 vpwr vgnd scs8hd_fill_2
XFILLER_8_149 vgnd vpwr scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_7_182 vgnd vpwr scs8hd_fill_1
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_9.LATCH_4_.latch data_in mem_bottom_track_9.LATCH_4_.latch/Q _140_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__220__A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _190_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__130__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_67 vpwr vgnd scs8hd_fill_2
XFILLER_4_23 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_251 vgnd vpwr scs8hd_decap_4
XANTENNA__215__A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XANTENNA__109__B _109_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_200 vpwr vgnd scs8hd_fill_2
XFILLER_9_222 vgnd vpwr scs8hd_decap_3
XFILLER_13_240 vpwr vgnd scs8hd_fill_2
XANTENNA__125__A address[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 bottom_left_grid_pin_9_ mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _143_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_170 vpwr vgnd scs8hd_fill_2
X_162_ _164_/A _164_/B _161_/C _164_/D _162_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_10_243 vpwr vgnd scs8hd_fill_2
X_093_ _093_/A address[2] address[0] _093_/X vgnd vpwr scs8hd_or3_4
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_10.LATCH_0_.latch data_in _180_/A _166_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_19_53 vgnd vpwr scs8hd_decap_4
XFILLER_10_88 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_162 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
XFILLER_35_96 vpwr vgnd scs8hd_fill_2
X_214_ chany_top_in[2] chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
X_145_ address[5] _160_/A vgnd vpwr scs8hd_inv_8
XANTENNA__106__C _163_/C vgnd vpwr scs8hd_diode_2
X_076_ address[0] _156_/A vgnd vpwr scs8hd_inv_8
XANTENNA__122__B _118_/X vgnd vpwr scs8hd_diode_2
XFILLER_18_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_195 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_165 vgnd vpwr scs8hd_decap_8
XFILLER_21_10 vgnd vpwr scs8hd_decap_12
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__223__A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_21_98 vpwr vgnd scs8hd_fill_2
XFILLER_30_135 vgnd vpwr scs8hd_fill_1
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_110 vpwr vgnd scs8hd_fill_2
XFILLER_15_132 vgnd vpwr scs8hd_decap_6
XFILLER_15_143 vpwr vgnd scs8hd_fill_2
X_128_ _127_/X _134_/B vgnd vpwr scs8hd_buf_1
XANTENNA__133__A _123_/A vgnd vpwr scs8hd_diode_2
XANTENNA__117__B address[6] vgnd vpwr scs8hd_diode_2
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XFILLER_23_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XFILLER_21_157 vpwr vgnd scs8hd_fill_2
XFILLER_21_146 vpwr vgnd scs8hd_fill_2
XFILLER_21_102 vgnd vpwr scs8hd_decap_6
Xmux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XANTENNA__218__A _218_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_16_65 vpwr vgnd scs8hd_fill_2
XFILLER_12_168 vgnd vpwr scs8hd_decap_8
XANTENNA__128__A _127_/X vgnd vpwr scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_17_227 vpwr vgnd scs8hd_fill_2
XANTENNA__130__B _134_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_bottom_track_17.LATCH_4_.latch data_in mem_bottom_track_17.LATCH_4_.latch/Q _149_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_219 vgnd vpwr scs8hd_decap_3
XFILLER_1_189 vpwr vgnd scs8hd_fill_2
XFILLER_1_101 vpwr vgnd scs8hd_fill_2
XFILLER_1_134 vpwr vgnd scs8hd_fill_2
Xmem_right_track_6.LATCH_0_.latch data_in _178_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__141__A _110_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_193 vgnd vpwr scs8hd_decap_4
XFILLER_39_182 vgnd vpwr scs8hd_fill_1
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
X_161_ _164_/A _164_/B _161_/C _163_/D _161_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_226 vpwr vgnd scs8hd_fill_2
XFILLER_6_248 vpwr vgnd scs8hd_fill_2
XFILLER_6_259 vgnd vpwr scs8hd_decap_12
X_092_ _095_/A _110_/A _092_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_1_14 vpwr vgnd scs8hd_fill_2
XFILLER_1_25 vgnd vpwr scs8hd_decap_6
XFILLER_1_36 vpwr vgnd scs8hd_fill_2
XANTENNA__136__A _136_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_152 vgnd vpwr scs8hd_fill_1
XFILLER_19_87 vpwr vgnd scs8hd_fill_2
XFILLER_19_65 vgnd vpwr scs8hd_decap_4
XFILLER_35_86 vgnd vpwr scs8hd_decap_3
Xmux_right_track_12.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_075_ address[2] _086_/B vgnd vpwr scs8hd_inv_8
X_213_ _213_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
X_144_ _113_/A _139_/B _144_/Y vgnd vpwr scs8hd_nor2_4
Xmux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _199_/HI mem_top_track_8.LATCH_2_.latch/Q
+ mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_2.tap_buf4_0_.scs8hd_inv_1 mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _207_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_273 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_174 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_1_ mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_22 vgnd vpwr scs8hd_decap_12
XFILLER_21_66 vgnd vpwr scs8hd_decap_4
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_15_199 vpwr vgnd scs8hd_fill_2
XANTENNA__117__C _170_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
X_127_ _117_/A _167_/B _170_/C _127_/X vgnd vpwr scs8hd_or3_4
XANTENNA__133__B _134_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _217_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[2] mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XFILLER_12_136 vpwr vgnd scs8hd_fill_2
XFILLER_16_44 vgnd vpwr scs8hd_decap_8
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA__144__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_180 vgnd vpwr scs8hd_decap_3
XFILLER_7_195 vgnd vpwr scs8hd_decap_3
Xmux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _174_/Y mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_76 vpwr vgnd scs8hd_fill_2
XFILLER_17_217 vgnd vpwr scs8hd_fill_1
XFILLER_17_239 vgnd vpwr scs8hd_decap_4
XFILLER_4_121 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vpwr vgnd scs8hd_fill_2
XFILLER_31_253 vpwr vgnd scs8hd_fill_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _139_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_78 vpwr vgnd scs8hd_fill_2
XFILLER_1_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__141__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_88 vpwr vgnd scs8hd_fill_2
XFILLER_24_44 vgnd vpwr scs8hd_decap_8
X_160_ _160_/A _164_/A vgnd vpwr scs8hd_buf_1
X_091_ _090_/X _110_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_238 vgnd vpwr scs8hd_fill_1
XANTENNA__152__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_120 vgnd vpwr scs8hd_decap_12
XFILLER_3_219 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_27_175 vpwr vgnd scs8hd_fill_2
X_212_ chany_top_in[4] chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB _129_/Y vgnd vpwr scs8hd_diode_2
X_143_ _123_/A _139_/B _143_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_33_134 vpwr vgnd scs8hd_fill_2
XFILLER_33_123 vpwr vgnd scs8hd_fill_2
XFILLER_33_112 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__147__A _146_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_34 vgnd vpwr scs8hd_decap_12
Xmux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ _180_/Y mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_36 vpwr vgnd scs8hd_fill_2
XFILLER_15_167 vpwr vgnd scs8hd_fill_2
XFILLER_15_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_126_ _125_/Y _167_/B vgnd vpwr scs8hd_buf_1
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[5] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_259 vgnd vpwr scs8hd_decap_12
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
Xmux_right_track_10.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_8_108 vgnd vpwr scs8hd_decap_4
XFILLER_12_104 vgnd vpwr scs8hd_fill_1
XFILLER_16_56 vgnd vpwr scs8hd_decap_6
XFILLER_20_170 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__144__B _139_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_163 vpwr vgnd scs8hd_fill_2
XFILLER_7_174 vpwr vgnd scs8hd_fill_2
X_109_ _109_/A _109_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__160__A _160_/A vgnd vpwr scs8hd_diode_2
XFILLER_34_251 vgnd vpwr scs8hd_decap_12
XFILLER_8_90 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_99 vpwr vgnd scs8hd_fill_2
XFILLER_27_44 vgnd vpwr scs8hd_decap_12
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_37 vpwr vgnd scs8hd_fill_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__155__A _165_/B vgnd vpwr scs8hd_diode_2
XANTENNA__139__B _139_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_1_114 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_13_221 vgnd vpwr scs8hd_fill_1
XFILLER_13_254 vgnd vpwr scs8hd_decap_4
XFILLER_13_265 vpwr vgnd scs8hd_fill_2
XFILLER_9_236 vpwr vgnd scs8hd_fill_2
XFILLER_9_258 vpwr vgnd scs8hd_fill_2
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_184 vgnd vpwr scs8hd_fill_1
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
X_090_ _093_/A address[2] _156_/A _090_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_206 vpwr vgnd scs8hd_fill_2
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_right_track_14.LATCH_0_.latch_SLEEPB _172_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__152__B _149_/B vgnd vpwr scs8hd_diode_2
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XFILLER_36_132 vgnd vpwr scs8hd_decap_12
Xmem_right_track_2.LATCH_0_.latch data_in _174_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_69 vpwr vgnd scs8hd_fill_2
XFILLER_27_143 vpwr vgnd scs8hd_fill_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_27_187 vgnd vpwr scs8hd_decap_12
X_211_ chany_top_in[5] chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
X_142_ _122_/A _139_/B _142_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A bottom_left_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_132 vgnd vpwr scs8hd_decap_4
XANTENNA__163__A _164_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_113 vpwr vgnd scs8hd_fill_2
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_46 vgnd vpwr scs8hd_decap_12
XFILLER_30_149 vgnd vpwr scs8hd_fill_1
XFILLER_30_105 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
X_125_ address[6] _125_/Y vgnd vpwr scs8hd_inv_8
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XFILLER_21_127 vpwr vgnd scs8hd_fill_2
XANTENNA__158__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_20_182 vgnd vpwr scs8hd_decap_3
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _095_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
X_108_ _139_/A _109_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_131 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_12.LATCH_1_.latch_SLEEPB _167_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _222_/A vgnd vpwr scs8hd_inv_1
XFILLER_27_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_12.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _191_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_145 vpwr vgnd scs8hd_fill_2
XFILLER_4_189 vpwr vgnd scs8hd_fill_2
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__171__A _159_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[5] mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__081__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_9_204 vgnd vpwr scs8hd_decap_3
XFILLER_13_200 vpwr vgnd scs8hd_fill_2
XFILLER_0_192 vpwr vgnd scs8hd_fill_2
XANTENNA__166__A _164_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_174 vgnd vpwr scs8hd_decap_8
XANTENNA__076__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_247 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_4_.latch data_in mem_bottom_track_1.LATCH_4_.latch/Q _130_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_144 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_4.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_37 vgnd vpwr scs8hd_decap_8
XFILLER_10_48 vgnd vpwr scs8hd_decap_6
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_27_199 vgnd vpwr scs8hd_decap_12
XFILLER_27_111 vgnd vpwr scs8hd_decap_4
XFILLER_19_57 vgnd vpwr scs8hd_fill_1
X_141_ _110_/A _139_/B _141_/Y vgnd vpwr scs8hd_nor2_4
X_210_ chany_top_in[6] chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_2_265 vgnd vpwr scs8hd_decap_8
XFILLER_2_254 vpwr vgnd scs8hd_fill_2
XFILLER_2_243 vpwr vgnd scs8hd_fill_2
XFILLER_2_221 vgnd vpwr scs8hd_decap_3
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_111 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_33_158 vpwr vgnd scs8hd_fill_2
XFILLER_33_147 vgnd vpwr scs8hd_decap_8
XANTENNA__163__B _164_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd vpwr
+ scs8hd_diode_2
Xmem_right_track_14.LATCH_1_.latch data_in _185_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_71 vpwr vgnd scs8hd_fill_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_58 vgnd vpwr scs8hd_decap_3
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_147 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_10.INVTX1_0_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_124_ _113_/A _118_/X _124_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_91 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_5_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_6 vgnd vpwr scs8hd_decap_12
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_117 vgnd vpwr scs8hd_decap_6
XFILLER_16_69 vpwr vgnd scs8hd_fill_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA__084__A _084_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_11_194 vpwr vgnd scs8hd_fill_2
X_107_ _106_/X _109_/B vgnd vpwr scs8hd_buf_1
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XANTENNA__169__A _160_/A vgnd vpwr scs8hd_diode_2
XANTENNA__079__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_25_275 vpwr vgnd scs8hd_fill_2
XFILLER_25_253 vpwr vgnd scs8hd_fill_2
XFILLER_25_231 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_4_102 vgnd vpwr scs8hd_decap_3
XFILLER_4_113 vpwr vgnd scs8hd_fill_2
XFILLER_4_179 vgnd vpwr scs8hd_fill_1
XFILLER_16_242 vgnd vpwr scs8hd_decap_3
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__171__B _167_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XANTENNA__081__B address[4] vgnd vpwr scs8hd_diode_2
XFILLER_1_138 vpwr vgnd scs8hd_fill_2
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
XANTENNA__166__B _165_/B vgnd vpwr scs8hd_diode_2
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_60 vgnd vpwr scs8hd_fill_1
XFILLER_5_82 vpwr vgnd scs8hd_fill_2
XFILLER_39_142 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vpwr vgnd scs8hd_fill_2
XFILLER_10_226 vpwr vgnd scs8hd_fill_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA__092__A _095_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_18 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_91 vgnd vpwr scs8hd_fill_1
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_10.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_69 vgnd vpwr scs8hd_fill_1
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_123 vgnd vpwr scs8hd_decap_3
XANTENNA__087__A _086_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_140_ _109_/A _139_/B _140_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_145 vgnd vpwr scs8hd_decap_4
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_178 vpwr vgnd scs8hd_fill_2
XANTENNA__163__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_2_50 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_192 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_123_ _123_/A _118_/X _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_118 vgnd vpwr scs8hd_fill_1
XFILLER_12_107 vgnd vpwr scs8hd_fill_1
Xmem_top_track_8.LATCH_3_.latch data_in mem_top_track_8.LATCH_3_.latch/Q _110_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_140 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XFILLER_11_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_144 vpwr vgnd scs8hd_fill_2
XFILLER_11_184 vgnd vpwr scs8hd_fill_1
X_106_ _117_/A _165_/B _163_/C _106_/X vgnd vpwr scs8hd_or3_4
XANTENNA__169__B _165_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XFILLER_25_243 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__095__A _095_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_136 vpwr vgnd scs8hd_fill_2
XFILLER_4_158 vgnd vpwr scs8hd_decap_4
XFILLER_16_232 vgnd vpwr scs8hd_fill_1
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XFILLER_17_80 vpwr vgnd scs8hd_fill_2
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XANTENNA__171__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_22_213 vgnd vpwr scs8hd_fill_1
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XANTENNA__081__C _104_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_13_224 vgnd vpwr scs8hd_fill_1
XFILLER_0_172 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[4] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__166__C _159_/C vgnd vpwr scs8hd_diode_2
XFILLER_39_110 vgnd vpwr scs8hd_decap_12
XFILLER_24_15 vgnd vpwr scs8hd_decap_12
XANTENNA__092__B _110_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_5_.latch data_in mem_bottom_track_9.LATCH_5_.latch/Q _139_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_81 vgnd vpwr scs8hd_decap_4
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _132_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_27_179 vgnd vpwr scs8hd_decap_4
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_201 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_33_116 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_top_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_157 vpwr vgnd scs8hd_fill_2
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__D _163_/D vgnd vpwr scs8hd_diode_2
X_199_ _199_/HI _199_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _192_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_24_138 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_9.LATCH_4_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__A _095_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_182 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_122_ _122_/A _118_/X _122_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_193 vgnd vpwr scs8hd_decap_8
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
Xmem_right_track_10.LATCH_1_.latch data_in _179_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_152 vgnd vpwr scs8hd_fill_1
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XFILLER_7_101 vpwr vgnd scs8hd_fill_2
XFILLER_7_123 vgnd vpwr scs8hd_fill_1
XFILLER_11_163 vgnd vpwr scs8hd_fill_1
X_105_ _105_/A _163_/C vgnd vpwr scs8hd_buf_1
XFILLER_7_167 vpwr vgnd scs8hd_fill_2
XFILLER_7_178 vpwr vgnd scs8hd_fill_2
XFILLER_21_6 vpwr vgnd scs8hd_fill_2
XFILLER_19_263 vpwr vgnd scs8hd_fill_2
XFILLER_19_252 vpwr vgnd scs8hd_fill_2
XFILLER_19_230 vpwr vgnd scs8hd_fill_2
XANTENNA__169__C _170_/C vgnd vpwr scs8hd_diode_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XFILLER_40_247 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__095__B _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_19 vgnd vpwr scs8hd_fill_1
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA__171__D _156_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_39 vgnd vpwr scs8hd_fill_1
XFILLER_1_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_236 vpwr vgnd scs8hd_fill_2
XFILLER_9_218 vpwr vgnd scs8hd_fill_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__166__D _164_/D vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_decap_4
XFILLER_8_273 vpwr vgnd scs8hd_fill_2
XFILLER_5_95 vpwr vgnd scs8hd_fill_2
XFILLER_24_27 vgnd vpwr scs8hd_decap_4
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_206 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_60 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_221 vgnd vpwr scs8hd_decap_4
XFILLER_5_254 vpwr vgnd scs8hd_fill_2
XFILLER_5_265 vpwr vgnd scs8hd_fill_2
XFILLER_14_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_4.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_5_.latch data_in mem_bottom_track_17.LATCH_5_.latch/Q _148_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
Xmux_right_track_6.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_158 vpwr vgnd scs8hd_fill_2
XFILLER_27_103 vpwr vgnd scs8hd_fill_2
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_2_235 vgnd vpwr scs8hd_decap_8
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _187_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/HI _198_/LO vgnd vpwr scs8hd_conb_1
XFILLER_24_117 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_6.LATCH_1_.latch data_in _177_/A _163_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__098__B _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_106 vpwr vgnd scs8hd_fill_2
XFILLER_30_109 vgnd vpwr scs8hd_decap_4
XFILLER_23_161 vpwr vgnd scs8hd_fill_2
X_121_ _110_/A _118_/X _121_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_72 vpwr vgnd scs8hd_fill_2
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XFILLER_22_71 vgnd vpwr scs8hd_fill_1
X_104_ _104_/A address[4] _104_/C _105_/A vgnd vpwr scs8hd_or3_4
XFILLER_11_175 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_275 vpwr vgnd scs8hd_fill_2
XANTENNA__169__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_8_84 vgnd vpwr scs8hd_decap_4
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_8
XFILLER_40_259 vgnd vpwr scs8hd_decap_12
XFILLER_4_149 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_201 vpwr vgnd scs8hd_fill_2
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_71 vpwr vgnd scs8hd_fill_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_22_259 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_204 vpwr vgnd scs8hd_fill_2
XFILLER_0_196 vpwr vgnd scs8hd_fill_2
XFILLER_0_130 vpwr vgnd scs8hd_fill_2
XFILLER_39_189 vpwr vgnd scs8hd_fill_2
XFILLER_39_123 vgnd vpwr scs8hd_decap_12
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_93 vgnd vpwr scs8hd_decap_3
XFILLER_5_200 vpwr vgnd scs8hd_fill_2
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XFILLER_27_115 vgnd vpwr scs8hd_fill_1
XFILLER_19_39 vgnd vpwr scs8hd_decap_3
XFILLER_35_181 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.tap_buf4_0_.scs8hd_inv_1 mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _201_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_258 vgnd vpwr scs8hd_decap_4
XFILLER_18_115 vpwr vgnd scs8hd_fill_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XFILLER_25_93 vpwr vgnd scs8hd_fill_2
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _197_/HI _197_/LO vgnd vpwr scs8hd_conb_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _218_/A vgnd vpwr scs8hd_inv_1
XFILLER_23_140 vpwr vgnd scs8hd_fill_2
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _109_/A _118_/X _120_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_4.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_62 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_18 vgnd vpwr scs8hd_decap_12
XFILLER_20_187 vgnd vpwr scs8hd_decap_3
XFILLER_20_165 vgnd vpwr scs8hd_decap_3
XFILLER_20_110 vgnd vpwr scs8hd_decap_3
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_11_110 vpwr vgnd scs8hd_fill_2
X_103_ address[3] _104_/A vgnd vpwr scs8hd_inv_8
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_198 vpwr vgnd scs8hd_fill_2
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_8_52 vgnd vpwr scs8hd_decap_4
XFILLER_6_191 vpwr vgnd scs8hd_fill_2
XFILLER_27_39 vgnd vpwr scs8hd_decap_3
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_4_117 vpwr vgnd scs8hd_fill_2
XFILLER_16_224 vpwr vgnd scs8hd_fill_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
XFILLER_22_205 vgnd vpwr scs8hd_decap_8
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_12.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vgnd vpwr scs8hd_fill_1
XFILLER_28_93 vgnd vpwr scs8hd_decap_8
XFILLER_5_20 vpwr vgnd scs8hd_fill_2
XFILLER_5_31 vpwr vgnd scs8hd_fill_2
XFILLER_5_42 vpwr vgnd scs8hd_fill_2
XFILLER_5_53 vgnd vpwr scs8hd_decap_4
XFILLER_39_146 vgnd vpwr scs8hd_decap_12
XFILLER_39_135 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _204_/A vgnd vpwr scs8hd_inv_1
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_2_.latch/Q mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__101__A _095_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_4
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_25_72 vgnd vpwr scs8hd_decap_4
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/HI _196_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_6
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_5_ mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_54 vgnd vpwr scs8hd_decap_4
XFILLER_32_163 vgnd vpwr scs8hd_decap_12
XFILLER_17_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_174 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _187_/HI mem_bottom_track_1.LATCH_2_.latch/Q
+ mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_3 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_163 vgnd vpwr scs8hd_decap_8
XFILLER_14_174 vpwr vgnd scs8hd_fill_2
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_2.LATCH_1_.latch data_in _173_/A _157_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_155 vpwr vgnd scs8hd_fill_2
XFILLER_7_148 vgnd vpwr scs8hd_decap_4
X_102_ address[6] _165_/B vgnd vpwr scs8hd_buf_1
Xmux_right_track_2.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_181 vgnd vpwr scs8hd_fill_1
XFILLER_40_239 vgnd vpwr scs8hd_decap_4
XFILLER_4_107 vgnd vpwr scs8hd_decap_3
XFILLER_16_247 vgnd vpwr scs8hd_decap_3
XFILLER_17_84 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_3
XFILLER_3_151 vpwr vgnd scs8hd_fill_2
XANTENNA__104__A _104_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_239 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_217 vgnd vpwr scs8hd_decap_4
XFILLER_28_83 vgnd vpwr scs8hd_fill_1
XFILLER_0_187 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_10 vgnd vpwr scs8hd_decap_6
XFILLER_8_254 vgnd vpwr scs8hd_decap_8
XFILLER_8_265 vgnd vpwr scs8hd_decap_8
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _092_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_0_.latch data_in mem_bottom_track_9.LATCH_0_.latch/Q _144_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_158 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_180 vgnd vpwr scs8hd_decap_3
XANTENNA__101__B _113_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_139 vpwr vgnd scs8hd_fill_2
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_6.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_205 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_9_ mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_128 vpwr vgnd scs8hd_fill_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_172 vpwr vgnd scs8hd_fill_2
XPHY_51 vgnd vpwr scs8hd_decap_3
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/HI _195_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__112__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_131 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_88 vgnd vpwr scs8hd_fill_1
XFILLER_32_175 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _106_/X vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_5_.latch data_in mem_bottom_track_1.LATCH_5_.latch/Q _129_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_127 vpwr vgnd scs8hd_fill_2
X_101_ _095_/A _113_/A _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_134 vgnd vpwr scs8hd_decap_6
XFILLER_22_85 vgnd vpwr scs8hd_fill_1
XFILLER_22_74 vpwr vgnd scs8hd_fill_2
XFILLER_22_63 vpwr vgnd scs8hd_fill_2
XFILLER_19_234 vpwr vgnd scs8hd_fill_2
XFILLER_19_201 vgnd vpwr scs8hd_fill_1
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_19_267 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_259 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__210__A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_16_259 vgnd vpwr scs8hd_decap_12
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_95 vpwr vgnd scs8hd_fill_2
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_3_130 vpwr vgnd scs8hd_fill_2
XANTENNA__104__B address[4] vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _153_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_6.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_240 vgnd vpwr scs8hd_decap_4
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
XFILLER_28_40 vpwr vgnd scs8hd_fill_2
XFILLER_8_211 vgnd vpwr scs8hd_decap_3
XANTENNA__115__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_8_244 vgnd vpwr scs8hd_fill_1
XFILLER_12_273 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_66 vgnd vpwr scs8hd_fill_1
XFILLER_5_99 vgnd vpwr scs8hd_decap_4
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_0_.latch data_in mem_bottom_track_17.LATCH_0_.latch/Q _153_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_236 vgnd vpwr scs8hd_decap_6
XFILLER_5_258 vgnd vpwr scs8hd_decap_4
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XFILLER_14_97 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_4_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_27_107 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_3_ vgnd vpwr scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_162 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_10.INVTX1_1_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr
+ scs8hd_diode_2
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_41 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/HI _194_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_67 vpwr vgnd scs8hd_fill_2
XFILLER_2_23 vgnd vpwr scs8hd_decap_8
XFILLER_2_12 vgnd vpwr scs8hd_decap_8
XANTENNA__112__B _109_/B vgnd vpwr scs8hd_diode_2
XFILLER_17_140 vgnd vpwr scs8hd_fill_1
XFILLER_17_173 vgnd vpwr scs8hd_decap_4
XFILLER_32_187 vgnd vpwr scs8hd_decap_12
XFILLER_23_198 vgnd vpwr scs8hd_decap_12
XFILLER_23_187 vgnd vpwr scs8hd_decap_3
XANTENNA__213__A _213_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_10 vgnd vpwr scs8hd_decap_12
XFILLER_11_87 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__A _123_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__208__A right_top_grid_pin_10_ vgnd vpwr scs8hd_diode_2
X_100_ _099_/X _113_/A vgnd vpwr scs8hd_buf_1
XFILLER_19_213 vpwr vgnd scs8hd_fill_2
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _118_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_16_205 vpwr vgnd scs8hd_fill_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_53 vpwr vgnd scs8hd_fill_2
XFILLER_17_75 vgnd vpwr scs8hd_decap_3
XFILLER_17_97 vpwr vgnd scs8hd_fill_2
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_175 vpwr vgnd scs8hd_fill_2
XFILLER_3_164 vpwr vgnd scs8hd_fill_2
XANTENNA__104__C _104_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA__120__B _118_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_6.INVTX1_1_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_21_263 vgnd vpwr scs8hd_decap_12
XANTENNA__221__A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_3
XFILLER_0_123 vgnd vpwr scs8hd_fill_1
XFILLER_0_134 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_63 vgnd vpwr scs8hd_fill_1
XFILLER_8_201 vpwr vgnd scs8hd_fill_2
Xmem_top_track_8.LATCH_4_.latch data_in mem_top_track_8.LATCH_4_.latch/Q _109_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_78 vpwr vgnd scs8hd_fill_2
XANTENNA__115__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA__131__A _110_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vgnd vpwr scs8hd_decap_8
XFILLER_14_43 vgnd vpwr scs8hd_decap_8
XFILLER_14_87 vpwr vgnd scs8hd_fill_2
XANTENNA__216__A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_5_204 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_36_108 vgnd vpwr scs8hd_decap_12
XANTENNA__126__A _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XFILLER_35_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vpwr vgnd scs8hd_fill_2
XPHY_42 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
X_193_ _193_/HI _193_/LO vgnd vpwr scs8hd_conb_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_199 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_144 vpwr vgnd scs8hd_fill_2
XFILLER_11_22 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_3_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_96 vgnd vpwr scs8hd_decap_12
XFILLER_14_122 vgnd vpwr scs8hd_fill_1
XFILLER_14_133 vgnd vpwr scs8hd_fill_1
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__B _118_/X vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XFILLER_20_136 vpwr vgnd scs8hd_fill_2
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XANTENNA__224__A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
X_159_ _159_/A _164_/B _159_/C _164_/D _159_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_195 vpwr vgnd scs8hd_fill_2
XANTENNA__134__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_228 vgnd vpwr scs8hd_decap_4
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__219__A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_6
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_198 vpwr vgnd scs8hd_fill_2
XANTENNA__129__A _139_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_275 vpwr vgnd scs8hd_fill_2
XFILLER_0_168 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_86 vgnd vpwr scs8hd_decap_6
XFILLER_28_75 vpwr vgnd scs8hd_fill_2
XANTENNA__131__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_24 vpwr vgnd scs8hd_fill_2
XFILLER_5_35 vpwr vgnd scs8hd_fill_2
XFILLER_5_46 vpwr vgnd scs8hd_fill_2
XFILLER_5_57 vgnd vpwr scs8hd_fill_1
XANTENNA__115__C _104_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_77 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XFILLER_29_172 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_2.LATCH_1_.latch_SLEEPB _157_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _122_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_120 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_bottom_track_9.LATCH_5_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_3_ mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_65 vgnd vpwr scs8hd_decap_4
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/HI _192_/LO vgnd vpwr scs8hd_conb_1
XFILLER_1_230 vpwr vgnd scs8hd_fill_2
Xmux_right_track_14.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_145 vgnd vpwr scs8hd_decap_8
XFILLER_32_123 vgnd vpwr scs8hd_decap_8
XANTENNA__137__A _117_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_197 vpwr vgnd scs8hd_fill_2
XFILLER_23_178 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_34 vgnd vpwr scs8hd_decap_8
XFILLER_14_101 vpwr vgnd scs8hd_fill_2
XFILLER_14_145 vgnd vpwr scs8hd_decap_6
XFILLER_14_178 vgnd vpwr scs8hd_decap_6
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XFILLER_20_115 vpwr vgnd scs8hd_fill_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XFILLER_28_204 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_4.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_104 vgnd vpwr scs8hd_decap_4
XFILLER_22_88 vpwr vgnd scs8hd_fill_2
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XFILLER_11_159 vgnd vpwr scs8hd_decap_4
Xmux_right_track_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ _178_/A mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_19_259 vpwr vgnd scs8hd_fill_2
XFILLER_19_248 vpwr vgnd scs8hd_fill_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_35 vpwr vgnd scs8hd_fill_2
XFILLER_8_79 vpwr vgnd scs8hd_fill_2
X_158_ address[0] _164_/D vgnd vpwr scs8hd_buf_1
X_089_ address[1] _093_/A vgnd vpwr scs8hd_inv_8
XFILLER_10_181 vpwr vgnd scs8hd_fill_2
XANTENNA__134__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA__150__A _110_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_207 vgnd vpwr scs8hd_decap_12
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_43 vgnd vpwr scs8hd_decap_12
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_251 vgnd vpwr scs8hd_decap_12
XANTENNA__129__B _134_/B vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_21_221 vpwr vgnd scs8hd_fill_2
XFILLER_21_210 vpwr vgnd scs8hd_fill_2
XFILLER_0_103 vpwr vgnd scs8hd_fill_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_8
XFILLER_0_147 vpwr vgnd scs8hd_fill_2
XFILLER_0_125 vgnd vpwr scs8hd_fill_1
XFILLER_12_210 vpwr vgnd scs8hd_fill_2
XFILLER_8_236 vgnd vpwr scs8hd_decap_8
XFILLER_12_243 vpwr vgnd scs8hd_fill_2
XFILLER_12_254 vpwr vgnd scs8hd_fill_2
XFILLER_12_265 vgnd vpwr scs8hd_decap_8
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_217 vpwr vgnd scs8hd_fill_2
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_39_86 vgnd vpwr scs8hd_decap_12
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XFILLER_29_151 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__142__B _139_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _197_/HI mem_top_track_0.LATCH_2_.latch/Q
+ mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_209 vgnd vpwr scs8hd_decap_3
XFILLER_26_110 vpwr vgnd scs8hd_fill_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_176 vgnd vpwr scs8hd_decap_4
XFILLER_26_154 vpwr vgnd scs8hd_fill_2
XFILLER_26_143 vgnd vpwr scs8hd_decap_4
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ _191_/HI _191_/LO vgnd vpwr scs8hd_conb_1
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XFILLER_17_165 vpwr vgnd scs8hd_fill_2
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__137__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA__153__A _113_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_157 vpwr vgnd scs8hd_fill_2
XFILLER_23_113 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XFILLER_11_68 vpwr vgnd scs8hd_fill_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_0_.latch data_in mem_bottom_track_1.LATCH_0_.latch/Q _134_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__148__A _139_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_12.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_12.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_36_271 vgnd vpwr scs8hd_decap_4
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_22_67 vgnd vpwr scs8hd_decap_4
XFILLER_22_56 vgnd vpwr scs8hd_decap_4
XFILLER_19_238 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_226_ _226_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
X_157_ _159_/A _164_/B _159_/C _163_/D _157_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_8_58 vpwr vgnd scs8hd_fill_2
XFILLER_8_69 vgnd vpwr scs8hd_decap_4
XFILLER_10_193 vpwr vgnd scs8hd_fill_2
XANTENNA__150__B _149_/B vgnd vpwr scs8hd_diode_2
X_088_ _095_/A _109_/A _088_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_219 vgnd vpwr scs8hd_decap_12
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_263 vgnd vpwr scs8hd_decap_12
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_99 vpwr vgnd scs8hd_fill_2
XFILLER_33_55 vgnd vpwr scs8hd_decap_6
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_134 vpwr vgnd scs8hd_fill_2
XFILLER_3_123 vgnd vpwr scs8hd_decap_3
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_211 vgnd vpwr scs8hd_decap_3
XANTENNA__161__A _164_/A vgnd vpwr scs8hd_diode_2
X_209_ _209_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_200 vpwr vgnd scs8hd_fill_2
XFILLER_12_222 vpwr vgnd scs8hd_fill_2
XFILLER_8_215 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_10.tap_buf4_0_.scs8hd_inv_1 mux_right_track_10.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vpwr scs8hd_inv_1
XANTENNA__156__A _156_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_270 vpwr vgnd scs8hd_fill_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_39_10 vgnd vpwr scs8hd_decap_12
XFILLER_39_98 vgnd vpwr scs8hd_decap_12
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 top_left_grid_pin_7_ mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_100 vgnd vpwr scs8hd_decap_12
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_25_89 vpwr vgnd scs8hd_fill_2
X_190_ _190_/HI _190_/LO vgnd vpwr scs8hd_conb_1
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_2_38 vgnd vpwr scs8hd_fill_1
XFILLER_1_265 vpwr vgnd scs8hd_fill_2
XFILLER_1_254 vpwr vgnd scs8hd_fill_2
XANTENNA__137__C _159_/C vgnd vpwr scs8hd_diode_2
XANTENNA__153__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
XFILLER_14_125 vpwr vgnd scs8hd_fill_2
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
XFILLER_20_106 vpwr vgnd scs8hd_fill_2
XANTENNA__148__B _149_/B vgnd vpwr scs8hd_diode_2
XANTENNA__164__A _164_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _130_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_151 vpwr vgnd scs8hd_fill_2
XFILLER_9_162 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_3
XFILLER_3_81 vpwr vgnd scs8hd_fill_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_22_79 vgnd vpwr scs8hd_decap_6
XFILLER_19_217 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_11_ mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_087_ _086_/X _109_/A vgnd vpwr scs8hd_buf_1
XFILLER_6_132 vpwr vgnd scs8hd_fill_2
XFILLER_6_165 vpwr vgnd scs8hd_fill_2
X_156_ _156_/A _163_/D vgnd vpwr scs8hd_buf_1
X_225_ chany_bottom_in[0] chany_top_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _159_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_10.INVTX1_1_.scs8hd_inv_1 chany_bottom_in[2] mux_right_track_10.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_209 vgnd vpwr scs8hd_decap_3
XFILLER_17_57 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_102 vpwr vgnd scs8hd_fill_2
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_168 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__161__B _164_/B vgnd vpwr scs8hd_diode_2
X_208_ right_top_grid_pin_10_ chanx_right_out[0] vgnd vpwr scs8hd_buf_2
X_139_ _139_/A _139_/B _139_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_4.tap_buf4_0_.scs8hd_inv_1 mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A
+ _206_/A vgnd vpwr scs8hd_inv_1
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_201 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_10.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_0_116 vgnd vpwr scs8hd_decap_4
XFILLER_28_45 vgnd vpwr scs8hd_decap_12
XFILLER_8_205 vgnd vpwr scs8hd_decap_4
XFILLER_5_16 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__A _159_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A _081_/X vgnd vpwr scs8hd_diode_2
XFILLER_39_22 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_4_230 vpwr vgnd scs8hd_fill_2
XFILLER_4_252 vpwr vgnd scs8hd_fill_2
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_35_112 vgnd vpwr scs8hd_decap_8
XFILLER_35_145 vgnd vpwr scs8hd_decap_12
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A _159_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_189 vgnd vpwr scs8hd_decap_12
XPHY_46 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A address[1] vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vpwr vgnd scs8hd_fill_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_101 vpwr vgnd scs8hd_fill_2
XFILLER_17_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_31_170 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _088_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _183_/A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_9.LATCH_1_.latch data_in mem_bottom_track_9.LATCH_1_.latch/Q _143_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_172_ _159_/A _167_/B _163_/C address[0] _172_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _193_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__164__B _164_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_130 vpwr vgnd scs8hd_fill_2
XFILLER_13_170 vgnd vpwr scs8hd_fill_1
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_196 vpwr vgnd scs8hd_fill_2
XFILLER_3_60 vgnd vpwr scs8hd_fill_1
XFILLER_36_251 vgnd vpwr scs8hd_decap_4
Xmux_right_track_6.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[5] mux_right_track_6.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
XANTENNA__090__A _093_/A vgnd vpwr scs8hd_diode_2
X_224_ chany_bottom_in[1] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_155_ _165_/B _164_/B vgnd vpwr scs8hd_buf_1
X_086_ address[1] _086_/B address[0] _086_/X vgnd vpwr scs8hd_or3_4
XFILLER_6_177 vpwr vgnd scs8hd_fill_2
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _164_/B vgnd vpwr scs8hd_diode_2
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_47 vgnd vpwr scs8hd_fill_1
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XANTENNA__085__A _139_/A vgnd vpwr scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_114 vpwr vgnd scs8hd_fill_2
XFILLER_3_147 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_210 vpwr vgnd scs8hd_fill_2
X_207_ _207_/A chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_15_254 vpwr vgnd scs8hd_fill_2
XFILLER_15_265 vpwr vgnd scs8hd_fill_2
XANTENNA__161__C _161_/C vgnd vpwr scs8hd_diode_2
X_138_ _137_/X _139_/B vgnd vpwr scs8hd_buf_1
XFILLER_24_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ _176_/A mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_0_72 vpwr vgnd scs8hd_fill_2
XFILLER_0_94 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_92 vpwr vgnd scs8hd_fill_2
XFILLER_28_79 vgnd vpwr scs8hd_decap_4
XFILLER_28_57 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_12.LATCH_0_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_12.LATCH_0_.latch data_in _182_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__172__B _167_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_34 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 chanx_right_in[2] mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_135 vgnd vpwr scs8hd_decap_3
XFILLER_35_157 vgnd vpwr scs8hd_decap_12
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
XANTENNA__167__B _167_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_71 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_26_135 vpwr vgnd scs8hd_fill_2
XFILLER_25_69 vgnd vpwr scs8hd_fill_1
XFILLER_25_47 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _086_/B vgnd vpwr scs8hd_diode_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA__093__A _093_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_234 vgnd vpwr scs8hd_decap_4
XFILLER_1_212 vgnd vpwr scs8hd_fill_1
XFILLER_17_179 vpwr vgnd scs8hd_fill_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_182 vgnd vpwr scs8hd_fill_1
XANTENNA__088__A _095_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_105 vgnd vpwr scs8hd_decap_4
X_171_ _159_/A _167_/B _163_/C _156_/A _171_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_10.LATCH_1_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_17.LATCH_1_.latch data_in mem_bottom_track_17.LATCH_1_.latch/Q _152_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__164__C _163_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_175 vpwr vgnd scs8hd_fill_2
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_6.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__090__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_263 vgnd vpwr scs8hd_decap_12
Xmux_right_track_12.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_12.INVTX1_2_.scs8hd_inv_1/Y
+ _182_/A mux_right_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
X_223_ chany_bottom_in[2] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_8_39 vpwr vgnd scs8hd_fill_2
XFILLER_6_112 vgnd vpwr scs8hd_fill_1
XFILLER_6_145 vgnd vpwr scs8hd_decap_8
XFILLER_10_163 vgnd vpwr scs8hd_decap_3
XFILLER_10_185 vpwr vgnd scs8hd_fill_2
X_085_ _139_/A _095_/A _085_/Y vgnd vpwr scs8hd_nor2_4
X_154_ _117_/A _159_/A vgnd vpwr scs8hd_buf_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__159__C _159_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_241 vgnd vpwr scs8hd_decap_8
XFILLER_18_252 vgnd vpwr scs8hd_decap_8
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__085__B _095_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_4.INVTX1_2_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_4.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_right_track_8.LATCH_0_.latch data_in _184_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_206_ _206_/A chanx_right_out[2] vgnd vpwr scs8hd_buf_2
X_137_ _117_/A _167_/B _159_/C _137_/X vgnd vpwr scs8hd_or3_4
XANTENNA__161__D _163_/D vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
XFILLER_21_225 vgnd vpwr scs8hd_decap_8
XFILLER_21_214 vgnd vpwr scs8hd_decap_4
XFILLER_9_71 vpwr vgnd scs8hd_fill_2
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_4.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__096__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_258 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_7_240 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__172__C _163_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_9_ vgnd vpwr scs8hd_diode_2
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_39_46 vgnd vpwr scs8hd_decap_12
XFILLER_29_155 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr
+ scs8hd_diode_2
XFILLER_4_210 vgnd vpwr scs8hd_decap_4
XFILLER_4_243 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_169 vgnd vpwr scs8hd_decap_12
XANTENNA__167__C _161_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_50 vpwr vgnd scs8hd_fill_2
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_26_158 vgnd vpwr scs8hd_decap_4
XFILLER_26_114 vpwr vgnd scs8hd_fill_2
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XPHY_48 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__077__C _156_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_136 vpwr vgnd scs8hd_fill_2
XFILLER_17_169 vpwr vgnd scs8hd_fill_2
XFILLER_32_106 vgnd vpwr scs8hd_decap_8
XFILLER_25_191 vpwr vgnd scs8hd_fill_2
XFILLER_15_81 vpwr vgnd scs8hd_fill_2
XFILLER_23_117 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_5_.latch data_in mem_top_track_8.LATCH_5_.latch/Q _108_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A bottom_left_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__088__B _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_194 vgnd vpwr scs8hd_decap_8
XFILLER_22_150 vgnd vpwr scs8hd_decap_3
X_170_ _160_/A _165_/B _170_/C _164_/D _170_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA__164__D _164_/D vgnd vpwr scs8hd_diode_2
XFILLER_3_40 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_4
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA__090__C _156_/A vgnd vpwr scs8hd_diode_2
XANTENNA__099__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_27_275 vpwr vgnd scs8hd_fill_2
XFILLER_27_253 vpwr vgnd scs8hd_fill_2
X_222_ _222_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_6_102 vpwr vgnd scs8hd_fill_2
X_153_ _113_/A _149_/B _153_/Y vgnd vpwr scs8hd_nor2_4
X_084_ _084_/A _095_/A vgnd vpwr scs8hd_buf_1
XFILLER_12_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA__159__D _164_/D vgnd vpwr scs8hd_diode_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_6.INVTX1_2_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _139_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_205_ _205_/A chanx_right_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_23_92 vpwr vgnd scs8hd_fill_2
XFILLER_23_81 vpwr vgnd scs8hd_fill_2
X_136_ _136_/A _159_/C vgnd vpwr scs8hd_buf_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_182 vgnd vpwr scs8hd_decap_4
XFILLER_0_63 vpwr vgnd scs8hd_fill_2
XFILLER_0_85 vpwr vgnd scs8hd_fill_2
XFILLER_21_259 vpwr vgnd scs8hd_fill_2
XFILLER_21_248 vgnd vpwr scs8hd_decap_6
XFILLER_21_204 vgnd vpwr scs8hd_decap_3
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XANTENNA__096__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_12_204 vgnd vpwr scs8hd_decap_4
XFILLER_20_270 vgnd vpwr scs8hd_decap_4
XFILLER_8_219 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _197_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_237 vgnd vpwr scs8hd_decap_4
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_12.INVTX1_0_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_7_274 vgnd vpwr scs8hd_decap_3
XANTENNA__172__D address[0] vgnd vpwr scs8hd_diode_2
X_119_ _139_/A _118_/X _119_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_2.INVTX1_2_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_58 vgnd vpwr scs8hd_decap_3
XFILLER_29_134 vpwr vgnd scs8hd_fill_2
XFILLER_29_123 vgnd vpwr scs8hd_decap_6
XFILLER_29_101 vpwr vgnd scs8hd_fill_2
XANTENNA__167__D _163_/D vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA__093__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
XFILLER_1_258 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_170 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XFILLER_14_118 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XFILLER_14_129 vgnd vpwr scs8hd_decap_4
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_13_151 vpwr vgnd scs8hd_fill_2
XFILLER_13_173 vgnd vpwr scs8hd_decap_4
XFILLER_13_184 vgnd vpwr scs8hd_decap_3
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_85 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__099__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_27_243 vgnd vpwr scs8hd_fill_1
X_221_ chany_bottom_in[4] chany_top_out[5] vgnd vpwr scs8hd_buf_2
X_083_ _117_/A address[6] _161_/C _084_/A vgnd vpwr scs8hd_or3_4
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_152_ _123_/A _149_/B _152_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_6_169 vgnd vpwr scs8hd_decap_8
Xmux_right_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _177_/A mux_right_track_6.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_213 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_39 vgnd vpwr scs8hd_decap_8
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XFILLER_3_106 vpwr vgnd scs8hd_fill_2
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
X_204_ _204_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_15_235 vpwr vgnd scs8hd_fill_2
X_135_ _104_/A _115_/B _104_/C _136_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XANTENNA__096__C _156_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_82 vgnd vpwr scs8hd_decap_4
XFILLER_18_93 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
X_118_ _118_/A _118_/X vgnd vpwr scs8hd_buf_1
Xmem_right_track_4.LATCH_0_.latch data_in _176_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_168 vpwr vgnd scs8hd_fill_2
Xmux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ _174_/A mux_right_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_70 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_26_149 vgnd vpwr scs8hd_decap_4
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_39 vgnd vpwr scs8hd_decap_8
XPHY_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XFILLER_1_215 vpwr vgnd scs8hd_fill_2
XFILLER_25_182 vgnd vpwr scs8hd_fill_1
XFILLER_17_149 vgnd vpwr scs8hd_decap_3
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_31_174 vgnd vpwr scs8hd_decap_8
XFILLER_31_163 vgnd vpwr scs8hd_decap_4
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
Xmux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _185_/A mux_right_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
XFILLER_22_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _195_/HI _178_/Y mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_123 vgnd vpwr scs8hd_decap_4
XFILLER_9_134 vpwr vgnd scs8hd_fill_2
XFILLER_13_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_53 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _194_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_211 vgnd vpwr scs8hd_decap_12
XANTENNA__099__C address[0] vgnd vpwr scs8hd_diode_2
X_220_ chany_bottom_in[5] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_115 vgnd vpwr scs8hd_decap_4
X_151_ _122_/A _149_/B _151_/Y vgnd vpwr scs8hd_nor2_4
X_082_ _081_/X _161_/C vgnd vpwr scs8hd_buf_1
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[0] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _198_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_33_39 vpwr vgnd scs8hd_fill_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_118 vpwr vgnd scs8hd_fill_2
XFILLER_15_214 vpwr vgnd scs8hd_fill_2
X_203_ _203_/A chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_258 vgnd vpwr scs8hd_decap_4
XFILLER_15_269 vgnd vpwr scs8hd_decap_8
XFILLER_2_140 vgnd vpwr scs8hd_fill_1
X_134_ _113_/A _134_/B _134_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ _180_/A mux_right_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_2_173 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_1.LATCH_1_.latch data_in mem_bottom_track_1.LATCH_1_.latch/Q _133_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_32 vpwr vgnd scs8hd_fill_2
XFILLER_0_43 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_6
XFILLER_7_221 vpwr vgnd scs8hd_fill_2
XFILLER_11_261 vpwr vgnd scs8hd_fill_2
X_117_ _117_/A address[6] _170_/C _118_/A vgnd vpwr scs8hd_or3_4
XFILLER_15_3 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _184_/A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_84 vpwr vgnd scs8hd_fill_2
XFILLER_28_180 vgnd vpwr scs8hd_decap_12
XFILLER_26_139 vpwr vgnd scs8hd_fill_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XANTENNA__102__A address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_142 vpwr vgnd scs8hd_fill_2
XFILLER_39_275 vpwr vgnd scs8hd_fill_2
XFILLER_39_231 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_6.LATCH_1_.latch_SLEEPB _163_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_98 vpwr vgnd scs8hd_fill_2
XFILLER_8_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_8
XFILLER_27_223 vgnd vpwr scs8hd_decap_12
X_150_ _110_/A _149_/B _150_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_081_ address[3] address[4] _104_/C _081_/X vgnd vpwr scs8hd_or3_4
XFILLER_10_145 vgnd vpwr scs8hd_decap_8
XFILLER_10_189 vpwr vgnd scs8hd_fill_2
XFILLER_12_63 vpwr vgnd scs8hd_fill_2
XFILLER_12_96 vpwr vgnd scs8hd_fill_2
XFILLER_5_171 vgnd vpwr scs8hd_decap_8
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A top_left_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd vpwr
+ scs8hd_diode_2
X_202_ _202_/A chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_23_73 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vpwr vgnd scs8hd_fill_2
XFILLER_23_51 vgnd vpwr scs8hd_decap_3
X_133_ _123_/A _134_/B _133_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_2_163 vpwr vgnd scs8hd_fill_2
XANTENNA__110__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_99 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_42 vgnd vpwr scs8hd_decap_3
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
XFILLER_9_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_218 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_10.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_10.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_116_ _115_/X _170_/C vgnd vpwr scs8hd_buf_1
XFILLER_7_200 vgnd vpwr scs8hd_decap_3
XFILLER_7_255 vpwr vgnd scs8hd_fill_2
XFILLER_7_266 vpwr vgnd scs8hd_fill_2
XANTENNA__105__A _105_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_240 vpwr vgnd scs8hd_fill_2
XFILLER_4_203 vgnd vpwr scs8hd_decap_4
XFILLER_4_247 vgnd vpwr scs8hd_decap_3
XFILLER_28_192 vgnd vpwr scs8hd_decap_12
XFILLER_6_32 vgnd vpwr scs8hd_decap_6
XFILLER_6_54 vpwr vgnd scs8hd_fill_2
XFILLER_34_151 vpwr vgnd scs8hd_fill_2
XPHY_19 vgnd vpwr scs8hd_decap_3
Xmem_top_track_8.LATCH_0_.latch data_in mem_top_track_8.LATCH_0_.latch/Q _113_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_195 vgnd vpwr scs8hd_decap_12
XFILLER_25_140 vpwr vgnd scs8hd_fill_2
XFILLER_15_85 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
XFILLER_0_261 vpwr vgnd scs8hd_fill_2
XFILLER_16_184 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_22_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vpwr vgnd scs8hd_fill_2
XFILLER_26_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_147 vpwr vgnd scs8hd_fill_2
XFILLER_9_158 vpwr vgnd scs8hd_fill_2
XFILLER_13_143 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A _113_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_235 vgnd vpwr scs8hd_decap_8
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
X_080_ enable _104_/C vgnd vpwr scs8hd_inv_8
XFILLER_6_106 vgnd vpwr scs8hd_decap_6
XFILLER_10_124 vpwr vgnd scs8hd_fill_2
XFILLER_10_168 vpwr vgnd scs8hd_fill_2
XFILLER_6_128 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 bottom_left_grid_pin_15_ mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_202 vpwr vgnd scs8hd_fill_2
XFILLER_18_224 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _139_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
XFILLER_24_205 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_12.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_12.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_271 vgnd vpwr scs8hd_decap_4
X_201_ _201_/A chanx_right_out[7] vgnd vpwr scs8hd_buf_2
X_132_ _122_/A _134_/B _132_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _085_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_2_197 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_2_.latch data_in mem_bottom_track_9.LATCH_2_.latch/Q _142_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__110__B _109_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_12 vpwr vgnd scs8hd_fill_2
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
Xmux_right_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _175_/A mux_right_track_4.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_274 vgnd vpwr scs8hd_fill_1
XANTENNA__211__A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_52 vpwr vgnd scs8hd_fill_2
XFILLER_18_63 vpwr vgnd scs8hd_fill_2
XFILLER_34_40 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
X_115_ address[3] _115_/B _104_/C _115_/X vgnd vpwr scs8hd_or3_4
XFILLER_7_245 vgnd vpwr scs8hd_fill_1
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA__121__A _110_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_138 vpwr vgnd scs8hd_fill_2
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_215 vpwr vgnd scs8hd_fill_2
XFILLER_4_226 vpwr vgnd scs8hd_fill_2
XFILLER_29_62 vgnd vpwr scs8hd_fill_1
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA__116__A _115_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_130 vgnd vpwr scs8hd_decap_8
XFILLER_19_193 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _196_/HI _183_/Y mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_174 vgnd vpwr scs8hd_decap_6
XFILLER_15_31 vgnd vpwr scs8hd_decap_12
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _189_/HI vgnd vpwr
+ scs8hd_diode_2
.ends

