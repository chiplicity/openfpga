VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_3__1_
  CLASS BLOCK ;
  FOREIGN cby_3__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 110.000 BY 110.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 4.120 110.000 4.720 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 12.960 110.000 13.560 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 22.480 110.000 23.080 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 31.320 110.000 31.920 ;
    END
  END address[6]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 107.600 4.510 110.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 107.600 13.250 110.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 40.840 110.000 41.440 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.170 107.600 22.450 110.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 107.600 31.650 110.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.400 13.560 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.570 107.600 40.850 110.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 2.400 23.080 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 49.680 110.000 50.280 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 59.200 110.000 59.800 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 49.770 107.600 50.050 110.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 107.600 59.250 110.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 107.600 68.450 110.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 2.400 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.400 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 2.400 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 107.600 77.650 110.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 2.400 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.400 41.440 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 107.600 68.040 110.000 68.640 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 2.400 50.280 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 2.400 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 77.560 110.000 78.160 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 86.400 110.000 87.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 2.400 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 2.400 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 95.920 110.000 96.520 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END enable
  PIN left_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 2.400 ;
    END
  END left_grid_pin_1_
  PIN left_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 86.570 107.600 86.850 110.000 ;
    END
  END left_grid_pin_5_
  PIN left_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 107.600 96.050 110.000 ;
    END
  END left_grid_pin_9_
  PIN right_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 2.400 78.160 ;
    END
  END right_grid_pin_0_
  PIN right_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END right_grid_pin_10_
  PIN right_grid_pin_12_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.970 107.600 105.250 110.000 ;
    END
  END right_grid_pin_12_
  PIN right_grid_pin_14_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 2.400 105.360 ;
    END
  END right_grid_pin_14_
  PIN right_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 2.400 87.000 ;
    END
  END right_grid_pin_2_
  PIN right_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 2.400 ;
    END
  END right_grid_pin_4_
  PIN right_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 2.400 96.520 ;
    END
  END right_grid_pin_6_
  PIN right_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 107.600 104.760 110.000 105.360 ;
    END
  END right_grid_pin_8_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 23.055 10.640 24.655 98.160 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 41.385 10.640 42.985 98.160 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 104.420 98.005 ;
      LAYER met1 ;
        RECT 0.530 0.040 108.030 107.740 ;
      LAYER met2 ;
        RECT 0.550 107.320 3.950 107.850 ;
        RECT 4.790 107.320 12.690 107.850 ;
        RECT 13.530 107.320 21.890 107.850 ;
        RECT 22.730 107.320 31.090 107.850 ;
        RECT 31.930 107.320 40.290 107.850 ;
        RECT 41.130 107.320 49.490 107.850 ;
        RECT 50.330 107.320 58.690 107.850 ;
        RECT 59.530 107.320 67.890 107.850 ;
        RECT 68.730 107.320 77.090 107.850 ;
        RECT 77.930 107.320 86.290 107.850 ;
        RECT 87.130 107.320 95.490 107.850 ;
        RECT 96.330 107.320 104.690 107.850 ;
        RECT 105.530 107.320 108.010 107.850 ;
        RECT 0.550 2.680 108.010 107.320 ;
        RECT 0.550 0.270 2.110 2.680 ;
        RECT 2.950 0.270 7.170 2.680 ;
        RECT 8.010 0.270 12.690 2.680 ;
        RECT 13.530 0.270 18.210 2.680 ;
        RECT 19.050 0.270 23.730 2.680 ;
        RECT 24.570 0.270 29.250 2.680 ;
        RECT 30.090 0.270 34.770 2.680 ;
        RECT 35.610 0.270 40.290 2.680 ;
        RECT 41.130 0.270 45.810 2.680 ;
        RECT 46.650 0.270 51.330 2.680 ;
        RECT 52.170 0.270 56.850 2.680 ;
        RECT 57.690 0.270 62.370 2.680 ;
        RECT 63.210 0.270 67.890 2.680 ;
        RECT 68.730 0.270 73.410 2.680 ;
        RECT 74.250 0.270 78.930 2.680 ;
        RECT 79.770 0.270 84.450 2.680 ;
        RECT 85.290 0.270 89.970 2.680 ;
        RECT 90.810 0.270 95.490 2.680 ;
        RECT 96.330 0.270 101.010 2.680 ;
        RECT 101.850 0.270 106.530 2.680 ;
        RECT 107.370 0.270 108.010 2.680 ;
      LAYER met3 ;
        RECT 2.800 104.360 107.200 104.760 ;
        RECT 0.270 96.920 108.290 104.360 ;
        RECT 2.800 95.520 107.200 96.920 ;
        RECT 0.270 87.400 108.290 95.520 ;
        RECT 2.800 86.000 107.200 87.400 ;
        RECT 0.270 78.560 108.290 86.000 ;
        RECT 2.800 77.160 107.200 78.560 ;
        RECT 0.270 69.040 108.290 77.160 ;
        RECT 2.800 67.640 107.200 69.040 ;
        RECT 0.270 60.200 108.290 67.640 ;
        RECT 2.800 58.800 107.200 60.200 ;
        RECT 0.270 50.680 108.290 58.800 ;
        RECT 2.800 49.280 107.200 50.680 ;
        RECT 0.270 41.840 108.290 49.280 ;
        RECT 2.800 40.440 107.200 41.840 ;
        RECT 0.270 32.320 108.290 40.440 ;
        RECT 2.800 30.920 107.200 32.320 ;
        RECT 0.270 23.480 108.290 30.920 ;
        RECT 2.800 22.080 107.200 23.480 ;
        RECT 0.270 13.960 108.290 22.080 ;
        RECT 2.800 12.560 107.200 13.960 ;
        RECT 0.270 5.120 108.290 12.560 ;
        RECT 2.800 4.720 107.200 5.120 ;
      LAYER met4 ;
        RECT 0.295 10.240 22.655 98.160 ;
        RECT 25.055 10.240 40.985 98.160 ;
        RECT 43.385 10.240 108.265 98.160 ;
        RECT 0.295 6.975 108.265 10.240 ;
  END
END cby_3__1_
END LIBRARY

