magic
tech sky130A
magscale 1 2
timestamp 1609025059
<< locali >>
rect 6653 9367 6687 9469
rect 2605 3451 2639 3689
<< viali >>
rect 5089 17289 5123 17323
rect 5917 17289 5951 17323
rect 6377 17289 6411 17323
rect 7113 17289 7147 17323
rect 7481 17289 7515 17323
rect 7757 17289 7791 17323
rect 8217 17289 8251 17323
rect 8677 17289 8711 17323
rect 9413 17289 9447 17323
rect 2697 17221 2731 17255
rect 10885 17221 10919 17255
rect 1685 17153 1719 17187
rect 2237 17153 2271 17187
rect 4813 17153 4847 17187
rect 9781 17153 9815 17187
rect 1501 17085 1535 17119
rect 2053 17085 2087 17119
rect 2789 17085 2823 17119
rect 4905 17085 4939 17119
rect 5273 17085 5307 17119
rect 5733 17085 5767 17119
rect 6929 17085 6963 17119
rect 7297 17085 7331 17119
rect 8033 17085 8067 17119
rect 8493 17085 8527 17119
rect 9045 17085 9079 17119
rect 9229 17085 9263 17119
rect 10701 17085 10735 17119
rect 14565 17085 14599 17119
rect 15117 17085 15151 17119
rect 8953 17017 8987 17051
rect 14841 17017 14875 17051
rect 3893 16949 3927 16983
rect 5457 16949 5491 16983
rect 6101 16949 6135 16983
rect 6469 16949 6503 16983
rect 6653 16949 6687 16983
rect 7941 16949 7975 16983
rect 10057 16949 10091 16983
rect 11161 16949 11195 16983
rect 2513 16745 2547 16779
rect 3249 16745 3283 16779
rect 4261 16745 4295 16779
rect 4997 16745 5031 16779
rect 7389 16745 7423 16779
rect 8217 16745 8251 16779
rect 13093 16745 13127 16779
rect 2145 16677 2179 16711
rect 9321 16677 9355 16711
rect 11682 16677 11716 16711
rect 14933 16677 14967 16711
rect 1869 16609 1903 16643
rect 3065 16609 3099 16643
rect 3433 16609 3467 16643
rect 4077 16609 4111 16643
rect 4445 16609 4479 16643
rect 4813 16609 4847 16643
rect 5632 16609 5666 16643
rect 6837 16609 6871 16643
rect 7205 16609 7239 16643
rect 7665 16609 7699 16643
rect 8033 16609 8067 16643
rect 8861 16609 8895 16643
rect 9956 16609 9990 16643
rect 11437 16609 11471 16643
rect 12909 16609 12943 16643
rect 13277 16609 13311 16643
rect 14381 16609 14415 16643
rect 14657 16609 14691 16643
rect 3801 16541 3835 16575
rect 5365 16541 5399 16575
rect 8953 16541 8987 16575
rect 9137 16541 9171 16575
rect 9689 16541 9723 16575
rect 11161 16541 11195 16575
rect 3617 16473 3651 16507
rect 4629 16473 4663 16507
rect 7021 16473 7055 16507
rect 7849 16473 7883 16507
rect 11069 16473 11103 16507
rect 12817 16473 12851 16507
rect 5181 16405 5215 16439
rect 6745 16405 6779 16439
rect 8493 16405 8527 16439
rect 6009 16201 6043 16235
rect 6653 16201 6687 16235
rect 10609 16201 10643 16235
rect 11805 16133 11839 16167
rect 1777 16065 1811 16099
rect 7389 16065 7423 16099
rect 10885 16065 10919 16099
rect 11437 16065 11471 16099
rect 11621 16065 11655 16099
rect 13001 16065 13035 16099
rect 1593 15997 1627 16031
rect 3157 15997 3191 16031
rect 4629 15997 4663 16031
rect 7757 15997 7791 16031
rect 9229 15997 9263 16031
rect 11345 15997 11379 16031
rect 3402 15929 3436 15963
rect 4874 15929 4908 15963
rect 6285 15929 6319 15963
rect 8024 15929 8058 15963
rect 9496 15929 9530 15963
rect 12909 15929 12943 15963
rect 2237 15861 2271 15895
rect 4537 15861 4571 15895
rect 6469 15861 6503 15895
rect 6837 15861 6871 15895
rect 7205 15861 7239 15895
rect 7297 15861 7331 15895
rect 9137 15861 9171 15895
rect 10977 15861 11011 15895
rect 12449 15861 12483 15895
rect 12817 15861 12851 15895
rect 2789 15657 2823 15691
rect 5917 15657 5951 15691
rect 8677 15657 8711 15691
rect 9045 15657 9079 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 10977 15657 11011 15691
rect 5181 15589 5215 15623
rect 6714 15589 6748 15623
rect 8125 15589 8159 15623
rect 12633 15589 12667 15623
rect 14381 15589 14415 15623
rect 1501 15521 1535 15555
rect 2605 15521 2639 15555
rect 2973 15521 3007 15555
rect 3525 15521 3559 15555
rect 4445 15521 4479 15555
rect 5825 15521 5859 15555
rect 8585 15521 8619 15555
rect 10057 15521 10091 15555
rect 11345 15521 11379 15555
rect 12173 15521 12207 15555
rect 12817 15521 12851 15555
rect 14105 15521 14139 15555
rect 1685 15453 1719 15487
rect 3617 15453 3651 15487
rect 3801 15453 3835 15487
rect 4537 15453 4571 15487
rect 4721 15453 4755 15487
rect 6101 15453 6135 15487
rect 6469 15453 6503 15487
rect 9137 15453 9171 15487
rect 9321 15453 9355 15487
rect 10241 15453 10275 15487
rect 10609 15453 10643 15487
rect 11437 15453 11471 15487
rect 11621 15453 11655 15487
rect 12265 15453 12299 15487
rect 12357 15453 12391 15487
rect 3157 15385 3191 15419
rect 4077 15385 4111 15419
rect 7941 15385 7975 15419
rect 8401 15385 8435 15419
rect 4997 15317 5031 15351
rect 5457 15317 5491 15351
rect 6285 15317 6319 15351
rect 7849 15317 7883 15351
rect 10793 15317 10827 15351
rect 11805 15317 11839 15351
rect 14749 15317 14783 15351
rect 3709 15113 3743 15147
rect 3801 15113 3835 15147
rect 5825 15113 5859 15147
rect 8493 15113 8527 15147
rect 10149 15113 10183 15147
rect 4997 15045 5031 15079
rect 10977 15045 11011 15079
rect 4353 14977 4387 15011
rect 5549 14977 5583 15011
rect 6377 14977 6411 15011
rect 7389 14977 7423 15011
rect 8217 14977 8251 15011
rect 9045 14977 9079 15011
rect 9873 14977 9907 15011
rect 10701 14977 10735 15011
rect 11437 14977 11471 15011
rect 11621 14977 11655 15011
rect 13001 14977 13035 15011
rect 1501 14909 1535 14943
rect 1777 14909 1811 14943
rect 2329 14909 2363 14943
rect 5365 14909 5399 14943
rect 6285 14909 6319 14943
rect 8033 14909 8067 14943
rect 9781 14909 9815 14943
rect 2596 14841 2630 14875
rect 4169 14841 4203 14875
rect 4813 14841 4847 14875
rect 6193 14841 6227 14875
rect 8953 14841 8987 14875
rect 10517 14841 10551 14875
rect 11989 14841 12023 14875
rect 12909 14841 12943 14875
rect 4261 14773 4295 14807
rect 4629 14773 4663 14807
rect 5457 14773 5491 14807
rect 6837 14773 6871 14807
rect 7205 14773 7239 14807
rect 7297 14773 7331 14807
rect 7665 14773 7699 14807
rect 8125 14773 8159 14807
rect 8861 14773 8895 14807
rect 9321 14773 9355 14807
rect 9689 14773 9723 14807
rect 10609 14773 10643 14807
rect 11345 14773 11379 14807
rect 11805 14773 11839 14807
rect 12449 14773 12483 14807
rect 12817 14773 12851 14807
rect 13277 14773 13311 14807
rect 3157 14569 3191 14603
rect 4077 14569 4111 14603
rect 4445 14569 4479 14603
rect 5365 14569 5399 14603
rect 5825 14569 5859 14603
rect 6193 14569 6227 14603
rect 6653 14569 6687 14603
rect 7021 14569 7055 14603
rect 8953 14569 8987 14603
rect 9321 14569 9355 14603
rect 12357 14569 12391 14603
rect 13185 14569 13219 14603
rect 13553 14569 13587 14603
rect 6561 14501 6595 14535
rect 7840 14501 7874 14535
rect 9137 14501 9171 14535
rect 10149 14501 10183 14535
rect 10876 14501 10910 14535
rect 13645 14501 13679 14535
rect 14381 14501 14415 14535
rect 1501 14433 1535 14467
rect 3065 14433 3099 14467
rect 5089 14433 5123 14467
rect 5733 14433 5767 14467
rect 7573 14433 7607 14467
rect 10057 14433 10091 14467
rect 12725 14433 12759 14467
rect 1685 14365 1719 14399
rect 3249 14365 3283 14399
rect 4537 14365 4571 14399
rect 4629 14365 4663 14399
rect 5917 14365 5951 14399
rect 6745 14365 6779 14399
rect 10241 14365 10275 14399
rect 10609 14365 10643 14399
rect 12817 14365 12851 14399
rect 12909 14365 12943 14399
rect 13737 14365 13771 14399
rect 7297 14297 7331 14331
rect 9689 14297 9723 14331
rect 14197 14297 14231 14331
rect 2697 14229 2731 14263
rect 4905 14229 4939 14263
rect 5181 14229 5215 14263
rect 11989 14229 12023 14263
rect 14013 14229 14047 14263
rect 4077 14025 4111 14059
rect 8309 14025 8343 14059
rect 10149 14025 10183 14059
rect 10793 14025 10827 14059
rect 6101 13957 6135 13991
rect 8769 13957 8803 13991
rect 2697 13889 2731 13923
rect 4721 13889 4755 13923
rect 5917 13889 5951 13923
rect 6929 13889 6963 13923
rect 11529 13889 11563 13923
rect 1593 13821 1627 13855
rect 1869 13821 1903 13855
rect 2964 13821 2998 13855
rect 4629 13821 4663 13855
rect 6377 13821 6411 13855
rect 8585 13821 8619 13855
rect 10517 13821 10551 13855
rect 12449 13821 12483 13855
rect 12705 13821 12739 13855
rect 5641 13753 5675 13787
rect 7196 13753 7230 13787
rect 8861 13753 8895 13787
rect 11253 13753 11287 13787
rect 4169 13685 4203 13719
rect 4537 13685 4571 13719
rect 4997 13685 5031 13719
rect 5273 13685 5307 13719
rect 5733 13685 5767 13719
rect 6561 13685 6595 13719
rect 10885 13685 10919 13719
rect 11345 13685 11379 13719
rect 13829 13685 13863 13719
rect 3157 13481 3191 13515
rect 4353 13481 4387 13515
rect 4813 13481 4847 13515
rect 9321 13481 9355 13515
rect 11161 13481 11195 13515
rect 11621 13481 11655 13515
rect 2044 13413 2078 13447
rect 5448 13413 5482 13447
rect 11529 13413 11563 13447
rect 1777 13345 1811 13379
rect 4721 13345 4755 13379
rect 6745 13345 6779 13379
rect 7012 13345 7046 13379
rect 8861 13345 8895 13379
rect 9505 13345 9539 13379
rect 10701 13345 10735 13379
rect 4077 13277 4111 13311
rect 4905 13277 4939 13311
rect 5181 13277 5215 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 9781 13277 9815 13311
rect 10793 13277 10827 13311
rect 10885 13277 10919 13311
rect 11805 13277 11839 13311
rect 6561 13141 6595 13175
rect 8125 13141 8159 13175
rect 8493 13141 8527 13175
rect 10333 13141 10367 13175
rect 3157 12937 3191 12971
rect 4997 12937 5031 12971
rect 5273 12937 5307 12971
rect 10885 12937 10919 12971
rect 11989 12937 12023 12971
rect 4813 12869 4847 12903
rect 3801 12801 3835 12835
rect 4445 12801 4479 12835
rect 4629 12801 4663 12835
rect 5825 12801 5859 12835
rect 6101 12801 6135 12835
rect 7389 12801 7423 12835
rect 8217 12801 8251 12835
rect 9137 12801 9171 12835
rect 11437 12801 11471 12835
rect 3617 12733 3651 12767
rect 4353 12733 4387 12767
rect 5181 12733 5215 12767
rect 7205 12733 7239 12767
rect 8033 12733 8067 12767
rect 9321 12733 9355 12767
rect 9577 12733 9611 12767
rect 3525 12665 3559 12699
rect 6285 12665 6319 12699
rect 8953 12665 8987 12699
rect 11345 12665 11379 12699
rect 3985 12597 4019 12631
rect 5641 12597 5675 12631
rect 5733 12597 5767 12631
rect 6837 12597 6871 12631
rect 7297 12597 7331 12631
rect 7665 12597 7699 12631
rect 8125 12597 8159 12631
rect 8493 12597 8527 12631
rect 8861 12597 8895 12631
rect 10701 12597 10735 12631
rect 11253 12597 11287 12631
rect 11805 12597 11839 12631
rect 7389 12393 7423 12427
rect 7941 12393 7975 12427
rect 8769 12393 8803 12427
rect 9137 12393 9171 12427
rect 9689 12393 9723 12427
rect 11345 12393 11379 12427
rect 12541 12393 12575 12427
rect 1777 12325 1811 12359
rect 8401 12325 8435 12359
rect 9229 12325 9263 12359
rect 1511 12257 1545 12291
rect 5457 12257 5491 12291
rect 6184 12257 6218 12291
rect 7573 12257 7607 12291
rect 7849 12257 7883 12291
rect 8309 12257 8343 12291
rect 10140 12257 10174 12291
rect 11713 12257 11747 12291
rect 12173 12257 12207 12291
rect 5549 12189 5583 12223
rect 5733 12189 5767 12223
rect 5917 12189 5951 12223
rect 8585 12189 8619 12223
rect 9321 12189 9355 12223
rect 9873 12189 9907 12223
rect 11805 12189 11839 12223
rect 11897 12189 11931 12223
rect 11253 12121 11287 12155
rect 5089 12053 5123 12087
rect 7297 12053 7331 12087
rect 9137 11849 9171 11883
rect 8585 11781 8619 11815
rect 9781 11713 9815 11747
rect 10241 11713 10275 11747
rect 1501 11645 1535 11679
rect 2053 11645 2087 11679
rect 3249 11645 3283 11679
rect 4721 11645 4755 11679
rect 7205 11645 7239 11679
rect 7461 11645 7495 11679
rect 8769 11645 8803 11679
rect 9045 11645 9079 11679
rect 9597 11645 9631 11679
rect 1777 11577 1811 11611
rect 2329 11577 2363 11611
rect 3516 11577 3550 11611
rect 4988 11577 5022 11611
rect 9965 11577 9999 11611
rect 3157 11509 3191 11543
rect 4629 11509 4663 11543
rect 6101 11509 6135 11543
rect 6653 11509 6687 11543
rect 6837 11509 6871 11543
rect 9505 11509 9539 11543
rect 1501 11305 1535 11339
rect 3801 11305 3835 11339
rect 4537 11305 4571 11339
rect 5181 11305 5215 11339
rect 5825 11305 5859 11339
rect 6377 11305 6411 11339
rect 6837 11305 6871 11339
rect 7665 11305 7699 11339
rect 8861 11305 8895 11339
rect 9689 11305 9723 11339
rect 8309 11237 8343 11271
rect 1869 11169 1903 11203
rect 2677 11169 2711 11203
rect 4445 11169 4479 11203
rect 5089 11169 5123 11203
rect 5917 11169 5951 11203
rect 7757 11169 7791 11203
rect 8769 11169 8803 11203
rect 9413 11169 9447 11203
rect 9873 11169 9907 11203
rect 10609 11169 10643 11203
rect 11345 11169 11379 11203
rect 11612 11169 11646 11203
rect 1961 11101 1995 11135
rect 2145 11101 2179 11135
rect 2421 11101 2455 11135
rect 4629 11101 4663 11135
rect 6101 11101 6135 11135
rect 6929 11101 6963 11135
rect 7113 11101 7147 11135
rect 7849 11101 7883 11135
rect 9045 11101 9079 11135
rect 10701 11101 10735 11135
rect 10885 11101 10919 11135
rect 4077 11033 4111 11067
rect 4905 11033 4939 11067
rect 5457 11033 5491 11067
rect 6469 11033 6503 11067
rect 10241 11033 10275 11067
rect 7297 10965 7331 10999
rect 8401 10965 8435 10999
rect 9229 10965 9263 10999
rect 12725 10965 12759 10999
rect 1501 10761 1535 10795
rect 3985 10761 4019 10795
rect 5181 10761 5215 10795
rect 6837 10761 6871 10795
rect 6377 10693 6411 10727
rect 11345 10693 11379 10727
rect 2145 10625 2179 10659
rect 2789 10625 2823 10659
rect 2973 10625 3007 10659
rect 3709 10625 3743 10659
rect 4445 10625 4479 10659
rect 4629 10625 4663 10659
rect 5825 10625 5859 10659
rect 7389 10625 7423 10659
rect 8217 10625 8251 10659
rect 8493 10625 8527 10659
rect 9965 10625 9999 10659
rect 11897 10625 11931 10659
rect 11989 10625 12023 10659
rect 13001 10625 13035 10659
rect 3525 10557 3559 10591
rect 5089 10557 5123 10591
rect 5549 10557 5583 10591
rect 7205 10557 7239 10591
rect 8125 10557 8159 10591
rect 10232 10557 10266 10591
rect 1869 10489 1903 10523
rect 2697 10489 2731 10523
rect 3617 10489 3651 10523
rect 5641 10489 5675 10523
rect 8760 10489 8794 10523
rect 11805 10489 11839 10523
rect 12909 10489 12943 10523
rect 1961 10421 1995 10455
rect 2329 10421 2363 10455
rect 3157 10421 3191 10455
rect 4353 10421 4387 10455
rect 4905 10421 4939 10455
rect 6101 10421 6135 10455
rect 6561 10421 6595 10455
rect 7297 10421 7331 10455
rect 7665 10421 7699 10455
rect 8033 10421 8067 10455
rect 9873 10421 9907 10455
rect 11437 10421 11471 10455
rect 12449 10421 12483 10455
rect 12817 10421 12851 10455
rect 13277 10421 13311 10455
rect 2973 10217 3007 10251
rect 3617 10217 3651 10251
rect 4261 10217 4295 10251
rect 4629 10217 4663 10251
rect 6837 10217 6871 10251
rect 12173 10217 12207 10251
rect 13001 10217 13035 10251
rect 13369 10217 13403 10251
rect 13461 10217 13495 10251
rect 14289 10217 14323 10251
rect 3525 10149 3559 10183
rect 4169 10149 4203 10183
rect 5610 10149 5644 10183
rect 10600 10149 10634 10183
rect 14013 10149 14047 10183
rect 1593 10081 1627 10115
rect 1860 10081 1894 10115
rect 4721 10081 4755 10115
rect 5365 10081 5399 10115
rect 7113 10081 7147 10115
rect 10333 10081 10367 10115
rect 12541 10081 12575 10115
rect 12633 10081 12667 10115
rect 3801 10013 3835 10047
rect 4905 10013 4939 10047
rect 12725 10013 12759 10047
rect 13553 10013 13587 10047
rect 13829 9945 13863 9979
rect 3157 9877 3191 9911
rect 5089 9877 5123 9911
rect 6745 9877 6779 9911
rect 8401 9877 8435 9911
rect 11713 9877 11747 9911
rect 11897 9673 11931 9707
rect 6469 9605 6503 9639
rect 8493 9605 8527 9639
rect 10057 9605 10091 9639
rect 10885 9605 10919 9639
rect 3709 9537 3743 9571
rect 4905 9537 4939 9571
rect 9137 9537 9171 9571
rect 10701 9537 10735 9571
rect 11529 9537 11563 9571
rect 15301 9537 15335 9571
rect 1501 9469 1535 9503
rect 2053 9469 2087 9503
rect 3525 9469 3559 9503
rect 4169 9469 4203 9503
rect 5089 9469 5123 9503
rect 5356 9469 5390 9503
rect 6653 9469 6687 9503
rect 6837 9469 6871 9503
rect 8953 9469 8987 9503
rect 9321 9469 9355 9503
rect 11253 9469 11287 9503
rect 15025 9469 15059 9503
rect 1777 9401 1811 9435
rect 2320 9401 2354 9435
rect 7104 9401 7138 9435
rect 8401 9401 8435 9435
rect 11345 9401 11379 9435
rect 11713 9401 11747 9435
rect 3433 9333 3467 9367
rect 4261 9333 4295 9367
rect 4629 9333 4663 9367
rect 4721 9333 4755 9367
rect 6653 9333 6687 9367
rect 8217 9333 8251 9367
rect 8861 9333 8895 9367
rect 9505 9333 9539 9367
rect 9781 9333 9815 9367
rect 9965 9333 9999 9367
rect 10425 9333 10459 9367
rect 10517 9333 10551 9367
rect 14841 9333 14875 9367
rect 1501 9129 1535 9163
rect 2329 9129 2363 9163
rect 3157 9129 3191 9163
rect 3525 9129 3559 9163
rect 4721 9129 4755 9163
rect 5181 9129 5215 9163
rect 5549 9129 5583 9163
rect 6837 9129 6871 9163
rect 7297 9129 7331 9163
rect 7665 9129 7699 9163
rect 10057 9129 10091 9163
rect 10425 9129 10459 9163
rect 11253 9129 11287 9163
rect 13093 9129 13127 9163
rect 1961 9061 1995 9095
rect 4077 9061 4111 9095
rect 5089 9061 5123 9095
rect 6929 9061 6963 9095
rect 1869 8993 1903 9027
rect 2697 8993 2731 9027
rect 2789 8993 2823 9027
rect 5917 8993 5951 9027
rect 8392 8993 8426 9027
rect 10517 8993 10551 9027
rect 11345 8993 11379 9027
rect 11980 8993 12014 9027
rect 2145 8925 2179 8959
rect 2927 8925 2961 8959
rect 3617 8925 3651 8959
rect 3709 8925 3743 8959
rect 5365 8925 5399 8959
rect 6009 8925 6043 8959
rect 6193 8925 6227 8959
rect 7113 8925 7147 8959
rect 7757 8925 7791 8959
rect 7941 8925 7975 8959
rect 8125 8925 8159 8959
rect 9689 8925 9723 8959
rect 10701 8925 10735 8959
rect 11529 8925 11563 8959
rect 11713 8925 11747 8959
rect 6469 8857 6503 8891
rect 10885 8857 10919 8891
rect 4353 8789 4387 8823
rect 4537 8789 4571 8823
rect 9505 8789 9539 8823
rect 8677 8585 8711 8619
rect 9505 8585 9539 8619
rect 10977 8585 11011 8619
rect 4445 8517 4479 8551
rect 6469 8517 6503 8551
rect 7021 8517 7055 8551
rect 7849 8517 7883 8551
rect 10333 8517 10367 8551
rect 10793 8517 10827 8551
rect 11805 8517 11839 8551
rect 12449 8517 12483 8551
rect 2145 8449 2179 8483
rect 5089 8449 5123 8483
rect 7665 8449 7699 8483
rect 8401 8449 8435 8483
rect 9229 8449 9263 8483
rect 10149 8449 10183 8483
rect 11437 8449 11471 8483
rect 11621 8449 11655 8483
rect 13001 8449 13035 8483
rect 1593 8381 1627 8415
rect 3065 8381 3099 8415
rect 4721 8381 4755 8415
rect 5356 8381 5390 8415
rect 7481 8381 7515 8415
rect 9965 8381 9999 8415
rect 10517 8381 10551 8415
rect 10701 8381 10735 8415
rect 12081 8381 12115 8415
rect 12817 8381 12851 8415
rect 3332 8313 3366 8347
rect 9137 8313 9171 8347
rect 9873 8313 9907 8347
rect 11345 8313 11379 8347
rect 12173 8313 12207 8347
rect 13369 8313 13403 8347
rect 4537 8245 4571 8279
rect 6653 8245 6687 8279
rect 6929 8245 6963 8279
rect 7389 8245 7423 8279
rect 8217 8245 8251 8279
rect 8309 8245 8343 8279
rect 9045 8245 9079 8279
rect 12909 8245 12943 8279
rect 1501 8041 1535 8075
rect 5549 8041 5583 8075
rect 8033 8041 8067 8075
rect 8125 8041 8159 8075
rect 8493 8041 8527 8075
rect 8953 8041 8987 8075
rect 9689 8041 9723 8075
rect 9965 8041 9999 8075
rect 14105 8041 14139 8075
rect 8585 7973 8619 8007
rect 1961 7905 1995 7939
rect 2228 7905 2262 7939
rect 4445 7905 4479 7939
rect 5917 7905 5951 7939
rect 6561 7905 6595 7939
rect 6920 7905 6954 7939
rect 9229 7905 9263 7939
rect 10701 7905 10735 7939
rect 11253 7905 11287 7939
rect 11509 7905 11543 7939
rect 12725 7905 12759 7939
rect 12981 7905 13015 7939
rect 4537 7837 4571 7871
rect 4629 7837 4663 7871
rect 4905 7837 4939 7871
rect 5457 7837 5491 7871
rect 6009 7837 6043 7871
rect 6193 7837 6227 7871
rect 6653 7837 6687 7871
rect 8769 7837 8803 7871
rect 10793 7837 10827 7871
rect 10977 7837 11011 7871
rect 3341 7769 3375 7803
rect 4077 7701 4111 7735
rect 5181 7701 5215 7735
rect 6377 7701 6411 7735
rect 9413 7701 9447 7735
rect 10333 7701 10367 7735
rect 12633 7701 12667 7735
rect 3893 7497 3927 7531
rect 4721 7497 4755 7531
rect 5825 7497 5859 7531
rect 11437 7497 11471 7531
rect 1685 7361 1719 7395
rect 3341 7361 3375 7395
rect 4445 7361 4479 7395
rect 5273 7361 5307 7395
rect 6469 7361 6503 7395
rect 7389 7361 7423 7395
rect 11161 7361 11195 7395
rect 11989 7361 12023 7395
rect 1501 7293 1535 7327
rect 5089 7293 5123 7327
rect 5181 7293 5215 7327
rect 5641 7293 5675 7327
rect 7205 7293 7239 7327
rect 7297 7293 7331 7327
rect 7665 7293 7699 7327
rect 7932 7293 7966 7327
rect 9137 7293 9171 7327
rect 11069 7293 11103 7327
rect 3065 7225 3099 7259
rect 4353 7225 4387 7259
rect 6193 7225 6227 7259
rect 9382 7225 9416 7259
rect 10977 7225 11011 7259
rect 11805 7225 11839 7259
rect 2697 7157 2731 7191
rect 3157 7157 3191 7191
rect 4261 7157 4295 7191
rect 6285 7157 6319 7191
rect 6837 7157 6871 7191
rect 9045 7157 9079 7191
rect 10517 7157 10551 7191
rect 10609 7157 10643 7191
rect 11897 7157 11931 7191
rect 2605 6953 2639 6987
rect 2973 6953 3007 6987
rect 3341 6953 3375 6987
rect 3801 6953 3835 6987
rect 4077 6953 4111 6987
rect 5457 6953 5491 6987
rect 6561 6953 6595 6987
rect 8125 6953 8159 6987
rect 8309 6953 8343 6987
rect 9229 6953 9263 6987
rect 11437 6953 11471 6987
rect 11621 6953 11655 6987
rect 12449 6953 12483 6987
rect 2513 6885 2547 6919
rect 4537 6885 4571 6919
rect 11253 6885 11287 6919
rect 11989 6885 12023 6919
rect 1501 6817 1535 6851
rect 3433 6817 3467 6851
rect 4445 6817 4479 6851
rect 5089 6817 5123 6851
rect 5917 6817 5951 6851
rect 6009 6817 6043 6851
rect 7012 6817 7046 6851
rect 8677 6817 8711 6851
rect 9137 6817 9171 6851
rect 9781 6817 9815 6851
rect 10037 6817 10071 6851
rect 12081 6817 12115 6851
rect 12817 6817 12851 6851
rect 13645 6817 13679 6851
rect 1685 6749 1719 6783
rect 2789 6749 2823 6783
rect 3525 6749 3559 6783
rect 4629 6749 4663 6783
rect 6101 6749 6135 6783
rect 6745 6749 6779 6783
rect 9321 6749 9355 6783
rect 12173 6749 12207 6783
rect 12909 6749 12943 6783
rect 13001 6749 13035 6783
rect 8493 6681 8527 6715
rect 13461 6681 13495 6715
rect 2145 6613 2179 6647
rect 4905 6613 4939 6647
rect 5273 6613 5307 6647
rect 5549 6613 5583 6647
rect 6377 6613 6411 6647
rect 8769 6613 8803 6647
rect 11161 6613 11195 6647
rect 13277 6613 13311 6647
rect 4537 6409 4571 6443
rect 6837 6409 6871 6443
rect 7849 6409 7883 6443
rect 8125 6409 8159 6443
rect 10241 6409 10275 6443
rect 6009 6341 6043 6375
rect 3157 6273 3191 6307
rect 6193 6273 6227 6307
rect 7481 6273 7515 6307
rect 8861 6273 8895 6307
rect 9045 6273 9079 6307
rect 9689 6273 9723 6307
rect 9873 6273 9907 6307
rect 10885 6273 10919 6307
rect 12081 6273 12115 6307
rect 1501 6205 1535 6239
rect 4629 6205 4663 6239
rect 4896 6205 4930 6239
rect 8769 6205 8803 6239
rect 9597 6205 9631 6239
rect 10609 6205 10643 6239
rect 1777 6137 1811 6171
rect 3424 6137 3458 6171
rect 6561 6137 6595 6171
rect 8217 6137 8251 6171
rect 10701 6137 10735 6171
rect 7205 6069 7239 6103
rect 7297 6069 7331 6103
rect 7757 6069 7791 6103
rect 8401 6069 8435 6103
rect 9229 6069 9263 6103
rect 10057 6069 10091 6103
rect 4077 5865 4111 5899
rect 4537 5865 4571 5899
rect 7021 5865 7055 5899
rect 7481 5865 7515 5899
rect 7849 5865 7883 5899
rect 8309 5865 8343 5899
rect 8677 5865 8711 5899
rect 9137 5865 9171 5899
rect 9689 5865 9723 5899
rect 10241 5865 10275 5899
rect 3617 5797 3651 5831
rect 5724 5797 5758 5831
rect 10149 5797 10183 5831
rect 10762 5797 10796 5831
rect 2053 5729 2087 5763
rect 2320 5729 2354 5763
rect 4445 5729 4479 5763
rect 5181 5729 5215 5763
rect 7389 5729 7423 5763
rect 8217 5729 8251 5763
rect 9045 5729 9079 5763
rect 10517 5729 10551 5763
rect 4629 5661 4663 5695
rect 5457 5661 5491 5695
rect 7573 5661 7607 5695
rect 8401 5661 8435 5695
rect 9321 5661 9355 5695
rect 3433 5593 3467 5627
rect 6837 5593 6871 5627
rect 4997 5525 5031 5559
rect 9873 5525 9907 5559
rect 11897 5525 11931 5559
rect 6101 5321 6135 5355
rect 6377 5321 6411 5355
rect 8217 5321 8251 5355
rect 8401 5321 8435 5355
rect 14841 5321 14875 5355
rect 6285 5253 6319 5287
rect 2237 5185 2271 5219
rect 6653 5185 6687 5219
rect 13093 5185 13127 5219
rect 1501 5117 1535 5151
rect 2053 5117 2087 5151
rect 2881 5117 2915 5151
rect 4537 5117 4571 5151
rect 4721 5117 4755 5151
rect 6837 5117 6871 5151
rect 8585 5117 8619 5151
rect 8852 5117 8886 5151
rect 10057 5117 10091 5151
rect 12909 5117 12943 5151
rect 13553 5117 13587 5151
rect 15025 5117 15059 5151
rect 1777 5049 1811 5083
rect 3148 5049 3182 5083
rect 4988 5049 5022 5083
rect 7104 5049 7138 5083
rect 10324 5049 10358 5083
rect 12817 5049 12851 5083
rect 13277 5049 13311 5083
rect 15301 5049 15335 5083
rect 4261 4981 4295 5015
rect 4353 4981 4387 5015
rect 9965 4981 9999 5015
rect 11437 4981 11471 5015
rect 12449 4981 12483 5015
rect 2789 4777 2823 4811
rect 3617 4777 3651 4811
rect 4353 4777 4387 4811
rect 4813 4777 4847 4811
rect 5181 4777 5215 4811
rect 5641 4777 5675 4811
rect 6561 4777 6595 4811
rect 6653 4777 6687 4811
rect 7941 4777 7975 4811
rect 8401 4777 8435 4811
rect 8769 4777 8803 4811
rect 9229 4777 9263 4811
rect 9965 4777 9999 4811
rect 10241 4777 10275 4811
rect 13185 4777 13219 4811
rect 13645 4777 13679 4811
rect 13921 4777 13955 4811
rect 3525 4709 3559 4743
rect 13277 4709 13311 4743
rect 1409 4641 1443 4675
rect 1676 4641 1710 4675
rect 4261 4641 4295 4675
rect 4721 4641 4755 4675
rect 5549 4641 5583 4675
rect 6101 4641 6135 4675
rect 7021 4641 7055 4675
rect 7849 4641 7883 4675
rect 8309 4641 8343 4675
rect 9137 4641 9171 4675
rect 9873 4641 9907 4675
rect 10793 4641 10827 4675
rect 11345 4641 11379 4675
rect 11612 4641 11646 4675
rect 3709 4573 3743 4607
rect 4905 4573 4939 4607
rect 5733 4573 5767 4607
rect 7113 4573 7147 4607
rect 7297 4573 7331 4607
rect 7481 4573 7515 4607
rect 8585 4573 8619 4607
rect 9321 4573 9355 4607
rect 10885 4573 10919 4607
rect 10977 4573 11011 4607
rect 13369 4573 13403 4607
rect 2973 4437 3007 4471
rect 3157 4437 3191 4471
rect 6285 4437 6319 4471
rect 9689 4437 9723 4471
rect 10425 4437 10459 4471
rect 12725 4437 12759 4471
rect 12817 4437 12851 4471
rect 2145 4233 2179 4267
rect 9965 4233 9999 4267
rect 10793 4233 10827 4267
rect 2421 4165 2455 4199
rect 9873 4165 9907 4199
rect 2973 4097 3007 4131
rect 3985 4097 4019 4131
rect 4997 4097 5031 4131
rect 5273 4097 5307 4131
rect 6469 4097 6503 4131
rect 7297 4097 7331 4131
rect 7481 4097 7515 4131
rect 8401 4097 8435 4131
rect 9137 4097 9171 4131
rect 10425 4097 10459 4131
rect 10609 4097 10643 4131
rect 11437 4097 11471 4131
rect 12909 4097 12943 4131
rect 13001 4097 13035 4131
rect 1501 4029 1535 4063
rect 2789 4029 2823 4063
rect 3341 4029 3375 4063
rect 4353 4029 4387 4063
rect 5549 4029 5583 4063
rect 7205 4029 7239 4063
rect 9689 4029 9723 4063
rect 11161 4029 11195 4063
rect 1777 3961 1811 3995
rect 2881 3961 2915 3995
rect 3801 3961 3835 3995
rect 6285 3961 6319 3995
rect 8217 3961 8251 3995
rect 10333 3961 10367 3995
rect 12817 3961 12851 3995
rect 2329 3893 2363 3927
rect 3433 3893 3467 3927
rect 3893 3893 3927 3927
rect 4445 3893 4479 3927
rect 4813 3893 4847 3927
rect 4905 3893 4939 3927
rect 5733 3893 5767 3927
rect 5917 3893 5951 3927
rect 6377 3893 6411 3927
rect 6837 3893 6871 3927
rect 7757 3893 7791 3927
rect 8125 3893 8159 3927
rect 8585 3893 8619 3927
rect 8953 3893 8987 3927
rect 9045 3893 9079 3927
rect 9413 3893 9447 3927
rect 11253 3893 11287 3927
rect 11713 3893 11747 3927
rect 12449 3893 12483 3927
rect 2605 3689 2639 3723
rect 3709 3689 3743 3723
rect 7573 3689 7607 3723
rect 9689 3689 9723 3723
rect 10149 3689 10183 3723
rect 10701 3689 10735 3723
rect 12909 3689 12943 3723
rect 1501 3553 1535 3587
rect 2053 3553 2087 3587
rect 1685 3485 1719 3519
rect 3893 3621 3927 3655
rect 5908 3621 5942 3655
rect 7481 3621 7515 3655
rect 8370 3621 8404 3655
rect 9873 3621 9907 3655
rect 3065 3553 3099 3587
rect 4353 3553 4387 3587
rect 4813 3553 4847 3587
rect 4905 3553 4939 3587
rect 5279 3553 5313 3587
rect 8125 3553 8159 3587
rect 11069 3553 11103 3587
rect 11529 3553 11563 3587
rect 11785 3553 11819 3587
rect 2973 3485 3007 3519
rect 4169 3485 4203 3519
rect 5089 3485 5123 3519
rect 5641 3485 5675 3519
rect 7757 3485 7791 3519
rect 10425 3485 10459 3519
rect 11161 3485 11195 3519
rect 11253 3485 11287 3519
rect 2421 3417 2455 3451
rect 2605 3417 2639 3451
rect 3249 3417 3283 3451
rect 3525 3417 3559 3451
rect 7113 3417 7147 3451
rect 7941 3417 7975 3451
rect 2237 3349 2271 3383
rect 2789 3349 2823 3383
rect 4445 3349 4479 3383
rect 5457 3349 5491 3383
rect 7021 3349 7055 3383
rect 9505 3349 9539 3383
rect 10333 3349 10367 3383
rect 4445 3145 4479 3179
rect 5365 3145 5399 3179
rect 6653 3145 6687 3179
rect 8309 3145 8343 3179
rect 9229 3145 9263 3179
rect 10977 3145 11011 3179
rect 12449 3145 12483 3179
rect 6377 3077 6411 3111
rect 8217 3077 8251 3111
rect 10793 3077 10827 3111
rect 5089 3009 5123 3043
rect 5917 3009 5951 3043
rect 6837 3009 6871 3043
rect 8861 3009 8895 3043
rect 9413 3009 9447 3043
rect 11529 3009 11563 3043
rect 13001 3009 13035 3043
rect 14565 3009 14599 3043
rect 1593 2941 1627 2975
rect 3065 2941 3099 2975
rect 4997 2941 5031 2975
rect 6193 2941 6227 2975
rect 7104 2941 7138 2975
rect 14289 2941 14323 2975
rect 14841 2941 14875 2975
rect 15393 2941 15427 2975
rect 1501 2873 1535 2907
rect 1838 2873 1872 2907
rect 3310 2873 3344 2907
rect 8677 2873 8711 2907
rect 9658 2873 9692 2907
rect 11437 2873 11471 2907
rect 11805 2873 11839 2907
rect 12173 2873 12207 2907
rect 12909 2873 12943 2907
rect 15117 2873 15151 2907
rect 2973 2805 3007 2839
rect 4537 2805 4571 2839
rect 4905 2805 4939 2839
rect 5733 2805 5767 2839
rect 5825 2805 5859 2839
rect 8769 2805 8803 2839
rect 11345 2805 11379 2839
rect 11989 2805 12023 2839
rect 12817 2805 12851 2839
rect 13277 2805 13311 2839
rect 15577 2805 15611 2839
rect 2145 2601 2179 2635
rect 2513 2601 2547 2635
rect 4077 2601 4111 2635
rect 4537 2601 4571 2635
rect 5825 2601 5859 2635
rect 6377 2601 6411 2635
rect 6929 2601 6963 2635
rect 7389 2601 7423 2635
rect 8217 2601 8251 2635
rect 8585 2601 8619 2635
rect 9045 2601 9079 2635
rect 10057 2601 10091 2635
rect 10977 2601 11011 2635
rect 12449 2601 12483 2635
rect 12817 2601 12851 2635
rect 13001 2601 13035 2635
rect 15485 2601 15519 2635
rect 4445 2533 4479 2567
rect 8125 2533 8159 2567
rect 9413 2533 9447 2567
rect 11989 2533 12023 2567
rect 14381 2533 14415 2567
rect 1501 2465 1535 2499
rect 1593 2465 1627 2499
rect 1961 2465 1995 2499
rect 2329 2465 2363 2499
rect 2697 2465 2731 2499
rect 3157 2465 3191 2499
rect 3525 2465 3559 2499
rect 4905 2465 4939 2499
rect 5273 2465 5307 2499
rect 5641 2465 5675 2499
rect 6009 2465 6043 2499
rect 6193 2465 6227 2499
rect 7297 2465 7331 2499
rect 8953 2465 8987 2499
rect 9873 2465 9907 2499
rect 10241 2465 10275 2499
rect 10609 2465 10643 2499
rect 11345 2465 11379 2499
rect 12173 2465 12207 2499
rect 12633 2465 12667 2499
rect 14105 2465 14139 2499
rect 14657 2465 14691 2499
rect 15209 2465 15243 2499
rect 4721 2397 4755 2431
rect 6561 2397 6595 2431
rect 7573 2397 7607 2431
rect 8309 2397 8343 2431
rect 9137 2397 9171 2431
rect 11437 2397 11471 2431
rect 11621 2397 11655 2431
rect 14933 2397 14967 2431
rect 1777 2329 1811 2363
rect 2881 2329 2915 2363
rect 3709 2329 3743 2363
rect 5457 2329 5491 2363
rect 3341 2261 3375 2295
rect 5089 2261 5123 2295
rect 7757 2261 7791 2295
rect 10425 2261 10459 2295
rect 10793 2261 10827 2295
rect 11805 2261 11839 2295
rect 13185 2261 13219 2295
<< metal1 >>
rect 7558 17688 7564 17740
rect 7616 17728 7622 17740
rect 15010 17728 15016 17740
rect 7616 17700 15016 17728
rect 7616 17688 7622 17700
rect 15010 17688 15016 17700
rect 15068 17688 15074 17740
rect 5258 17620 5264 17672
rect 5316 17660 5322 17672
rect 6362 17660 6368 17672
rect 5316 17632 6368 17660
rect 5316 17620 5322 17632
rect 6362 17620 6368 17632
rect 6420 17660 6426 17672
rect 11974 17660 11980 17672
rect 6420 17632 11980 17660
rect 6420 17620 6426 17632
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 1302 17552 1308 17604
rect 1360 17592 1366 17604
rect 14642 17592 14648 17604
rect 1360 17564 14648 17592
rect 1360 17552 1366 17564
rect 14642 17552 14648 17564
rect 14700 17552 14706 17604
rect 6822 17484 6828 17536
rect 6880 17524 6886 17536
rect 7742 17524 7748 17536
rect 6880 17496 7748 17524
rect 6880 17484 6886 17496
rect 7742 17484 7748 17496
rect 7800 17524 7806 17536
rect 10042 17524 10048 17536
rect 7800 17496 10048 17524
rect 7800 17484 7806 17496
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 1104 17434 16008 17456
rect 1104 17382 3480 17434
rect 3532 17382 3544 17434
rect 3596 17382 3608 17434
rect 3660 17382 3672 17434
rect 3724 17382 8478 17434
rect 8530 17382 8542 17434
rect 8594 17382 8606 17434
rect 8658 17382 8670 17434
rect 8722 17382 13475 17434
rect 13527 17382 13539 17434
rect 13591 17382 13603 17434
rect 13655 17382 13667 17434
rect 13719 17382 16008 17434
rect 1104 17360 16008 17382
rect 4614 17280 4620 17332
rect 4672 17320 4678 17332
rect 5077 17323 5135 17329
rect 5077 17320 5089 17323
rect 4672 17292 5089 17320
rect 4672 17280 4678 17292
rect 5077 17289 5089 17292
rect 5123 17289 5135 17323
rect 5077 17283 5135 17289
rect 5718 17280 5724 17332
rect 5776 17320 5782 17332
rect 5905 17323 5963 17329
rect 5905 17320 5917 17323
rect 5776 17292 5917 17320
rect 5776 17280 5782 17292
rect 5905 17289 5917 17292
rect 5951 17289 5963 17323
rect 6362 17320 6368 17332
rect 6323 17292 6368 17320
rect 5905 17283 5963 17289
rect 6362 17280 6368 17292
rect 6420 17280 6426 17332
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 7101 17323 7159 17329
rect 7101 17320 7113 17323
rect 6972 17292 7113 17320
rect 6972 17280 6978 17292
rect 7101 17289 7113 17292
rect 7147 17289 7159 17323
rect 7101 17283 7159 17289
rect 7282 17280 7288 17332
rect 7340 17320 7346 17332
rect 7469 17323 7527 17329
rect 7469 17320 7481 17323
rect 7340 17292 7481 17320
rect 7340 17280 7346 17292
rect 7469 17289 7481 17292
rect 7515 17289 7527 17323
rect 7742 17320 7748 17332
rect 7703 17292 7748 17320
rect 7469 17283 7527 17289
rect 7742 17280 7748 17292
rect 7800 17280 7806 17332
rect 8205 17323 8263 17329
rect 8205 17289 8217 17323
rect 8251 17320 8263 17323
rect 8294 17320 8300 17332
rect 8251 17292 8300 17320
rect 8251 17289 8263 17292
rect 8205 17283 8263 17289
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 8665 17323 8723 17329
rect 8665 17289 8677 17323
rect 8711 17320 8723 17323
rect 8846 17320 8852 17332
rect 8711 17292 8852 17320
rect 8711 17289 8723 17292
rect 8665 17283 8723 17289
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 9122 17280 9128 17332
rect 9180 17320 9186 17332
rect 9401 17323 9459 17329
rect 9401 17320 9413 17323
rect 9180 17292 9413 17320
rect 9180 17280 9186 17292
rect 9401 17289 9413 17292
rect 9447 17289 9459 17323
rect 9401 17283 9459 17289
rect 934 17212 940 17264
rect 992 17252 998 17264
rect 992 17224 2268 17252
rect 992 17212 998 17224
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 2240 17193 2268 17224
rect 2498 17212 2504 17264
rect 2556 17252 2562 17264
rect 2685 17255 2743 17261
rect 2685 17252 2697 17255
rect 2556 17224 2697 17252
rect 2556 17212 2562 17224
rect 2685 17221 2697 17224
rect 2731 17252 2743 17255
rect 7558 17252 7564 17264
rect 2731 17224 7564 17252
rect 2731 17221 2743 17224
rect 2685 17215 2743 17221
rect 7558 17212 7564 17224
rect 7616 17212 7622 17264
rect 8018 17212 8024 17264
rect 8076 17252 8082 17264
rect 10873 17255 10931 17261
rect 10873 17252 10885 17255
rect 8076 17224 10885 17252
rect 8076 17212 8082 17224
rect 10873 17221 10885 17224
rect 10919 17221 10931 17255
rect 10873 17215 10931 17221
rect 2225 17187 2283 17193
rect 2225 17153 2237 17187
rect 2271 17153 2283 17187
rect 2225 17147 2283 17153
rect 4430 17144 4436 17196
rect 4488 17184 4494 17196
rect 4801 17187 4859 17193
rect 4801 17184 4813 17187
rect 4488 17156 4813 17184
rect 4488 17144 4494 17156
rect 4801 17153 4813 17156
rect 4847 17184 4859 17187
rect 7926 17184 7932 17196
rect 4847 17156 7932 17184
rect 4847 17153 4859 17156
rect 4801 17147 4859 17153
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 8502 17156 9781 17184
rect 8502 17128 8530 17156
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 1489 17119 1547 17125
rect 1489 17085 1501 17119
rect 1535 17085 1547 17119
rect 1489 17079 1547 17085
rect 1504 17048 1532 17079
rect 1578 17076 1584 17128
rect 1636 17116 1642 17128
rect 1946 17116 1952 17128
rect 1636 17088 1952 17116
rect 1636 17076 1642 17088
rect 1946 17076 1952 17088
rect 2004 17116 2010 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 2004 17088 2053 17116
rect 2004 17076 2010 17088
rect 2041 17085 2053 17088
rect 2087 17116 2099 17119
rect 2777 17119 2835 17125
rect 2777 17116 2789 17119
rect 2087 17088 2789 17116
rect 2087 17085 2099 17088
rect 2041 17079 2099 17085
rect 2777 17085 2789 17088
rect 2823 17085 2835 17119
rect 2777 17079 2835 17085
rect 4893 17119 4951 17125
rect 4893 17085 4905 17119
rect 4939 17085 4951 17119
rect 5258 17116 5264 17128
rect 5219 17088 5264 17116
rect 4893 17079 4951 17085
rect 2498 17048 2504 17060
rect 1504 17020 2504 17048
rect 2498 17008 2504 17020
rect 2556 17008 2562 17060
rect 4908 17048 4936 17079
rect 5258 17076 5264 17088
rect 5316 17076 5322 17128
rect 5721 17119 5779 17125
rect 5721 17085 5733 17119
rect 5767 17116 5779 17119
rect 6917 17119 6975 17125
rect 6917 17116 6929 17119
rect 5767 17088 6316 17116
rect 5767 17085 5779 17088
rect 5721 17079 5779 17085
rect 4908 17020 5856 17048
rect 5828 16992 5856 17020
rect 6288 16992 6316 17088
rect 6656 17088 6929 17116
rect 6656 16992 6684 17088
rect 6917 17085 6929 17088
rect 6963 17085 6975 17119
rect 6917 17079 6975 17085
rect 7285 17119 7343 17125
rect 7285 17085 7297 17119
rect 7331 17085 7343 17119
rect 7285 17079 7343 17085
rect 7300 17048 7328 17079
rect 7466 17076 7472 17128
rect 7524 17116 7530 17128
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7524 17088 8033 17116
rect 7524 17076 7530 17088
rect 8021 17085 8033 17088
rect 8067 17116 8079 17119
rect 8386 17116 8392 17128
rect 8067 17088 8392 17116
rect 8067 17085 8079 17088
rect 8021 17079 8079 17085
rect 8386 17076 8392 17088
rect 8444 17076 8450 17128
rect 8478 17076 8484 17128
rect 8536 17116 8542 17128
rect 8536 17088 8581 17116
rect 8536 17076 8542 17088
rect 8662 17076 8668 17128
rect 8720 17116 8726 17128
rect 9033 17119 9091 17125
rect 9033 17116 9045 17119
rect 8720 17088 9045 17116
rect 8720 17076 8726 17088
rect 9033 17085 9045 17088
rect 9079 17085 9091 17119
rect 9033 17079 9091 17085
rect 9217 17119 9275 17125
rect 9217 17085 9229 17119
rect 9263 17116 9275 17119
rect 10689 17119 10747 17125
rect 9263 17088 10088 17116
rect 9263 17085 9275 17088
rect 9217 17079 9275 17085
rect 8938 17048 8944 17060
rect 7300 17020 8944 17048
rect 8938 17008 8944 17020
rect 8996 17008 9002 17060
rect 3881 16983 3939 16989
rect 3881 16949 3893 16983
rect 3927 16980 3939 16983
rect 3970 16980 3976 16992
rect 3927 16952 3976 16980
rect 3927 16949 3939 16952
rect 3881 16943 3939 16949
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 4982 16940 4988 16992
rect 5040 16980 5046 16992
rect 5445 16983 5503 16989
rect 5445 16980 5457 16983
rect 5040 16952 5457 16980
rect 5040 16940 5046 16952
rect 5445 16949 5457 16952
rect 5491 16949 5503 16983
rect 5445 16943 5503 16949
rect 5810 16940 5816 16992
rect 5868 16980 5874 16992
rect 6089 16983 6147 16989
rect 6089 16980 6101 16983
rect 5868 16952 6101 16980
rect 5868 16940 5874 16952
rect 6089 16949 6101 16952
rect 6135 16949 6147 16983
rect 6089 16943 6147 16949
rect 6270 16940 6276 16992
rect 6328 16980 6334 16992
rect 6457 16983 6515 16989
rect 6457 16980 6469 16983
rect 6328 16952 6469 16980
rect 6328 16940 6334 16952
rect 6457 16949 6469 16952
rect 6503 16949 6515 16983
rect 6638 16980 6644 16992
rect 6599 16952 6644 16980
rect 6457 16943 6515 16949
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 7742 16940 7748 16992
rect 7800 16980 7806 16992
rect 7929 16983 7987 16989
rect 7929 16980 7941 16983
rect 7800 16952 7941 16980
rect 7800 16940 7806 16952
rect 7929 16949 7941 16952
rect 7975 16980 7987 16983
rect 9398 16980 9404 16992
rect 7975 16952 9404 16980
rect 7975 16949 7987 16952
rect 7929 16943 7987 16949
rect 9398 16940 9404 16952
rect 9456 16940 9462 16992
rect 10060 16989 10088 17088
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 10735 17088 11192 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 10045 16983 10103 16989
rect 10045 16949 10057 16983
rect 10091 16980 10103 16983
rect 10318 16980 10324 16992
rect 10091 16952 10324 16980
rect 10091 16949 10103 16952
rect 10045 16943 10103 16949
rect 10318 16940 10324 16952
rect 10376 16940 10382 16992
rect 11164 16989 11192 17088
rect 14274 17076 14280 17128
rect 14332 17116 14338 17128
rect 14553 17119 14611 17125
rect 14553 17116 14565 17119
rect 14332 17088 14565 17116
rect 14332 17076 14338 17088
rect 14553 17085 14565 17088
rect 14599 17116 14611 17119
rect 15105 17119 15163 17125
rect 15105 17116 15117 17119
rect 14599 17088 15117 17116
rect 14599 17085 14611 17088
rect 14553 17079 14611 17085
rect 15105 17085 15117 17088
rect 15151 17085 15163 17119
rect 15105 17079 15163 17085
rect 14826 17048 14832 17060
rect 14787 17020 14832 17048
rect 14826 17008 14832 17020
rect 14884 17008 14890 17060
rect 11149 16983 11207 16989
rect 11149 16949 11161 16983
rect 11195 16980 11207 16983
rect 11698 16980 11704 16992
rect 11195 16952 11704 16980
rect 11195 16949 11207 16952
rect 11149 16943 11207 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 1104 16890 16008 16912
rect 1104 16838 5979 16890
rect 6031 16838 6043 16890
rect 6095 16838 6107 16890
rect 6159 16838 6171 16890
rect 6223 16838 10976 16890
rect 11028 16838 11040 16890
rect 11092 16838 11104 16890
rect 11156 16838 11168 16890
rect 11220 16838 16008 16890
rect 1104 16816 16008 16838
rect 2498 16776 2504 16788
rect 2459 16748 2504 16776
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 3237 16779 3295 16785
rect 3237 16776 3249 16779
rect 2832 16748 3249 16776
rect 2832 16736 2838 16748
rect 3237 16745 3249 16748
rect 3283 16745 3295 16779
rect 3237 16739 3295 16745
rect 3786 16736 3792 16788
rect 3844 16776 3850 16788
rect 4249 16779 4307 16785
rect 4249 16776 4261 16779
rect 3844 16748 4261 16776
rect 3844 16736 3850 16748
rect 4249 16745 4261 16748
rect 4295 16745 4307 16779
rect 4249 16739 4307 16745
rect 4338 16736 4344 16788
rect 4396 16776 4402 16788
rect 4985 16779 5043 16785
rect 4985 16776 4997 16779
rect 4396 16748 4997 16776
rect 4396 16736 4402 16748
rect 4985 16745 4997 16748
rect 5031 16745 5043 16779
rect 4985 16739 5043 16745
rect 6546 16736 6552 16788
rect 6604 16776 6610 16788
rect 7377 16779 7435 16785
rect 7377 16776 7389 16779
rect 6604 16748 7389 16776
rect 6604 16736 6610 16748
rect 7377 16745 7389 16748
rect 7423 16745 7435 16779
rect 7377 16739 7435 16745
rect 7650 16736 7656 16788
rect 7708 16776 7714 16788
rect 8205 16779 8263 16785
rect 8205 16776 8217 16779
rect 7708 16748 8217 16776
rect 7708 16736 7714 16748
rect 8205 16745 8217 16748
rect 8251 16745 8263 16779
rect 8205 16739 8263 16745
rect 10134 16736 10140 16788
rect 10192 16776 10198 16788
rect 13081 16779 13139 16785
rect 13081 16776 13093 16779
rect 10192 16748 13093 16776
rect 10192 16736 10198 16748
rect 13081 16745 13093 16748
rect 13127 16745 13139 16779
rect 13081 16739 13139 16745
rect 2038 16668 2044 16720
rect 2096 16708 2102 16720
rect 2133 16711 2191 16717
rect 2133 16708 2145 16711
rect 2096 16680 2145 16708
rect 2096 16668 2102 16680
rect 2133 16677 2145 16680
rect 2179 16677 2191 16711
rect 2133 16671 2191 16677
rect 1857 16643 1915 16649
rect 1857 16609 1869 16643
rect 1903 16640 1915 16643
rect 2516 16640 2544 16736
rect 5534 16668 5540 16720
rect 5592 16708 5598 16720
rect 9309 16711 9367 16717
rect 9309 16708 9321 16711
rect 5592 16680 7880 16708
rect 5592 16668 5598 16680
rect 1903 16612 2544 16640
rect 3053 16643 3111 16649
rect 1903 16609 1915 16612
rect 1857 16603 1915 16609
rect 3053 16609 3065 16643
rect 3099 16609 3111 16643
rect 3053 16603 3111 16609
rect 3068 16572 3096 16603
rect 3418 16600 3424 16652
rect 3476 16640 3482 16652
rect 4065 16643 4123 16649
rect 3476 16612 3521 16640
rect 3476 16600 3482 16612
rect 4065 16609 4077 16643
rect 4111 16609 4123 16643
rect 4430 16640 4436 16652
rect 4391 16612 4436 16640
rect 4065 16603 4123 16609
rect 3786 16572 3792 16584
rect 3068 16544 3792 16572
rect 3786 16532 3792 16544
rect 3844 16532 3850 16584
rect 4080 16572 4108 16603
rect 4430 16600 4436 16612
rect 4488 16600 4494 16652
rect 4798 16640 4804 16652
rect 4759 16612 4804 16640
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 5620 16643 5678 16649
rect 5620 16609 5632 16643
rect 5666 16640 5678 16643
rect 5994 16640 6000 16652
rect 5666 16612 6000 16640
rect 5666 16609 5678 16612
rect 5620 16603 5678 16609
rect 5994 16600 6000 16612
rect 6052 16600 6058 16652
rect 6822 16640 6828 16652
rect 6783 16612 6828 16640
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16640 7251 16643
rect 7558 16640 7564 16652
rect 7239 16612 7564 16640
rect 7239 16609 7251 16612
rect 7193 16603 7251 16609
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 7653 16643 7711 16649
rect 7653 16609 7665 16643
rect 7699 16640 7711 16643
rect 7699 16612 7788 16640
rect 7699 16609 7711 16612
rect 7653 16603 7711 16609
rect 7760 16584 7788 16612
rect 5350 16572 5356 16584
rect 4080 16544 5028 16572
rect 5311 16544 5356 16572
rect 3142 16464 3148 16516
rect 3200 16504 3206 16516
rect 3605 16507 3663 16513
rect 3605 16504 3617 16507
rect 3200 16476 3617 16504
rect 3200 16464 3206 16476
rect 3605 16473 3617 16476
rect 3651 16473 3663 16507
rect 3605 16467 3663 16473
rect 3878 16464 3884 16516
rect 3936 16504 3942 16516
rect 4617 16507 4675 16513
rect 4617 16504 4629 16507
rect 3936 16476 4629 16504
rect 3936 16464 3942 16476
rect 4617 16473 4629 16476
rect 4663 16473 4675 16507
rect 4617 16467 4675 16473
rect 5000 16448 5028 16544
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 7742 16532 7748 16584
rect 7800 16532 7806 16584
rect 6362 16464 6368 16516
rect 6420 16504 6426 16516
rect 7852 16513 7880 16680
rect 8128 16680 9321 16708
rect 8128 16652 8156 16680
rect 9309 16677 9321 16680
rect 9355 16677 9367 16711
rect 9309 16671 9367 16677
rect 9674 16668 9680 16720
rect 9732 16708 9738 16720
rect 9732 16680 10088 16708
rect 9732 16668 9738 16680
rect 8021 16643 8079 16649
rect 8021 16609 8033 16643
rect 8067 16640 8079 16643
rect 8110 16640 8116 16652
rect 8067 16612 8116 16640
rect 8067 16609 8079 16612
rect 8021 16603 8079 16609
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 8849 16643 8907 16649
rect 8849 16609 8861 16643
rect 8895 16640 8907 16643
rect 9490 16640 9496 16652
rect 8895 16612 9496 16640
rect 8895 16609 8907 16612
rect 8849 16603 8907 16609
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 9950 16649 9956 16652
rect 9944 16640 9956 16649
rect 9600 16612 9956 16640
rect 8938 16572 8944 16584
rect 8899 16544 8944 16572
rect 8938 16532 8944 16544
rect 8996 16532 9002 16584
rect 9125 16575 9183 16581
rect 9125 16541 9137 16575
rect 9171 16572 9183 16575
rect 9600 16572 9628 16612
rect 9944 16603 9956 16612
rect 9950 16600 9956 16603
rect 10008 16600 10014 16652
rect 10060 16640 10088 16680
rect 10226 16668 10232 16720
rect 10284 16708 10290 16720
rect 11146 16708 11152 16720
rect 10284 16680 11152 16708
rect 10284 16668 10290 16680
rect 11146 16668 11152 16680
rect 11204 16668 11210 16720
rect 11606 16668 11612 16720
rect 11664 16717 11670 16720
rect 11664 16711 11728 16717
rect 11664 16677 11682 16711
rect 11716 16677 11728 16711
rect 14921 16711 14979 16717
rect 14921 16708 14933 16711
rect 11664 16671 11728 16677
rect 14384 16680 14933 16708
rect 11664 16668 11670 16671
rect 11425 16643 11483 16649
rect 11425 16640 11437 16643
rect 10060 16612 11437 16640
rect 11425 16609 11437 16612
rect 11471 16640 11483 16643
rect 12066 16640 12072 16652
rect 11471 16612 12072 16640
rect 11471 16609 11483 16612
rect 11425 16603 11483 16609
rect 12066 16600 12072 16612
rect 12124 16600 12130 16652
rect 12897 16643 12955 16649
rect 12897 16609 12909 16643
rect 12943 16640 12955 16643
rect 13262 16640 13268 16652
rect 12943 16612 13268 16640
rect 12943 16609 12955 16612
rect 12897 16603 12955 16609
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 14090 16600 14096 16652
rect 14148 16640 14154 16652
rect 14384 16649 14412 16680
rect 14921 16677 14933 16680
rect 14967 16677 14979 16711
rect 14921 16671 14979 16677
rect 14369 16643 14427 16649
rect 14369 16640 14381 16643
rect 14148 16612 14381 16640
rect 14148 16600 14154 16612
rect 14369 16609 14381 16612
rect 14415 16609 14427 16643
rect 14642 16640 14648 16652
rect 14603 16612 14648 16640
rect 14369 16603 14427 16609
rect 14642 16600 14648 16612
rect 14700 16600 14706 16652
rect 9171 16544 9628 16572
rect 9171 16541 9183 16544
rect 9125 16535 9183 16541
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 11146 16572 11152 16584
rect 9732 16544 9777 16572
rect 11107 16544 11152 16572
rect 9732 16532 9738 16544
rect 11146 16532 11152 16544
rect 11204 16532 11210 16584
rect 7009 16507 7067 16513
rect 7009 16504 7021 16507
rect 6420 16476 7021 16504
rect 6420 16464 6426 16476
rect 7009 16473 7021 16476
rect 7055 16473 7067 16507
rect 7009 16467 7067 16473
rect 7837 16507 7895 16513
rect 7837 16473 7849 16507
rect 7883 16473 7895 16507
rect 7837 16467 7895 16473
rect 11057 16507 11115 16513
rect 11057 16473 11069 16507
rect 11103 16504 11115 16507
rect 11422 16504 11428 16516
rect 11103 16476 11428 16504
rect 11103 16473 11115 16476
rect 11057 16467 11115 16473
rect 11422 16464 11428 16476
rect 11480 16464 11486 16516
rect 12805 16507 12863 16513
rect 12805 16473 12817 16507
rect 12851 16504 12863 16507
rect 12986 16504 12992 16516
rect 12851 16476 12992 16504
rect 12851 16473 12863 16476
rect 12805 16467 12863 16473
rect 12986 16464 12992 16476
rect 13044 16464 13050 16516
rect 4982 16396 4988 16448
rect 5040 16436 5046 16448
rect 5169 16439 5227 16445
rect 5169 16436 5181 16439
rect 5040 16408 5181 16436
rect 5040 16396 5046 16408
rect 5169 16405 5181 16408
rect 5215 16405 5227 16439
rect 6730 16436 6736 16448
rect 6691 16408 6736 16436
rect 5169 16399 5227 16405
rect 6730 16396 6736 16408
rect 6788 16396 6794 16448
rect 8294 16396 8300 16448
rect 8352 16436 8358 16448
rect 8481 16439 8539 16445
rect 8481 16436 8493 16439
rect 8352 16408 8493 16436
rect 8352 16396 8358 16408
rect 8481 16405 8493 16408
rect 8527 16405 8539 16439
rect 8481 16399 8539 16405
rect 1104 16346 16008 16368
rect 1104 16294 3480 16346
rect 3532 16294 3544 16346
rect 3596 16294 3608 16346
rect 3660 16294 3672 16346
rect 3724 16294 8478 16346
rect 8530 16294 8542 16346
rect 8594 16294 8606 16346
rect 8658 16294 8670 16346
rect 8722 16294 13475 16346
rect 13527 16294 13539 16346
rect 13591 16294 13603 16346
rect 13655 16294 13667 16346
rect 13719 16294 16008 16346
rect 1104 16272 16008 16294
rect 1486 16192 1492 16244
rect 1544 16232 1550 16244
rect 1544 16204 5580 16232
rect 1544 16192 1550 16204
rect 5552 16164 5580 16204
rect 5626 16192 5632 16244
rect 5684 16232 5690 16244
rect 5994 16232 6000 16244
rect 5684 16204 6000 16232
rect 5684 16192 5690 16204
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 6641 16235 6699 16241
rect 6641 16201 6653 16235
rect 6687 16232 6699 16235
rect 7742 16232 7748 16244
rect 6687 16204 7748 16232
rect 6687 16201 6699 16204
rect 6641 16195 6699 16201
rect 7742 16192 7748 16204
rect 7800 16232 7806 16244
rect 8846 16232 8852 16244
rect 7800 16204 8852 16232
rect 7800 16192 7806 16204
rect 8846 16192 8852 16204
rect 8904 16192 8910 16244
rect 9950 16192 9956 16244
rect 10008 16232 10014 16244
rect 10597 16235 10655 16241
rect 10597 16232 10609 16235
rect 10008 16204 10609 16232
rect 10008 16192 10014 16204
rect 10597 16201 10609 16204
rect 10643 16201 10655 16235
rect 10597 16195 10655 16201
rect 10870 16192 10876 16244
rect 10928 16232 10934 16244
rect 15102 16232 15108 16244
rect 10928 16204 15108 16232
rect 10928 16192 10934 16204
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 5552 16136 7512 16164
rect 198 16056 204 16108
rect 256 16096 262 16108
rect 1765 16099 1823 16105
rect 1765 16096 1777 16099
rect 256 16068 1777 16096
rect 256 16056 262 16068
rect 1765 16065 1777 16068
rect 1811 16065 1823 16099
rect 7374 16096 7380 16108
rect 7335 16068 7380 16096
rect 1765 16059 1823 16065
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 7484 16096 7512 16136
rect 10226 16124 10232 16176
rect 10284 16164 10290 16176
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 10284 16136 11805 16164
rect 10284 16124 10290 16136
rect 11793 16133 11805 16136
rect 11839 16164 11851 16167
rect 12250 16164 12256 16176
rect 11839 16136 12256 16164
rect 11839 16133 11851 16136
rect 11793 16127 11851 16133
rect 12250 16124 12256 16136
rect 12308 16124 12314 16176
rect 7484 16068 7880 16096
rect 1581 16031 1639 16037
rect 1581 15997 1593 16031
rect 1627 16028 1639 16031
rect 1627 16000 2268 16028
rect 1627 15997 1639 16000
rect 1581 15991 1639 15997
rect 2240 15901 2268 16000
rect 2682 15988 2688 16040
rect 2740 16028 2746 16040
rect 3145 16031 3203 16037
rect 3145 16028 3157 16031
rect 2740 16000 3157 16028
rect 2740 15988 2746 16000
rect 3145 15997 3157 16000
rect 3191 16028 3203 16031
rect 4614 16028 4620 16040
rect 3191 16000 4620 16028
rect 3191 15997 3203 16000
rect 3145 15991 3203 15997
rect 4614 15988 4620 16000
rect 4672 16028 4678 16040
rect 5350 16028 5356 16040
rect 4672 16000 5356 16028
rect 4672 15988 4678 16000
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 7742 16028 7748 16040
rect 7703 16000 7748 16028
rect 7742 15988 7748 16000
rect 7800 15988 7806 16040
rect 7852 16028 7880 16068
rect 10778 16056 10784 16108
rect 10836 16096 10842 16108
rect 10873 16099 10931 16105
rect 10873 16096 10885 16099
rect 10836 16068 10885 16096
rect 10836 16056 10842 16068
rect 10873 16065 10885 16068
rect 10919 16096 10931 16099
rect 11425 16099 11483 16105
rect 11425 16096 11437 16099
rect 10919 16068 11437 16096
rect 10919 16065 10931 16068
rect 10873 16059 10931 16065
rect 11425 16065 11437 16068
rect 11471 16065 11483 16099
rect 11606 16096 11612 16108
rect 11567 16068 11612 16096
rect 11425 16059 11483 16065
rect 11606 16056 11612 16068
rect 11664 16056 11670 16108
rect 12986 16096 12992 16108
rect 12947 16068 12992 16096
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 8294 16028 8300 16040
rect 7852 16000 8300 16028
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 9217 16031 9275 16037
rect 9217 15997 9229 16031
rect 9263 16028 9275 16031
rect 9766 16028 9772 16040
rect 9263 16000 9772 16028
rect 9263 15997 9275 16000
rect 9217 15991 9275 15997
rect 9766 15988 9772 16000
rect 9824 15988 9830 16040
rect 11146 16028 11152 16040
rect 10879 16000 11152 16028
rect 3326 15920 3332 15972
rect 3384 15969 3390 15972
rect 3384 15963 3448 15969
rect 3384 15929 3402 15963
rect 3436 15929 3448 15963
rect 4862 15963 4920 15969
rect 4862 15960 4874 15963
rect 3384 15923 3448 15929
rect 4724 15932 4874 15960
rect 3384 15920 3390 15923
rect 4724 15904 4752 15932
rect 4862 15929 4874 15932
rect 4908 15929 4920 15963
rect 4862 15923 4920 15929
rect 6273 15963 6331 15969
rect 6273 15929 6285 15963
rect 6319 15960 6331 15963
rect 8012 15963 8070 15969
rect 6319 15932 7328 15960
rect 6319 15929 6331 15932
rect 6273 15923 6331 15929
rect 7300 15904 7328 15932
rect 8012 15929 8024 15963
rect 8058 15960 8070 15963
rect 9030 15960 9036 15972
rect 8058 15932 9036 15960
rect 8058 15929 8070 15932
rect 8012 15923 8070 15929
rect 9030 15920 9036 15932
rect 9088 15920 9094 15972
rect 9484 15963 9542 15969
rect 9484 15960 9496 15963
rect 9140 15932 9496 15960
rect 2225 15895 2283 15901
rect 2225 15861 2237 15895
rect 2271 15892 2283 15895
rect 2314 15892 2320 15904
rect 2271 15864 2320 15892
rect 2271 15861 2283 15864
rect 2225 15855 2283 15861
rect 2314 15852 2320 15864
rect 2372 15852 2378 15904
rect 4525 15895 4583 15901
rect 4525 15861 4537 15895
rect 4571 15892 4583 15895
rect 4706 15892 4712 15904
rect 4571 15864 4712 15892
rect 4571 15861 4583 15864
rect 4525 15855 4583 15861
rect 4706 15852 4712 15864
rect 4764 15852 4770 15904
rect 6454 15892 6460 15904
rect 6415 15864 6460 15892
rect 6454 15852 6460 15864
rect 6512 15852 6518 15904
rect 6822 15892 6828 15904
rect 6783 15864 6828 15892
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7190 15892 7196 15904
rect 7151 15864 7196 15892
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 7282 15852 7288 15904
rect 7340 15892 7346 15904
rect 9140 15901 9168 15932
rect 9484 15929 9496 15932
rect 9530 15960 9542 15963
rect 9950 15960 9956 15972
rect 9530 15932 9956 15960
rect 9530 15929 9542 15932
rect 9484 15923 9542 15929
rect 9950 15920 9956 15932
rect 10008 15920 10014 15972
rect 9125 15895 9183 15901
rect 7340 15864 7385 15892
rect 7340 15852 7346 15864
rect 9125 15861 9137 15895
rect 9171 15861 9183 15895
rect 9125 15855 9183 15861
rect 9582 15852 9588 15904
rect 9640 15892 9646 15904
rect 10134 15892 10140 15904
rect 9640 15864 10140 15892
rect 9640 15852 9646 15864
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 10879 15892 10907 16000
rect 11146 15988 11152 16000
rect 11204 16028 11210 16040
rect 11333 16031 11391 16037
rect 11333 16028 11345 16031
rect 11204 16000 11345 16028
rect 11204 15988 11210 16000
rect 11333 15997 11345 16000
rect 11379 15997 11391 16031
rect 11333 15991 11391 15997
rect 11882 15988 11888 16040
rect 11940 16028 11946 16040
rect 13354 16028 13360 16040
rect 11940 16000 13360 16028
rect 11940 15988 11946 16000
rect 13354 15988 13360 16000
rect 13412 15988 13418 16040
rect 12897 15963 12955 15969
rect 12897 15960 12909 15963
rect 10980 15932 12909 15960
rect 10980 15901 11008 15932
rect 12897 15929 12909 15932
rect 12943 15929 12955 15963
rect 12897 15923 12955 15929
rect 10560 15864 10907 15892
rect 10965 15895 11023 15901
rect 10560 15852 10566 15864
rect 10965 15861 10977 15895
rect 11011 15861 11023 15895
rect 10965 15855 11023 15861
rect 12437 15895 12495 15901
rect 12437 15861 12449 15895
rect 12483 15892 12495 15895
rect 12618 15892 12624 15904
rect 12483 15864 12624 15892
rect 12483 15861 12495 15864
rect 12437 15855 12495 15861
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 12802 15892 12808 15904
rect 12763 15864 12808 15892
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 1104 15802 16008 15824
rect 1104 15750 5979 15802
rect 6031 15750 6043 15802
rect 6095 15750 6107 15802
rect 6159 15750 6171 15802
rect 6223 15750 10976 15802
rect 11028 15750 11040 15802
rect 11092 15750 11104 15802
rect 11156 15750 11168 15802
rect 11220 15750 16008 15802
rect 1104 15728 16008 15750
rect 2406 15648 2412 15700
rect 2464 15688 2470 15700
rect 2777 15691 2835 15697
rect 2777 15688 2789 15691
rect 2464 15660 2789 15688
rect 2464 15648 2470 15660
rect 2777 15657 2789 15660
rect 2823 15657 2835 15691
rect 5905 15691 5963 15697
rect 2777 15651 2835 15657
rect 4172 15660 5764 15688
rect 4172 15620 4200 15660
rect 3804 15592 4200 15620
rect 1486 15552 1492 15564
rect 1447 15524 1492 15552
rect 1486 15512 1492 15524
rect 1544 15512 1550 15564
rect 2593 15555 2651 15561
rect 2593 15521 2605 15555
rect 2639 15552 2651 15555
rect 2958 15552 2964 15564
rect 2639 15524 2964 15552
rect 2639 15521 2651 15524
rect 2593 15515 2651 15521
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 3513 15555 3571 15561
rect 3513 15521 3525 15555
rect 3559 15521 3571 15555
rect 3513 15515 3571 15521
rect 1670 15484 1676 15496
rect 1631 15456 1676 15484
rect 1670 15444 1676 15456
rect 1728 15444 1734 15496
rect 2866 15376 2872 15428
rect 2924 15416 2930 15428
rect 3145 15419 3203 15425
rect 3145 15416 3157 15419
rect 2924 15388 3157 15416
rect 2924 15376 2930 15388
rect 3145 15385 3157 15388
rect 3191 15385 3203 15419
rect 3145 15379 3203 15385
rect 3528 15348 3556 15515
rect 3804 15493 3832 15592
rect 4798 15580 4804 15632
rect 4856 15620 4862 15632
rect 5169 15623 5227 15629
rect 5169 15620 5181 15623
rect 4856 15592 5181 15620
rect 4856 15580 4862 15592
rect 5169 15589 5181 15592
rect 5215 15620 5227 15623
rect 5258 15620 5264 15632
rect 5215 15592 5264 15620
rect 5215 15589 5227 15592
rect 5169 15583 5227 15589
rect 5258 15580 5264 15592
rect 5316 15580 5322 15632
rect 5736 15620 5764 15660
rect 5905 15657 5917 15691
rect 5951 15688 5963 15691
rect 6454 15688 6460 15700
rect 5951 15660 6460 15688
rect 5951 15657 5963 15660
rect 5905 15651 5963 15657
rect 6454 15648 6460 15660
rect 6512 15648 6518 15700
rect 6546 15648 6552 15700
rect 6604 15688 6610 15700
rect 8665 15691 8723 15697
rect 6604 15660 8616 15688
rect 6604 15648 6610 15660
rect 6730 15629 6736 15632
rect 6702 15623 6736 15629
rect 6702 15620 6714 15623
rect 5736 15592 6714 15620
rect 6702 15589 6714 15592
rect 6788 15620 6794 15632
rect 6788 15592 6850 15620
rect 6702 15583 6736 15589
rect 6730 15580 6736 15583
rect 6788 15580 6794 15592
rect 7190 15580 7196 15632
rect 7248 15620 7254 15632
rect 8113 15623 8171 15629
rect 8113 15620 8125 15623
rect 7248 15592 8125 15620
rect 7248 15580 7254 15592
rect 8113 15589 8125 15592
rect 8159 15620 8171 15623
rect 8202 15620 8208 15632
rect 8159 15592 8208 15620
rect 8159 15589 8171 15592
rect 8113 15583 8171 15589
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 8588 15620 8616 15660
rect 8665 15657 8677 15691
rect 8711 15688 8723 15691
rect 8938 15688 8944 15700
rect 8711 15660 8944 15688
rect 8711 15657 8723 15660
rect 8665 15651 8723 15657
rect 8938 15648 8944 15660
rect 8996 15648 9002 15700
rect 9033 15691 9091 15697
rect 9033 15657 9045 15691
rect 9079 15688 9091 15691
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 9079 15660 9689 15688
rect 9079 15657 9091 15660
rect 9033 15651 9091 15657
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 10137 15691 10195 15697
rect 10137 15688 10149 15691
rect 9677 15651 9735 15657
rect 9784 15660 10149 15688
rect 8588 15592 9352 15620
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 4982 15552 4988 15564
rect 4479 15524 4988 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 4982 15512 4988 15524
rect 5040 15512 5046 15564
rect 5813 15555 5871 15561
rect 5813 15521 5825 15555
rect 5859 15552 5871 15555
rect 5902 15552 5908 15564
rect 5859 15524 5908 15552
rect 5859 15521 5871 15524
rect 5813 15515 5871 15521
rect 5902 15512 5908 15524
rect 5960 15512 5966 15564
rect 7282 15552 7288 15564
rect 6104 15524 7288 15552
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15453 3663 15487
rect 3605 15447 3663 15453
rect 3789 15487 3847 15493
rect 3789 15453 3801 15487
rect 3835 15453 3847 15487
rect 4338 15484 4344 15496
rect 3789 15447 3847 15453
rect 3988 15456 4344 15484
rect 3620 15416 3648 15447
rect 3988 15416 4016 15456
rect 4338 15444 4344 15456
rect 4396 15444 4402 15496
rect 4522 15484 4528 15496
rect 4483 15456 4528 15484
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 4706 15484 4712 15496
rect 4619 15456 4712 15484
rect 4706 15444 4712 15456
rect 4764 15484 4770 15496
rect 6104 15493 6132 15524
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 8573 15555 8631 15561
rect 8573 15521 8585 15555
rect 8619 15552 8631 15555
rect 9214 15552 9220 15564
rect 8619 15524 9220 15552
rect 8619 15521 8631 15524
rect 8573 15515 8631 15521
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 9324 15552 9352 15592
rect 9582 15580 9588 15632
rect 9640 15620 9646 15632
rect 9784 15620 9812 15660
rect 10137 15657 10149 15660
rect 10183 15688 10195 15691
rect 10410 15688 10416 15700
rect 10183 15660 10416 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 10410 15648 10416 15660
rect 10468 15688 10474 15700
rect 10686 15688 10692 15700
rect 10468 15660 10692 15688
rect 10468 15648 10474 15660
rect 10686 15648 10692 15660
rect 10744 15648 10750 15700
rect 10965 15691 11023 15697
rect 10965 15657 10977 15691
rect 11011 15688 11023 15691
rect 12802 15688 12808 15700
rect 11011 15660 12808 15688
rect 11011 15657 11023 15660
rect 10965 15651 11023 15657
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 10226 15620 10232 15632
rect 9640 15592 9812 15620
rect 9883 15592 10232 15620
rect 9640 15580 9646 15592
rect 9883 15552 9911 15592
rect 10226 15580 10232 15592
rect 10284 15580 10290 15632
rect 10594 15580 10600 15632
rect 10652 15620 10658 15632
rect 11790 15620 11796 15632
rect 10652 15592 11796 15620
rect 10652 15580 10658 15592
rect 11790 15580 11796 15592
rect 11848 15580 11854 15632
rect 12621 15623 12679 15629
rect 12621 15620 12633 15623
rect 11900 15592 12633 15620
rect 10042 15552 10048 15564
rect 9324 15524 9911 15552
rect 9955 15524 10048 15552
rect 10042 15512 10048 15524
rect 10100 15552 10106 15564
rect 11330 15552 11336 15564
rect 10100 15524 10640 15552
rect 11291 15524 11336 15552
rect 10100 15512 10106 15524
rect 6089 15487 6147 15493
rect 6089 15484 6101 15487
rect 4764 15456 6101 15484
rect 4764 15444 4770 15456
rect 6089 15453 6101 15456
rect 6135 15453 6147 15487
rect 6089 15447 6147 15453
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15453 6515 15487
rect 6457 15447 6515 15453
rect 3620 15388 4016 15416
rect 4065 15419 4123 15425
rect 4065 15385 4077 15419
rect 4111 15416 4123 15419
rect 5350 15416 5356 15428
rect 4111 15388 5356 15416
rect 4111 15385 4123 15388
rect 4065 15379 4123 15385
rect 5350 15376 5356 15388
rect 5408 15376 5414 15428
rect 5534 15376 5540 15428
rect 5592 15416 5598 15428
rect 6472 15416 6500 15447
rect 7742 15444 7748 15496
rect 7800 15484 7806 15496
rect 9122 15484 9128 15496
rect 7800 15456 8432 15484
rect 9083 15456 9128 15484
rect 7800 15444 7806 15456
rect 7926 15416 7932 15428
rect 5592 15388 6500 15416
rect 7392 15388 7932 15416
rect 5592 15376 5598 15388
rect 4798 15348 4804 15360
rect 3528 15320 4804 15348
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 4982 15348 4988 15360
rect 4943 15320 4988 15348
rect 4982 15308 4988 15320
rect 5040 15308 5046 15360
rect 5442 15348 5448 15360
rect 5403 15320 5448 15348
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 5902 15308 5908 15360
rect 5960 15348 5966 15360
rect 6270 15348 6276 15360
rect 5960 15320 6276 15348
rect 5960 15308 5966 15320
rect 6270 15308 6276 15320
rect 6328 15308 6334 15360
rect 6362 15308 6368 15360
rect 6420 15348 6426 15360
rect 7392 15348 7420 15388
rect 7926 15376 7932 15388
rect 7984 15376 7990 15428
rect 8404 15425 8432 15456
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9309 15487 9367 15493
rect 9309 15453 9321 15487
rect 9355 15484 9367 15487
rect 9950 15484 9956 15496
rect 9355 15456 9956 15484
rect 9355 15453 9367 15456
rect 9309 15447 9367 15453
rect 9950 15444 9956 15456
rect 10008 15444 10014 15496
rect 10134 15444 10140 15496
rect 10192 15484 10198 15496
rect 10612 15493 10640 15524
rect 11330 15512 11336 15524
rect 11388 15552 11394 15564
rect 11900 15552 11928 15592
rect 12621 15589 12633 15592
rect 12667 15589 12679 15623
rect 14366 15620 14372 15632
rect 14327 15592 14372 15620
rect 12621 15583 12679 15589
rect 14366 15580 14372 15592
rect 14424 15580 14430 15632
rect 12161 15555 12219 15561
rect 12161 15552 12173 15555
rect 11388 15524 11928 15552
rect 11983 15524 12173 15552
rect 11388 15512 11394 15524
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 10192 15456 10241 15484
rect 10192 15444 10198 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 10597 15487 10655 15493
rect 10597 15453 10609 15487
rect 10643 15484 10655 15487
rect 10962 15484 10968 15496
rect 10643 15456 10968 15484
rect 10643 15453 10655 15456
rect 10597 15447 10655 15453
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11425 15487 11483 15493
rect 11425 15484 11437 15487
rect 11072 15456 11437 15484
rect 8389 15419 8447 15425
rect 8389 15385 8401 15419
rect 8435 15416 8447 15419
rect 9674 15416 9680 15428
rect 8435 15388 9680 15416
rect 8435 15385 8447 15388
rect 8389 15379 8447 15385
rect 9674 15376 9680 15388
rect 9732 15376 9738 15428
rect 10042 15376 10048 15428
rect 10100 15416 10106 15428
rect 10870 15416 10876 15428
rect 10100 15388 10876 15416
rect 10100 15376 10106 15388
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 7834 15348 7840 15360
rect 6420 15320 7420 15348
rect 7795 15320 7840 15348
rect 6420 15308 6426 15320
rect 7834 15308 7840 15320
rect 7892 15308 7898 15360
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 8996 15320 10793 15348
rect 8996 15308 9002 15320
rect 10781 15317 10793 15320
rect 10827 15348 10839 15351
rect 11072 15348 11100 15456
rect 11425 15453 11437 15456
rect 11471 15453 11483 15487
rect 11606 15484 11612 15496
rect 11519 15456 11612 15484
rect 11425 15447 11483 15453
rect 11606 15444 11612 15456
rect 11664 15444 11670 15496
rect 11790 15444 11796 15496
rect 11848 15484 11854 15496
rect 11983 15484 12011 15524
rect 12161 15521 12173 15524
rect 12207 15552 12219 15555
rect 12805 15555 12863 15561
rect 12805 15552 12817 15555
rect 12207 15524 12817 15552
rect 12207 15521 12219 15524
rect 12161 15515 12219 15521
rect 12805 15521 12817 15524
rect 12851 15552 12863 15555
rect 13170 15552 13176 15564
rect 12851 15524 13176 15552
rect 12851 15521 12863 15524
rect 12805 15515 12863 15521
rect 13170 15512 13176 15524
rect 13228 15512 13234 15564
rect 14093 15555 14151 15561
rect 14093 15521 14105 15555
rect 14139 15552 14151 15555
rect 14139 15524 14780 15552
rect 14139 15521 14151 15524
rect 14093 15515 14151 15521
rect 12250 15484 12256 15496
rect 11848 15456 12011 15484
rect 12211 15456 12256 15484
rect 11848 15444 11854 15456
rect 12250 15444 12256 15456
rect 12308 15444 12314 15496
rect 12345 15487 12403 15493
rect 12345 15453 12357 15487
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 11624 15416 11652 15444
rect 12360 15416 12388 15447
rect 11624 15388 12388 15416
rect 10827 15320 11100 15348
rect 10827 15317 10839 15320
rect 10781 15311 10839 15317
rect 11422 15308 11428 15360
rect 11480 15348 11486 15360
rect 14752 15357 14780 15524
rect 11793 15351 11851 15357
rect 11793 15348 11805 15351
rect 11480 15320 11805 15348
rect 11480 15308 11486 15320
rect 11793 15317 11805 15320
rect 11839 15317 11851 15351
rect 11793 15311 11851 15317
rect 14737 15351 14795 15357
rect 14737 15317 14749 15351
rect 14783 15348 14795 15351
rect 14918 15348 14924 15360
rect 14783 15320 14924 15348
rect 14783 15317 14795 15320
rect 14737 15311 14795 15317
rect 14918 15308 14924 15320
rect 14976 15308 14982 15360
rect 1104 15258 16008 15280
rect 1104 15206 3480 15258
rect 3532 15206 3544 15258
rect 3596 15206 3608 15258
rect 3660 15206 3672 15258
rect 3724 15206 8478 15258
rect 8530 15206 8542 15258
rect 8594 15206 8606 15258
rect 8658 15206 8670 15258
rect 8722 15206 13475 15258
rect 13527 15206 13539 15258
rect 13591 15206 13603 15258
rect 13655 15206 13667 15258
rect 13719 15206 16008 15258
rect 1104 15184 16008 15206
rect 3326 15104 3332 15156
rect 3384 15144 3390 15156
rect 3697 15147 3755 15153
rect 3697 15144 3709 15147
rect 3384 15116 3709 15144
rect 3384 15104 3390 15116
rect 3697 15113 3709 15116
rect 3743 15113 3755 15147
rect 3697 15107 3755 15113
rect 3789 15147 3847 15153
rect 3789 15113 3801 15147
rect 3835 15144 3847 15147
rect 4522 15144 4528 15156
rect 3835 15116 4528 15144
rect 3835 15113 3847 15116
rect 3789 15107 3847 15113
rect 3712 15008 3740 15107
rect 4522 15104 4528 15116
rect 4580 15104 4586 15156
rect 4798 15104 4804 15156
rect 4856 15144 4862 15156
rect 5813 15147 5871 15153
rect 5813 15144 5825 15147
rect 4856 15116 5825 15144
rect 4856 15104 4862 15116
rect 5813 15113 5825 15116
rect 5859 15113 5871 15147
rect 5813 15107 5871 15113
rect 8481 15147 8539 15153
rect 8481 15113 8493 15147
rect 8527 15144 8539 15147
rect 9122 15144 9128 15156
rect 8527 15116 9128 15144
rect 8527 15113 8539 15116
rect 8481 15107 8539 15113
rect 9122 15104 9128 15116
rect 9180 15104 9186 15156
rect 9490 15104 9496 15156
rect 9548 15144 9554 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 9548 15116 10149 15144
rect 9548 15104 9554 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 13170 15144 13176 15156
rect 10137 15107 10195 15113
rect 10796 15116 13176 15144
rect 4430 15036 4436 15088
rect 4488 15076 4494 15088
rect 4985 15079 5043 15085
rect 4985 15076 4997 15079
rect 4488 15048 4997 15076
rect 4488 15036 4494 15048
rect 4985 15045 4997 15048
rect 5031 15045 5043 15079
rect 9766 15076 9772 15088
rect 4985 15039 5043 15045
rect 5276 15048 9772 15076
rect 4341 15011 4399 15017
rect 4341 15008 4353 15011
rect 1504 14980 2452 15008
rect 3712 14980 4353 15008
rect 1504 14949 1532 14980
rect 1489 14943 1547 14949
rect 1489 14909 1501 14943
rect 1535 14909 1547 14943
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1489 14903 1547 14909
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 2317 14943 2375 14949
rect 2317 14909 2329 14943
rect 2363 14909 2375 14943
rect 2424 14940 2452 14980
rect 4341 14977 4353 14980
rect 4387 14977 4399 15011
rect 4341 14971 4399 14977
rect 5276 14940 5304 15048
rect 9766 15036 9772 15048
rect 9824 15036 9830 15088
rect 10226 15076 10232 15088
rect 9876 15048 10232 15076
rect 5534 15008 5540 15020
rect 5495 14980 5540 15008
rect 5534 14968 5540 14980
rect 5592 15008 5598 15020
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 5592 14980 6377 15008
rect 5592 14968 5598 14980
rect 6365 14977 6377 14980
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 7374 15008 7380 15020
rect 6788 14980 7236 15008
rect 7335 14980 7380 15008
rect 6788 14968 6794 14980
rect 2424 14912 5304 14940
rect 5353 14943 5411 14949
rect 2317 14903 2375 14909
rect 5353 14909 5365 14943
rect 5399 14940 5411 14943
rect 5442 14940 5448 14952
rect 5399 14912 5448 14940
rect 5399 14909 5411 14912
rect 5353 14903 5411 14909
rect 2332 14804 2360 14903
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 6273 14943 6331 14949
rect 6273 14909 6285 14943
rect 6319 14940 6331 14943
rect 6822 14940 6828 14952
rect 6319 14912 6828 14940
rect 6319 14909 6331 14912
rect 6273 14903 6331 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 7208 14940 7236 14980
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 7834 14968 7840 15020
rect 7892 15008 7898 15020
rect 8205 15011 8263 15017
rect 8205 15008 8217 15011
rect 7892 14980 8217 15008
rect 7892 14968 7898 14980
rect 8205 14977 8217 14980
rect 8251 14977 8263 15011
rect 9030 15008 9036 15020
rect 8991 14980 9036 15008
rect 8205 14971 8263 14977
rect 9030 14968 9036 14980
rect 9088 15008 9094 15020
rect 9876 15017 9904 15048
rect 10226 15036 10232 15048
rect 10284 15036 10290 15088
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 9088 14980 9873 15008
rect 9088 14968 9094 14980
rect 9861 14977 9873 14980
rect 9907 14977 9919 15011
rect 9861 14971 9919 14977
rect 9950 14968 9956 15020
rect 10008 15008 10014 15020
rect 10689 15011 10747 15017
rect 10689 15008 10701 15011
rect 10008 14980 10701 15008
rect 10008 14968 10014 14980
rect 10689 14977 10701 14980
rect 10735 14977 10747 15011
rect 10689 14971 10747 14977
rect 8021 14943 8079 14949
rect 8021 14940 8033 14943
rect 7208 14912 8033 14940
rect 8021 14909 8033 14912
rect 8067 14909 8079 14943
rect 8021 14903 8079 14909
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14940 9827 14943
rect 10134 14940 10140 14952
rect 9815 14912 10140 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 10134 14900 10140 14912
rect 10192 14940 10198 14952
rect 10796 14940 10824 15116
rect 13170 15104 13176 15116
rect 13228 15144 13234 15156
rect 16574 15144 16580 15156
rect 13228 15116 16580 15144
rect 13228 15104 13234 15116
rect 16574 15104 16580 15116
rect 16632 15104 16638 15156
rect 10965 15079 11023 15085
rect 10965 15045 10977 15079
rect 11011 15076 11023 15079
rect 11330 15076 11336 15088
rect 11011 15048 11336 15076
rect 11011 15045 11023 15048
rect 10965 15039 11023 15045
rect 11330 15036 11336 15048
rect 11388 15036 11394 15088
rect 12894 15036 12900 15088
rect 12952 15076 12958 15088
rect 13078 15076 13084 15088
rect 12952 15048 13084 15076
rect 12952 15036 12958 15048
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 11422 15008 11428 15020
rect 11383 14980 11428 15008
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 11606 15008 11612 15020
rect 11567 14980 11612 15008
rect 11606 14968 11612 14980
rect 11664 14968 11670 15020
rect 12250 14968 12256 15020
rect 12308 15008 12314 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12308 14980 13001 15008
rect 12308 14968 12314 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 10192 14912 10824 14940
rect 10192 14900 10198 14912
rect 2584 14875 2642 14881
rect 2584 14841 2596 14875
rect 2630 14872 2642 14875
rect 3234 14872 3240 14884
rect 2630 14844 3240 14872
rect 2630 14841 2642 14844
rect 2584 14835 2642 14841
rect 3234 14832 3240 14844
rect 3292 14832 3298 14884
rect 4157 14875 4215 14881
rect 4157 14841 4169 14875
rect 4203 14872 4215 14875
rect 4430 14872 4436 14884
rect 4203 14844 4436 14872
rect 4203 14841 4215 14844
rect 4157 14835 4215 14841
rect 4430 14832 4436 14844
rect 4488 14872 4494 14884
rect 4801 14875 4859 14881
rect 4801 14872 4813 14875
rect 4488 14844 4813 14872
rect 4488 14832 4494 14844
rect 4801 14841 4813 14844
rect 4847 14841 4859 14875
rect 4801 14835 4859 14841
rect 6181 14875 6239 14881
rect 6181 14841 6193 14875
rect 6227 14872 6239 14875
rect 8941 14875 8999 14881
rect 8941 14872 8953 14875
rect 6227 14844 6868 14872
rect 6227 14841 6239 14844
rect 6181 14835 6239 14841
rect 2682 14804 2688 14816
rect 2332 14776 2688 14804
rect 2682 14764 2688 14776
rect 2740 14764 2746 14816
rect 3786 14764 3792 14816
rect 3844 14804 3850 14816
rect 4246 14804 4252 14816
rect 3844 14776 4252 14804
rect 3844 14764 3850 14776
rect 4246 14764 4252 14776
rect 4304 14804 4310 14816
rect 4617 14807 4675 14813
rect 4617 14804 4629 14807
rect 4304 14776 4629 14804
rect 4304 14764 4310 14776
rect 4617 14773 4629 14776
rect 4663 14773 4675 14807
rect 4617 14767 4675 14773
rect 5350 14764 5356 14816
rect 5408 14804 5414 14816
rect 6840 14813 6868 14844
rect 7668 14844 8953 14872
rect 5445 14807 5503 14813
rect 5445 14804 5457 14807
rect 5408 14776 5457 14804
rect 5408 14764 5414 14776
rect 5445 14773 5457 14776
rect 5491 14773 5503 14807
rect 5445 14767 5503 14773
rect 6825 14807 6883 14813
rect 6825 14773 6837 14807
rect 6871 14773 6883 14807
rect 6825 14767 6883 14773
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 7064 14776 7205 14804
rect 7064 14764 7070 14776
rect 7193 14773 7205 14776
rect 7239 14773 7251 14807
rect 7193 14767 7251 14773
rect 7285 14807 7343 14813
rect 7285 14773 7297 14807
rect 7331 14804 7343 14807
rect 7466 14804 7472 14816
rect 7331 14776 7472 14804
rect 7331 14773 7343 14776
rect 7285 14767 7343 14773
rect 7466 14764 7472 14776
rect 7524 14764 7530 14816
rect 7668 14813 7696 14844
rect 8941 14841 8953 14844
rect 8987 14841 8999 14875
rect 10505 14875 10563 14881
rect 10505 14872 10517 14875
rect 8941 14835 8999 14841
rect 9324 14844 10517 14872
rect 7653 14807 7711 14813
rect 7653 14773 7665 14807
rect 7699 14773 7711 14807
rect 7653 14767 7711 14773
rect 7926 14764 7932 14816
rect 7984 14804 7990 14816
rect 8113 14807 8171 14813
rect 8113 14804 8125 14807
rect 7984 14776 8125 14804
rect 7984 14764 7990 14776
rect 8113 14773 8125 14776
rect 8159 14773 8171 14807
rect 8113 14767 8171 14773
rect 8754 14764 8760 14816
rect 8812 14804 8818 14816
rect 9324 14813 9352 14844
rect 10505 14841 10517 14844
rect 10551 14841 10563 14875
rect 10505 14835 10563 14841
rect 10686 14832 10692 14884
rect 10744 14872 10750 14884
rect 11977 14875 12035 14881
rect 11977 14872 11989 14875
rect 10744 14844 11989 14872
rect 10744 14832 10750 14844
rect 11977 14841 11989 14844
rect 12023 14841 12035 14875
rect 11977 14835 12035 14841
rect 12342 14832 12348 14884
rect 12400 14872 12406 14884
rect 12897 14875 12955 14881
rect 12897 14872 12909 14875
rect 12400 14844 12909 14872
rect 12400 14832 12406 14844
rect 12897 14841 12909 14844
rect 12943 14841 12955 14875
rect 12897 14835 12955 14841
rect 8849 14807 8907 14813
rect 8849 14804 8861 14807
rect 8812 14776 8861 14804
rect 8812 14764 8818 14776
rect 8849 14773 8861 14776
rect 8895 14773 8907 14807
rect 8849 14767 8907 14773
rect 9309 14807 9367 14813
rect 9309 14773 9321 14807
rect 9355 14773 9367 14807
rect 9674 14804 9680 14816
rect 9635 14776 9680 14804
rect 9309 14767 9367 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 10410 14764 10416 14816
rect 10468 14804 10474 14816
rect 10597 14807 10655 14813
rect 10597 14804 10609 14807
rect 10468 14776 10609 14804
rect 10468 14764 10474 14776
rect 10597 14773 10609 14776
rect 10643 14773 10655 14807
rect 10597 14767 10655 14773
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14804 11391 14807
rect 11790 14804 11796 14816
rect 11379 14776 11796 14804
rect 11379 14773 11391 14776
rect 11333 14767 11391 14773
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 12434 14804 12440 14816
rect 12395 14776 12440 14804
rect 12434 14764 12440 14776
rect 12492 14764 12498 14816
rect 12802 14804 12808 14816
rect 12763 14776 12808 14804
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 13265 14807 13323 14813
rect 13265 14773 13277 14807
rect 13311 14804 13323 14807
rect 13538 14804 13544 14816
rect 13311 14776 13544 14804
rect 13311 14773 13323 14776
rect 13265 14767 13323 14773
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 1104 14714 16008 14736
rect 1104 14662 5979 14714
rect 6031 14662 6043 14714
rect 6095 14662 6107 14714
rect 6159 14662 6171 14714
rect 6223 14662 10976 14714
rect 11028 14662 11040 14714
rect 11092 14662 11104 14714
rect 11156 14662 11168 14714
rect 11220 14662 16008 14714
rect 1104 14640 16008 14662
rect 3145 14603 3203 14609
rect 3145 14569 3157 14603
rect 3191 14600 3203 14603
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 3191 14572 4077 14600
rect 3191 14569 3203 14572
rect 3145 14563 3203 14569
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4065 14563 4123 14569
rect 4433 14603 4491 14609
rect 4433 14569 4445 14603
rect 4479 14600 4491 14603
rect 5353 14603 5411 14609
rect 5353 14600 5365 14603
rect 4479 14572 5365 14600
rect 4479 14569 4491 14572
rect 4433 14563 4491 14569
rect 5353 14569 5365 14572
rect 5399 14569 5411 14603
rect 5353 14563 5411 14569
rect 5813 14603 5871 14609
rect 5813 14569 5825 14603
rect 5859 14600 5871 14603
rect 6181 14603 6239 14609
rect 6181 14600 6193 14603
rect 5859 14572 6193 14600
rect 5859 14569 5871 14572
rect 5813 14563 5871 14569
rect 6181 14569 6193 14572
rect 6227 14569 6239 14603
rect 6641 14603 6699 14609
rect 6641 14600 6653 14603
rect 6181 14563 6239 14569
rect 6380 14572 6653 14600
rect 1489 14467 1547 14473
rect 1489 14433 1501 14467
rect 1535 14464 1547 14467
rect 2866 14464 2872 14476
rect 1535 14436 2872 14464
rect 1535 14433 1547 14436
rect 1489 14427 1547 14433
rect 2866 14424 2872 14436
rect 2924 14424 2930 14476
rect 3050 14464 3056 14476
rect 3011 14436 3056 14464
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 5074 14464 5080 14476
rect 5035 14436 5080 14464
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5718 14464 5724 14476
rect 5679 14436 5724 14464
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 5810 14424 5816 14476
rect 5868 14464 5874 14476
rect 6380 14464 6408 14572
rect 6641 14569 6653 14572
rect 6687 14569 6699 14603
rect 7006 14600 7012 14612
rect 6967 14572 7012 14600
rect 6641 14563 6699 14569
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 8941 14603 8999 14609
rect 7156 14572 7972 14600
rect 7156 14560 7162 14572
rect 7834 14541 7840 14544
rect 6549 14535 6607 14541
rect 6549 14501 6561 14535
rect 6595 14532 6607 14535
rect 7828 14532 7840 14541
rect 6595 14504 6868 14532
rect 7795 14504 7840 14532
rect 6595 14501 6607 14504
rect 6549 14495 6607 14501
rect 5868 14436 6408 14464
rect 5868 14424 5874 14436
rect 1670 14396 1676 14408
rect 1631 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 3234 14396 3240 14408
rect 3195 14368 3240 14396
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 4522 14396 4528 14408
rect 4483 14368 4528 14396
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 4617 14399 4675 14405
rect 4617 14365 4629 14399
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 4062 14288 4068 14340
rect 4120 14328 4126 14340
rect 4632 14328 4660 14359
rect 4890 14356 4896 14408
rect 4948 14396 4954 14408
rect 5905 14399 5963 14405
rect 5905 14396 5917 14399
rect 4948 14368 5917 14396
rect 4948 14356 4954 14368
rect 5905 14365 5917 14368
rect 5951 14365 5963 14399
rect 5905 14359 5963 14365
rect 4120 14300 4660 14328
rect 6196 14328 6224 14436
rect 6638 14424 6644 14476
rect 6696 14464 6702 14476
rect 6696 14436 6776 14464
rect 6696 14424 6702 14436
rect 6748 14405 6776 14436
rect 6733 14399 6791 14405
rect 6733 14365 6745 14399
rect 6779 14365 6791 14399
rect 6840 14396 6868 14504
rect 7828 14495 7840 14504
rect 7834 14492 7840 14495
rect 7892 14492 7898 14544
rect 7944 14532 7972 14572
rect 8941 14569 8953 14603
rect 8987 14600 8999 14603
rect 9030 14600 9036 14612
rect 8987 14572 9036 14600
rect 8987 14569 8999 14572
rect 8941 14563 8999 14569
rect 9030 14560 9036 14572
rect 9088 14600 9094 14612
rect 9309 14603 9367 14609
rect 9088 14572 9260 14600
rect 9088 14560 9094 14572
rect 8754 14532 8760 14544
rect 7944 14504 8760 14532
rect 8754 14492 8760 14504
rect 8812 14532 8818 14544
rect 9125 14535 9183 14541
rect 9125 14532 9137 14535
rect 8812 14504 9137 14532
rect 8812 14492 8818 14504
rect 9125 14501 9137 14504
rect 9171 14501 9183 14535
rect 9125 14495 9183 14501
rect 6914 14424 6920 14476
rect 6972 14464 6978 14476
rect 7561 14467 7619 14473
rect 7561 14464 7573 14467
rect 6972 14436 7573 14464
rect 6972 14424 6978 14436
rect 7561 14433 7573 14436
rect 7607 14464 7619 14467
rect 7650 14464 7656 14476
rect 7607 14436 7656 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 7098 14396 7104 14408
rect 6840 14368 7104 14396
rect 6733 14359 6791 14365
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 9232 14396 9260 14572
rect 9309 14569 9321 14603
rect 9355 14600 9367 14603
rect 9674 14600 9680 14612
rect 9355 14572 9680 14600
rect 9355 14569 9367 14572
rect 9309 14563 9367 14569
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 11422 14600 11428 14612
rect 9824 14572 11428 14600
rect 9824 14560 9830 14572
rect 11422 14560 11428 14572
rect 11480 14560 11486 14612
rect 12342 14600 12348 14612
rect 12303 14572 12348 14600
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 13173 14603 13231 14609
rect 13173 14600 13185 14603
rect 12860 14572 13185 14600
rect 12860 14560 12866 14572
rect 13173 14569 13185 14572
rect 13219 14569 13231 14603
rect 13538 14600 13544 14612
rect 13499 14572 13544 14600
rect 13173 14563 13231 14569
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 10137 14535 10195 14541
rect 10137 14501 10149 14535
rect 10183 14532 10195 14535
rect 10864 14535 10922 14541
rect 10183 14504 10824 14532
rect 10183 14501 10195 14504
rect 10137 14495 10195 14501
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 10318 14464 10324 14476
rect 10091 14436 10324 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 10796 14464 10824 14504
rect 10864 14501 10876 14535
rect 10910 14532 10922 14535
rect 11606 14532 11612 14544
rect 10910 14504 11612 14532
rect 10910 14501 10922 14504
rect 10864 14495 10922 14501
rect 11606 14492 11612 14504
rect 11664 14532 11670 14544
rect 11664 14504 12848 14532
rect 11664 14492 11670 14504
rect 11146 14464 11152 14476
rect 10796 14436 11152 14464
rect 11146 14424 11152 14436
rect 11204 14464 11210 14476
rect 11882 14464 11888 14476
rect 11204 14436 11888 14464
rect 11204 14424 11210 14436
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 12710 14464 12716 14476
rect 12671 14436 12716 14464
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 12820 14464 12848 14504
rect 12894 14492 12900 14544
rect 12952 14532 12958 14544
rect 13633 14535 13691 14541
rect 13633 14532 13645 14535
rect 12952 14504 13645 14532
rect 12952 14492 12958 14504
rect 13633 14501 13645 14504
rect 13679 14532 13691 14535
rect 14369 14535 14427 14541
rect 14369 14532 14381 14535
rect 13679 14504 14381 14532
rect 13679 14501 13691 14504
rect 13633 14495 13691 14501
rect 14369 14501 14381 14504
rect 14415 14532 14427 14535
rect 16942 14532 16948 14544
rect 14415 14504 16948 14532
rect 14415 14501 14427 14504
rect 14369 14495 14427 14501
rect 16942 14492 16948 14504
rect 17000 14492 17006 14544
rect 12986 14464 12992 14476
rect 12820 14436 12992 14464
rect 12912 14405 12940 14436
rect 12986 14424 12992 14436
rect 13044 14464 13050 14476
rect 13044 14436 13768 14464
rect 13044 14424 13050 14436
rect 13740 14405 13768 14436
rect 10229 14399 10287 14405
rect 10229 14396 10241 14399
rect 9232 14368 10241 14396
rect 10229 14365 10241 14368
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14365 10655 14399
rect 10597 14359 10655 14365
rect 12805 14399 12863 14405
rect 12805 14365 12817 14399
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 12897 14399 12955 14405
rect 12897 14365 12909 14399
rect 12943 14365 12955 14399
rect 12897 14359 12955 14365
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14365 13783 14399
rect 13725 14359 13783 14365
rect 7285 14331 7343 14337
rect 7285 14328 7297 14331
rect 6196 14300 7297 14328
rect 4120 14288 4126 14300
rect 7285 14297 7297 14300
rect 7331 14297 7343 14331
rect 7285 14291 7343 14297
rect 9677 14331 9735 14337
rect 9677 14297 9689 14331
rect 9723 14328 9735 14331
rect 10410 14328 10416 14340
rect 9723 14300 10416 14328
rect 9723 14297 9735 14300
rect 9677 14291 9735 14297
rect 10410 14288 10416 14300
rect 10468 14288 10474 14340
rect 1578 14220 1584 14272
rect 1636 14260 1642 14272
rect 2685 14263 2743 14269
rect 2685 14260 2697 14263
rect 1636 14232 2697 14260
rect 1636 14220 1642 14232
rect 2685 14229 2697 14232
rect 2731 14229 2743 14263
rect 2685 14223 2743 14229
rect 4614 14220 4620 14272
rect 4672 14260 4678 14272
rect 4893 14263 4951 14269
rect 4893 14260 4905 14263
rect 4672 14232 4905 14260
rect 4672 14220 4678 14232
rect 4893 14229 4905 14232
rect 4939 14260 4951 14263
rect 4982 14260 4988 14272
rect 4939 14232 4988 14260
rect 4939 14229 4951 14232
rect 4893 14223 4951 14229
rect 4982 14220 4988 14232
rect 5040 14220 5046 14272
rect 5166 14260 5172 14272
rect 5127 14232 5172 14260
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 5258 14220 5264 14272
rect 5316 14260 5322 14272
rect 7374 14260 7380 14272
rect 5316 14232 7380 14260
rect 5316 14220 5322 14232
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 10612 14260 10640 14359
rect 12066 14328 12072 14340
rect 11532 14300 12072 14328
rect 11532 14260 11560 14300
rect 12066 14288 12072 14300
rect 12124 14288 12130 14340
rect 12710 14288 12716 14340
rect 12768 14328 12774 14340
rect 12820 14328 12848 14359
rect 14185 14331 14243 14337
rect 14185 14328 14197 14331
rect 12768 14300 14197 14328
rect 12768 14288 12774 14300
rect 14185 14297 14197 14300
rect 14231 14328 14243 14331
rect 15470 14328 15476 14340
rect 14231 14300 15476 14328
rect 14231 14297 14243 14300
rect 14185 14291 14243 14297
rect 15470 14288 15476 14300
rect 15528 14288 15534 14340
rect 10612 14232 11560 14260
rect 11977 14263 12035 14269
rect 11977 14229 11989 14263
rect 12023 14260 12035 14263
rect 12250 14260 12256 14272
rect 12023 14232 12256 14260
rect 12023 14229 12035 14232
rect 11977 14223 12035 14229
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 13262 14260 13268 14272
rect 12860 14232 13268 14260
rect 12860 14220 12866 14232
rect 13262 14220 13268 14232
rect 13320 14260 13326 14272
rect 14001 14263 14059 14269
rect 14001 14260 14013 14263
rect 13320 14232 14013 14260
rect 13320 14220 13326 14232
rect 14001 14229 14013 14232
rect 14047 14229 14059 14263
rect 14001 14223 14059 14229
rect 1104 14170 16008 14192
rect 1104 14118 3480 14170
rect 3532 14118 3544 14170
rect 3596 14118 3608 14170
rect 3660 14118 3672 14170
rect 3724 14118 8478 14170
rect 8530 14118 8542 14170
rect 8594 14118 8606 14170
rect 8658 14118 8670 14170
rect 8722 14118 13475 14170
rect 13527 14118 13539 14170
rect 13591 14118 13603 14170
rect 13655 14118 13667 14170
rect 13719 14118 16008 14170
rect 1104 14096 16008 14118
rect 2958 14016 2964 14068
rect 3016 14056 3022 14068
rect 4062 14056 4068 14068
rect 3016 14028 3924 14056
rect 4023 14028 4068 14056
rect 3016 14016 3022 14028
rect 3896 13988 3924 14028
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 4706 14016 4712 14068
rect 4764 14016 4770 14068
rect 8297 14059 8355 14065
rect 8297 14056 8309 14059
rect 6932 14028 8309 14056
rect 4724 13988 4752 14016
rect 6089 13991 6147 13997
rect 6089 13988 6101 13991
rect 3896 13960 6101 13988
rect 2682 13920 2688 13932
rect 2643 13892 2688 13920
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 4709 13923 4767 13929
rect 4709 13920 4721 13923
rect 4540 13892 4721 13920
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 1854 13852 1860 13864
rect 1815 13824 1860 13852
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 2952 13855 3010 13861
rect 2952 13821 2964 13855
rect 2998 13852 3010 13855
rect 4540 13852 4568 13892
rect 4709 13889 4721 13892
rect 4755 13920 4767 13923
rect 4890 13920 4896 13932
rect 4755 13892 4896 13920
rect 4755 13889 4767 13892
rect 4709 13883 4767 13889
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 2998 13824 4568 13852
rect 4617 13855 4675 13861
rect 2998 13821 3010 13824
rect 2952 13815 3010 13821
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 5166 13852 5172 13864
rect 4663 13824 5172 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 3970 13744 3976 13796
rect 4028 13784 4034 13796
rect 4632 13784 4660 13815
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 5258 13812 5264 13864
rect 5316 13812 5322 13864
rect 5276 13784 5304 13812
rect 4028 13756 4660 13784
rect 5000 13756 5304 13784
rect 4028 13744 4034 13756
rect 4154 13676 4160 13728
rect 4212 13716 4218 13728
rect 4525 13719 4583 13725
rect 4212 13688 4257 13716
rect 4212 13676 4218 13688
rect 4525 13685 4537 13719
rect 4571 13716 4583 13719
rect 4614 13716 4620 13728
rect 4571 13688 4620 13716
rect 4571 13685 4583 13688
rect 4525 13679 4583 13685
rect 4614 13676 4620 13688
rect 4672 13716 4678 13728
rect 5000 13725 5028 13756
rect 4985 13719 5043 13725
rect 4985 13716 4997 13719
rect 4672 13688 4997 13716
rect 4672 13676 4678 13688
rect 4985 13685 4997 13688
rect 5031 13685 5043 13719
rect 5258 13716 5264 13728
rect 5219 13688 5264 13716
rect 4985 13679 5043 13685
rect 5258 13676 5264 13688
rect 5316 13676 5322 13728
rect 5460 13716 5488 13960
rect 6089 13957 6101 13960
rect 6135 13988 6147 13991
rect 6362 13988 6368 14000
rect 6135 13960 6368 13988
rect 6135 13957 6147 13960
rect 6089 13951 6147 13957
rect 6362 13948 6368 13960
rect 6420 13948 6426 14000
rect 6638 13988 6644 14000
rect 6472 13960 6644 13988
rect 5534 13880 5540 13932
rect 5592 13920 5598 13932
rect 5905 13923 5963 13929
rect 5905 13920 5917 13923
rect 5592 13892 5917 13920
rect 5592 13880 5598 13892
rect 5905 13889 5917 13892
rect 5951 13920 5963 13923
rect 6472 13920 6500 13960
rect 6638 13948 6644 13960
rect 6696 13988 6702 14000
rect 6932 13988 6960 14028
rect 8297 14025 8309 14028
rect 8343 14025 8355 14059
rect 8297 14019 8355 14025
rect 8846 14016 8852 14068
rect 8904 14056 8910 14068
rect 9766 14056 9772 14068
rect 8904 14028 9772 14056
rect 8904 14016 8910 14028
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10134 14056 10140 14068
rect 10095 14028 10140 14056
rect 10134 14016 10140 14028
rect 10192 14016 10198 14068
rect 10781 14059 10839 14065
rect 10781 14025 10793 14059
rect 10827 14056 10839 14059
rect 11146 14056 11152 14068
rect 10827 14028 11152 14056
rect 10827 14025 10839 14028
rect 10781 14019 10839 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 12250 14056 12256 14068
rect 11808 14028 12256 14056
rect 8757 13991 8815 13997
rect 8757 13988 8769 13991
rect 6696 13960 6960 13988
rect 7944 13960 8769 13988
rect 6696 13948 6702 13960
rect 5951 13892 6500 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 6914 13880 6920 13932
rect 6972 13920 6978 13932
rect 6972 13892 7017 13920
rect 6972 13880 6978 13892
rect 5718 13812 5724 13864
rect 5776 13852 5782 13864
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 5776 13824 6377 13852
rect 5776 13812 5782 13824
rect 6365 13821 6377 13824
rect 6411 13852 6423 13855
rect 6546 13852 6552 13864
rect 6411 13824 6552 13852
rect 6411 13821 6423 13824
rect 6365 13815 6423 13821
rect 6546 13812 6552 13824
rect 6604 13812 6610 13864
rect 7466 13812 7472 13864
rect 7524 13852 7530 13864
rect 7944 13852 7972 13960
rect 8757 13957 8769 13960
rect 8803 13988 8815 13991
rect 8803 13960 11008 13988
rect 8803 13957 8815 13960
rect 8757 13951 8815 13957
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 10778 13920 10784 13932
rect 8996 13892 10784 13920
rect 8996 13880 9002 13892
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 10980 13920 11008 13960
rect 11054 13948 11060 14000
rect 11112 13988 11118 14000
rect 11606 13988 11612 14000
rect 11112 13960 11612 13988
rect 11112 13948 11118 13960
rect 11606 13948 11612 13960
rect 11664 13948 11670 14000
rect 11517 13923 11575 13929
rect 10980 13892 11468 13920
rect 8018 13852 8024 13864
rect 7524 13824 8024 13852
rect 7524 13812 7530 13824
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13852 8631 13855
rect 9858 13852 9864 13864
rect 8619 13824 9864 13852
rect 8619 13821 8631 13824
rect 8573 13815 8631 13821
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 10410 13812 10416 13864
rect 10468 13852 10474 13864
rect 10505 13855 10563 13861
rect 10505 13852 10517 13855
rect 10468 13824 10517 13852
rect 10468 13812 10474 13824
rect 10505 13821 10517 13824
rect 10551 13821 10563 13855
rect 11330 13852 11336 13864
rect 10505 13815 10563 13821
rect 11256 13824 11336 13852
rect 5629 13787 5687 13793
rect 5629 13753 5641 13787
rect 5675 13784 5687 13787
rect 7184 13787 7242 13793
rect 5675 13756 6592 13784
rect 5675 13753 5687 13756
rect 5629 13747 5687 13753
rect 6564 13725 6592 13756
rect 7184 13753 7196 13787
rect 7230 13784 7242 13787
rect 7374 13784 7380 13796
rect 7230 13756 7380 13784
rect 7230 13753 7242 13756
rect 7184 13747 7242 13753
rect 7374 13744 7380 13756
rect 7432 13744 7438 13796
rect 8846 13784 8852 13796
rect 7484 13756 8852 13784
rect 5721 13719 5779 13725
rect 5721 13716 5733 13719
rect 5460 13688 5733 13716
rect 5721 13685 5733 13688
rect 5767 13685 5779 13719
rect 5721 13679 5779 13685
rect 6549 13719 6607 13725
rect 6549 13685 6561 13719
rect 6595 13716 6607 13719
rect 6730 13716 6736 13728
rect 6595 13688 6736 13716
rect 6595 13685 6607 13688
rect 6549 13679 6607 13685
rect 6730 13676 6736 13688
rect 6788 13676 6794 13728
rect 7098 13676 7104 13728
rect 7156 13716 7162 13728
rect 7484 13716 7512 13756
rect 8846 13744 8852 13756
rect 8904 13744 8910 13796
rect 11054 13744 11060 13796
rect 11112 13744 11118 13796
rect 11256 13793 11284 13824
rect 11330 13812 11336 13824
rect 11388 13812 11394 13864
rect 11241 13787 11299 13793
rect 11241 13753 11253 13787
rect 11287 13753 11299 13787
rect 11440 13784 11468 13892
rect 11517 13889 11529 13923
rect 11563 13920 11575 13923
rect 11808 13920 11836 14028
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 11563 13892 11836 13920
rect 11563 13889 11575 13892
rect 11517 13883 11575 13889
rect 12250 13880 12256 13932
rect 12308 13920 12314 13932
rect 12308 13892 12572 13920
rect 12308 13880 12314 13892
rect 12066 13812 12072 13864
rect 12124 13852 12130 13864
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12124 13824 12449 13852
rect 12124 13812 12130 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12544 13852 12572 13892
rect 12693 13855 12751 13861
rect 12693 13852 12705 13855
rect 12544 13824 12705 13852
rect 12437 13815 12495 13821
rect 12693 13821 12705 13824
rect 12739 13821 12751 13855
rect 12693 13815 12751 13821
rect 16206 13784 16212 13796
rect 11440 13756 16212 13784
rect 11241 13747 11299 13753
rect 16206 13744 16212 13756
rect 16264 13744 16270 13796
rect 7156 13688 7512 13716
rect 10873 13719 10931 13725
rect 7156 13676 7162 13688
rect 10873 13685 10885 13719
rect 10919 13716 10931 13719
rect 11072 13716 11100 13744
rect 10919 13688 11100 13716
rect 11333 13719 11391 13725
rect 10919 13685 10931 13688
rect 10873 13679 10931 13685
rect 11333 13685 11345 13719
rect 11379 13716 11391 13719
rect 12618 13716 12624 13728
rect 11379 13688 12624 13716
rect 11379 13685 11391 13688
rect 11333 13679 11391 13685
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 13262 13676 13268 13728
rect 13320 13716 13326 13728
rect 13817 13719 13875 13725
rect 13817 13716 13829 13719
rect 13320 13688 13829 13716
rect 13320 13676 13326 13688
rect 13817 13685 13829 13688
rect 13863 13685 13875 13719
rect 13817 13679 13875 13685
rect 1104 13626 16008 13648
rect 1104 13574 5979 13626
rect 6031 13574 6043 13626
rect 6095 13574 6107 13626
rect 6159 13574 6171 13626
rect 6223 13574 10976 13626
rect 11028 13574 11040 13626
rect 11092 13574 11104 13626
rect 11156 13574 11168 13626
rect 11220 13574 16008 13626
rect 1104 13552 16008 13574
rect 3145 13515 3203 13521
rect 3145 13481 3157 13515
rect 3191 13512 3203 13515
rect 3234 13512 3240 13524
rect 3191 13484 3240 13512
rect 3191 13481 3203 13484
rect 3145 13475 3203 13481
rect 3234 13472 3240 13484
rect 3292 13472 3298 13524
rect 4341 13515 4399 13521
rect 4341 13481 4353 13515
rect 4387 13512 4399 13515
rect 4522 13512 4528 13524
rect 4387 13484 4528 13512
rect 4387 13481 4399 13484
rect 4341 13475 4399 13481
rect 4522 13472 4528 13484
rect 4580 13472 4586 13524
rect 4801 13515 4859 13521
rect 4801 13481 4813 13515
rect 4847 13512 4859 13515
rect 5258 13512 5264 13524
rect 4847 13484 5264 13512
rect 4847 13481 4859 13484
rect 4801 13475 4859 13481
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 6638 13472 6644 13524
rect 6696 13512 6702 13524
rect 6696 13484 7052 13512
rect 6696 13472 6702 13484
rect 2032 13447 2090 13453
rect 2032 13413 2044 13447
rect 2078 13444 2090 13447
rect 4062 13444 4068 13456
rect 2078 13416 4068 13444
rect 2078 13413 2090 13416
rect 2032 13407 2090 13413
rect 4062 13404 4068 13416
rect 4120 13404 4126 13456
rect 5436 13447 5494 13453
rect 5436 13413 5448 13447
rect 5482 13444 5494 13447
rect 5534 13444 5540 13456
rect 5482 13416 5540 13444
rect 5482 13413 5494 13416
rect 5436 13407 5494 13413
rect 5534 13404 5540 13416
rect 5592 13404 5598 13456
rect 6914 13444 6920 13456
rect 6748 13416 6920 13444
rect 1765 13379 1823 13385
rect 1765 13345 1777 13379
rect 1811 13376 1823 13379
rect 2590 13376 2596 13388
rect 1811 13348 2596 13376
rect 1811 13345 1823 13348
rect 1765 13339 1823 13345
rect 2590 13336 2596 13348
rect 2648 13336 2654 13388
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 5258 13376 5264 13388
rect 4755 13348 5264 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 6748 13385 6776 13416
rect 6914 13404 6920 13416
rect 6972 13404 6978 13456
rect 7024 13444 7052 13484
rect 9214 13472 9220 13524
rect 9272 13512 9278 13524
rect 9309 13515 9367 13521
rect 9309 13512 9321 13515
rect 9272 13484 9321 13512
rect 9272 13472 9278 13484
rect 9309 13481 9321 13484
rect 9355 13481 9367 13515
rect 9309 13475 9367 13481
rect 11149 13515 11207 13521
rect 11149 13481 11161 13515
rect 11195 13512 11207 13515
rect 11422 13512 11428 13524
rect 11195 13484 11428 13512
rect 11195 13481 11207 13484
rect 11149 13475 11207 13481
rect 11422 13472 11428 13484
rect 11480 13472 11486 13524
rect 11606 13512 11612 13524
rect 11567 13484 11612 13512
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 11517 13447 11575 13453
rect 7024 13416 11468 13444
rect 6733 13379 6791 13385
rect 6733 13345 6745 13379
rect 6779 13345 6791 13379
rect 6733 13339 6791 13345
rect 7000 13379 7058 13385
rect 7000 13345 7012 13379
rect 7046 13376 7058 13379
rect 8202 13376 8208 13388
rect 7046 13348 8208 13376
rect 7046 13345 7058 13348
rect 7000 13339 7058 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 8849 13379 8907 13385
rect 8849 13376 8861 13379
rect 8772 13348 8861 13376
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13308 4123 13311
rect 4338 13308 4344 13320
rect 4111 13280 4344 13308
rect 4111 13277 4123 13280
rect 4065 13271 4123 13277
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 4890 13308 4896 13320
rect 4851 13280 4896 13308
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 4982 13268 4988 13320
rect 5040 13308 5046 13320
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 5040 13280 5181 13308
rect 5040 13268 5046 13280
rect 5169 13277 5181 13280
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 4890 13132 4896 13184
rect 4948 13172 4954 13184
rect 6549 13175 6607 13181
rect 6549 13172 6561 13175
rect 4948 13144 6561 13172
rect 4948 13132 4954 13144
rect 6549 13141 6561 13144
rect 6595 13141 6607 13175
rect 6549 13135 6607 13141
rect 7374 13132 7380 13184
rect 7432 13172 7438 13184
rect 8113 13175 8171 13181
rect 8113 13172 8125 13175
rect 7432 13144 8125 13172
rect 7432 13132 7438 13144
rect 8113 13141 8125 13144
rect 8159 13141 8171 13175
rect 8113 13135 8171 13141
rect 8294 13132 8300 13184
rect 8352 13172 8358 13184
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 8352 13144 8493 13172
rect 8352 13132 8358 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 8772 13172 8800 13348
rect 8849 13345 8861 13348
rect 8895 13345 8907 13379
rect 9490 13376 9496 13388
rect 9451 13348 9496 13376
rect 8849 13339 8907 13345
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 10689 13379 10747 13385
rect 10689 13345 10701 13379
rect 10735 13376 10747 13379
rect 11330 13376 11336 13388
rect 10735 13348 11336 13376
rect 10735 13345 10747 13348
rect 10689 13339 10747 13345
rect 11330 13336 11336 13348
rect 11388 13336 11394 13388
rect 11440 13376 11468 13416
rect 11517 13413 11529 13447
rect 11563 13444 11575 13447
rect 12434 13444 12440 13456
rect 11563 13416 12440 13444
rect 11563 13413 11575 13416
rect 11517 13407 11575 13413
rect 12434 13404 12440 13416
rect 12492 13404 12498 13456
rect 15838 13376 15844 13388
rect 11440 13348 15844 13376
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13308 9183 13311
rect 9306 13308 9312 13320
rect 9171 13280 9312 13308
rect 9171 13277 9183 13280
rect 9125 13271 9183 13277
rect 8846 13200 8852 13252
rect 8904 13240 8910 13252
rect 8956 13240 8984 13271
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 9398 13268 9404 13320
rect 9456 13308 9462 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 9456 13280 9781 13308
rect 9456 13268 9462 13280
rect 9769 13277 9781 13280
rect 9815 13308 9827 13311
rect 10226 13308 10232 13320
rect 9815 13280 10232 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 10778 13308 10784 13320
rect 10739 13280 10784 13308
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 10870 13268 10876 13320
rect 10928 13308 10934 13320
rect 11793 13311 11851 13317
rect 10928 13280 10973 13308
rect 10928 13268 10934 13280
rect 11793 13277 11805 13311
rect 11839 13308 11851 13311
rect 13262 13308 13268 13320
rect 11839 13280 13268 13308
rect 11839 13277 11851 13280
rect 11793 13271 11851 13277
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 8904 13212 8984 13240
rect 8904 13200 8910 13212
rect 9398 13172 9404 13184
rect 8772 13144 9404 13172
rect 8481 13135 8539 13141
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 10318 13172 10324 13184
rect 10279 13144 10324 13172
rect 10318 13132 10324 13144
rect 10376 13132 10382 13184
rect 1104 13082 16008 13104
rect 1104 13030 3480 13082
rect 3532 13030 3544 13082
rect 3596 13030 3608 13082
rect 3660 13030 3672 13082
rect 3724 13030 8478 13082
rect 8530 13030 8542 13082
rect 8594 13030 8606 13082
rect 8658 13030 8670 13082
rect 8722 13030 13475 13082
rect 13527 13030 13539 13082
rect 13591 13030 13603 13082
rect 13655 13030 13667 13082
rect 13719 13030 16008 13082
rect 1104 13008 16008 13030
rect 3050 12928 3056 12980
rect 3108 12968 3114 12980
rect 3145 12971 3203 12977
rect 3145 12968 3157 12971
rect 3108 12940 3157 12968
rect 3108 12928 3114 12940
rect 3145 12937 3157 12940
rect 3191 12937 3203 12971
rect 3145 12931 3203 12937
rect 4985 12971 5043 12977
rect 4985 12937 4997 12971
rect 5031 12968 5043 12971
rect 5074 12968 5080 12980
rect 5031 12940 5080 12968
rect 5031 12937 5043 12940
rect 4985 12931 5043 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5258 12968 5264 12980
rect 5219 12940 5264 12968
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 10318 12968 10324 12980
rect 7208 12940 10324 12968
rect 4801 12903 4859 12909
rect 4801 12900 4813 12903
rect 4448 12872 4813 12900
rect 3789 12835 3847 12841
rect 3789 12801 3801 12835
rect 3835 12832 3847 12835
rect 4062 12832 4068 12844
rect 3835 12804 4068 12832
rect 3835 12801 3847 12804
rect 3789 12795 3847 12801
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4448 12841 4476 12872
rect 4801 12869 4813 12872
rect 4847 12900 4859 12903
rect 6638 12900 6644 12912
rect 4847 12872 6644 12900
rect 4847 12869 4859 12872
rect 4801 12863 4859 12869
rect 6638 12860 6644 12872
rect 6696 12860 6702 12912
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12801 4491 12835
rect 4433 12795 4491 12801
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4890 12832 4896 12844
rect 4663 12804 4896 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5592 12804 5825 12832
rect 5592 12792 5598 12804
rect 5813 12801 5825 12804
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 6089 12835 6147 12841
rect 6089 12801 6101 12835
rect 6135 12832 6147 12835
rect 6454 12832 6460 12844
rect 6135 12804 6460 12832
rect 6135 12801 6147 12804
rect 6089 12795 6147 12801
rect 6454 12792 6460 12804
rect 6512 12832 6518 12844
rect 6914 12832 6920 12844
rect 6512 12804 6920 12832
rect 6512 12792 6518 12804
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12764 3663 12767
rect 4154 12764 4160 12776
rect 3651 12736 4160 12764
rect 3651 12733 3663 12736
rect 3605 12727 3663 12733
rect 4154 12724 4160 12736
rect 4212 12724 4218 12776
rect 4338 12764 4344 12776
rect 4299 12736 4344 12764
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 7208 12773 7236 12940
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 10778 12928 10784 12980
rect 10836 12968 10842 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 10836 12940 10885 12968
rect 10836 12928 10842 12940
rect 10873 12937 10885 12940
rect 10919 12937 10931 12971
rect 10873 12931 10931 12937
rect 11977 12971 12035 12977
rect 11977 12937 11989 12971
rect 12023 12968 12035 12971
rect 12434 12968 12440 12980
rect 12023 12940 12440 12968
rect 12023 12937 12035 12940
rect 11977 12931 12035 12937
rect 9030 12860 9036 12912
rect 9088 12900 9094 12912
rect 9306 12900 9312 12912
rect 9088 12872 9312 12900
rect 9088 12860 9094 12872
rect 9306 12860 9312 12872
rect 9364 12860 9370 12912
rect 7374 12832 7380 12844
rect 7335 12804 7380 12832
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 8202 12832 8208 12844
rect 8163 12804 8208 12832
rect 8202 12792 8208 12804
rect 8260 12832 8266 12844
rect 9125 12835 9183 12841
rect 8260 12804 9076 12832
rect 8260 12792 8266 12804
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12764 5227 12767
rect 7193 12767 7251 12773
rect 5215 12736 6776 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 3513 12699 3571 12705
rect 3513 12665 3525 12699
rect 3559 12696 3571 12699
rect 3559 12668 4016 12696
rect 3559 12665 3571 12668
rect 3513 12659 3571 12665
rect 3988 12637 4016 12668
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 4614 12696 4620 12708
rect 4120 12668 4620 12696
rect 4120 12656 4126 12668
rect 4614 12656 4620 12668
rect 4672 12656 4678 12708
rect 6273 12699 6331 12705
rect 6273 12696 6285 12699
rect 5644 12668 6285 12696
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12597 4031 12631
rect 3973 12591 4031 12597
rect 5534 12588 5540 12640
rect 5592 12628 5598 12640
rect 5644 12637 5672 12668
rect 6273 12665 6285 12668
rect 6319 12665 6331 12699
rect 6748 12696 6776 12736
rect 7193 12733 7205 12767
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 8294 12764 8300 12776
rect 8067 12736 8300 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 7374 12696 7380 12708
rect 6748 12668 7380 12696
rect 6273 12659 6331 12665
rect 7374 12656 7380 12668
rect 7432 12656 7438 12708
rect 8754 12656 8760 12708
rect 8812 12696 8818 12708
rect 8941 12699 8999 12705
rect 8941 12696 8953 12699
rect 8812 12668 8953 12696
rect 8812 12656 8818 12668
rect 8941 12665 8953 12668
rect 8987 12665 8999 12699
rect 8941 12659 8999 12665
rect 5629 12631 5687 12637
rect 5629 12628 5641 12631
rect 5592 12600 5641 12628
rect 5592 12588 5598 12600
rect 5629 12597 5641 12600
rect 5675 12597 5687 12631
rect 5629 12591 5687 12597
rect 5721 12631 5779 12637
rect 5721 12597 5733 12631
rect 5767 12628 5779 12631
rect 6454 12628 6460 12640
rect 5767 12600 6460 12628
rect 5767 12597 5779 12600
rect 5721 12591 5779 12597
rect 6454 12588 6460 12600
rect 6512 12588 6518 12640
rect 6822 12628 6828 12640
rect 6783 12600 6828 12628
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7285 12631 7343 12637
rect 7285 12597 7297 12631
rect 7331 12628 7343 12631
rect 7653 12631 7711 12637
rect 7653 12628 7665 12631
rect 7331 12600 7665 12628
rect 7331 12597 7343 12600
rect 7285 12591 7343 12597
rect 7653 12597 7665 12600
rect 7699 12597 7711 12631
rect 7653 12591 7711 12597
rect 8113 12631 8171 12637
rect 8113 12597 8125 12631
rect 8159 12628 8171 12631
rect 8481 12631 8539 12637
rect 8481 12628 8493 12631
rect 8159 12600 8493 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8481 12597 8493 12600
rect 8527 12597 8539 12631
rect 8846 12628 8852 12640
rect 8807 12600 8852 12628
rect 8481 12591 8539 12597
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9048 12628 9076 12804
rect 9125 12801 9137 12835
rect 9171 12832 9183 12835
rect 11422 12832 11428 12844
rect 9171 12804 9444 12832
rect 11383 12804 11428 12832
rect 9171 12801 9183 12804
rect 9125 12795 9183 12801
rect 9416 12776 9444 12804
rect 11422 12792 11428 12804
rect 11480 12792 11486 12844
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 9122 12656 9128 12708
rect 9180 12696 9186 12708
rect 9324 12696 9352 12727
rect 9398 12724 9404 12776
rect 9456 12764 9462 12776
rect 9565 12767 9623 12773
rect 9565 12764 9577 12767
rect 9456 12736 9577 12764
rect 9456 12724 9462 12736
rect 9565 12733 9577 12736
rect 9611 12764 9623 12767
rect 11440 12764 11468 12792
rect 9611 12736 11468 12764
rect 9611 12733 9623 12736
rect 9565 12727 9623 12733
rect 9180 12668 9352 12696
rect 9180 12656 9186 12668
rect 9674 12656 9680 12708
rect 9732 12696 9738 12708
rect 9858 12696 9864 12708
rect 9732 12668 9864 12696
rect 9732 12656 9738 12668
rect 9858 12656 9864 12668
rect 9916 12656 9922 12708
rect 11333 12699 11391 12705
rect 11333 12665 11345 12699
rect 11379 12696 11391 12699
rect 11992 12696 12020 12931
rect 12434 12928 12440 12940
rect 12492 12968 12498 12980
rect 13814 12968 13820 12980
rect 12492 12940 13820 12968
rect 12492 12928 12498 12940
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 11379 12668 12020 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 10689 12631 10747 12637
rect 10689 12628 10701 12631
rect 9048 12600 10701 12628
rect 10689 12597 10701 12600
rect 10735 12628 10747 12631
rect 10870 12628 10876 12640
rect 10735 12600 10876 12628
rect 10735 12597 10747 12600
rect 10689 12591 10747 12597
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 11241 12631 11299 12637
rect 11241 12597 11253 12631
rect 11287 12628 11299 12631
rect 11790 12628 11796 12640
rect 11287 12600 11796 12628
rect 11287 12597 11299 12600
rect 11241 12591 11299 12597
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 1104 12538 16008 12560
rect 1104 12486 5979 12538
rect 6031 12486 6043 12538
rect 6095 12486 6107 12538
rect 6159 12486 6171 12538
rect 6223 12486 10976 12538
rect 11028 12486 11040 12538
rect 11092 12486 11104 12538
rect 11156 12486 11168 12538
rect 11220 12486 16008 12538
rect 1104 12464 16008 12486
rect 1504 12396 2176 12424
rect 1504 12297 1532 12396
rect 1762 12356 1768 12368
rect 1723 12328 1768 12356
rect 1762 12316 1768 12328
rect 1820 12316 1826 12368
rect 2148 12356 2176 12396
rect 5350 12384 5356 12436
rect 5408 12424 5414 12436
rect 7374 12424 7380 12436
rect 5408 12396 6960 12424
rect 7335 12396 7380 12424
rect 5408 12384 5414 12396
rect 6822 12356 6828 12368
rect 2148 12328 6828 12356
rect 6822 12316 6828 12328
rect 6880 12316 6886 12368
rect 6932 12356 6960 12396
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 7929 12427 7987 12433
rect 7929 12393 7941 12427
rect 7975 12424 7987 12427
rect 8662 12424 8668 12436
rect 7975 12396 8668 12424
rect 7975 12393 7987 12396
rect 7929 12387 7987 12393
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 8812 12396 8857 12424
rect 8812 12384 8818 12396
rect 9030 12384 9036 12436
rect 9088 12424 9094 12436
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 9088 12396 9137 12424
rect 9088 12384 9094 12396
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 9125 12387 9183 12393
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 9677 12427 9735 12433
rect 9677 12424 9689 12427
rect 9456 12396 9689 12424
rect 9456 12384 9462 12396
rect 9677 12393 9689 12396
rect 9723 12393 9735 12427
rect 11330 12424 11336 12436
rect 11291 12396 11336 12424
rect 9677 12387 9735 12393
rect 11330 12384 11336 12396
rect 11388 12384 11394 12436
rect 12529 12427 12587 12433
rect 12529 12393 12541 12427
rect 12575 12424 12587 12427
rect 12710 12424 12716 12436
rect 12575 12396 12716 12424
rect 12575 12393 12587 12396
rect 12529 12387 12587 12393
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 8386 12356 8392 12368
rect 6932 12328 8392 12356
rect 8386 12316 8392 12328
rect 8444 12316 8450 12368
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 9217 12359 9275 12365
rect 9217 12356 9229 12359
rect 8996 12328 9229 12356
rect 8996 12316 9002 12328
rect 9217 12325 9229 12328
rect 9263 12325 9275 12359
rect 9217 12319 9275 12325
rect 9582 12316 9588 12368
rect 9640 12356 9646 12368
rect 9858 12356 9864 12368
rect 9640 12328 9864 12356
rect 9640 12316 9646 12328
rect 9858 12316 9864 12328
rect 9916 12316 9922 12368
rect 6178 12297 6184 12300
rect 1499 12291 1557 12297
rect 1499 12257 1511 12291
rect 1545 12257 1557 12291
rect 1499 12251 1557 12257
rect 5445 12291 5503 12297
rect 5445 12257 5457 12291
rect 5491 12288 5503 12291
rect 6172 12288 6184 12297
rect 5491 12260 5856 12288
rect 6139 12260 6184 12288
rect 5491 12257 5503 12260
rect 5445 12251 5503 12257
rect 5166 12180 5172 12232
rect 5224 12220 5230 12232
rect 5537 12223 5595 12229
rect 5537 12220 5549 12223
rect 5224 12192 5549 12220
rect 5224 12180 5230 12192
rect 5537 12189 5549 12192
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12189 5779 12223
rect 5721 12183 5779 12189
rect 1486 12044 1492 12096
rect 1544 12084 1550 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 1544 12056 5089 12084
rect 1544 12044 1550 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5736 12084 5764 12183
rect 5828 12164 5856 12260
rect 6172 12251 6184 12260
rect 6178 12248 6184 12251
rect 6236 12248 6242 12300
rect 6454 12248 6460 12300
rect 6512 12288 6518 12300
rect 6730 12288 6736 12300
rect 6512 12260 6736 12288
rect 6512 12248 6518 12260
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 7558 12288 7564 12300
rect 7519 12260 7564 12288
rect 7558 12248 7564 12260
rect 7616 12248 7622 12300
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12288 7895 12291
rect 8202 12288 8208 12300
rect 7883 12260 8208 12288
rect 7883 12257 7895 12260
rect 7837 12251 7895 12257
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 5960 12192 6005 12220
rect 5960 12180 5966 12192
rect 7006 12180 7012 12232
rect 7064 12220 7070 12232
rect 7852 12220 7880 12251
rect 8202 12248 8208 12260
rect 8260 12288 8266 12300
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 8260 12260 8309 12288
rect 8260 12248 8266 12260
rect 8297 12257 8309 12260
rect 8343 12257 8355 12291
rect 9950 12288 9956 12300
rect 8297 12251 8355 12257
rect 9876 12260 9956 12288
rect 9876 12229 9904 12260
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 10134 12297 10140 12300
rect 10128 12251 10140 12297
rect 10192 12288 10198 12300
rect 11701 12291 11759 12297
rect 10192 12260 10228 12288
rect 10134 12248 10140 12251
rect 10192 12248 10198 12260
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 11747 12260 12173 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 12161 12251 12219 12257
rect 7064 12192 7880 12220
rect 8573 12223 8631 12229
rect 7064 12180 7070 12192
rect 8573 12189 8585 12223
rect 8619 12189 8631 12223
rect 8573 12183 8631 12189
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 5810 12112 5816 12164
rect 5868 12112 5874 12164
rect 8588 12152 8616 12183
rect 9324 12152 9352 12183
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 11793 12223 11851 12229
rect 11793 12220 11805 12223
rect 11664 12192 11805 12220
rect 11664 12180 11670 12192
rect 11793 12189 11805 12192
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 11885 12223 11943 12229
rect 11885 12189 11897 12223
rect 11931 12189 11943 12223
rect 11885 12183 11943 12189
rect 11241 12155 11299 12161
rect 8588 12124 9904 12152
rect 7282 12084 7288 12096
rect 5736 12056 7288 12084
rect 5077 12047 5135 12053
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 9030 12044 9036 12096
rect 9088 12084 9094 12096
rect 9766 12084 9772 12096
rect 9088 12056 9772 12084
rect 9088 12044 9094 12056
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 9876 12084 9904 12124
rect 11241 12121 11253 12155
rect 11287 12152 11299 12155
rect 11422 12152 11428 12164
rect 11287 12124 11428 12152
rect 11287 12121 11299 12124
rect 11241 12115 11299 12121
rect 11422 12112 11428 12124
rect 11480 12152 11486 12164
rect 11900 12152 11928 12183
rect 11480 12124 11928 12152
rect 11480 12112 11486 12124
rect 10134 12084 10140 12096
rect 9876 12056 10140 12084
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 11698 12044 11704 12096
rect 11756 12084 11762 12096
rect 12710 12084 12716 12096
rect 11756 12056 12716 12084
rect 11756 12044 11762 12056
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 1104 11994 16008 12016
rect 1104 11942 3480 11994
rect 3532 11942 3544 11994
rect 3596 11942 3608 11994
rect 3660 11942 3672 11994
rect 3724 11942 8478 11994
rect 8530 11942 8542 11994
rect 8594 11942 8606 11994
rect 8658 11942 8670 11994
rect 8722 11942 13475 11994
rect 13527 11942 13539 11994
rect 13591 11942 13603 11994
rect 13655 11942 13667 11994
rect 13719 11942 16008 11994
rect 1104 11920 16008 11942
rect 6730 11840 6736 11892
rect 6788 11880 6794 11892
rect 7098 11880 7104 11892
rect 6788 11852 7104 11880
rect 6788 11840 6794 11852
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 8404 11852 8708 11880
rect 8202 11772 8208 11824
rect 8260 11812 8266 11824
rect 8404 11812 8432 11852
rect 8260 11784 8432 11812
rect 8573 11815 8631 11821
rect 8260 11772 8266 11784
rect 8573 11781 8585 11815
rect 8619 11781 8631 11815
rect 8680 11812 8708 11852
rect 8846 11840 8852 11892
rect 8904 11880 8910 11892
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 8904 11852 9137 11880
rect 8904 11840 8910 11852
rect 9125 11849 9137 11852
rect 9171 11849 9183 11883
rect 9125 11843 9183 11849
rect 9766 11840 9772 11892
rect 9824 11880 9830 11892
rect 10502 11880 10508 11892
rect 9824 11852 10508 11880
rect 9824 11840 9830 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 10594 11812 10600 11824
rect 8680 11784 10600 11812
rect 8573 11775 8631 11781
rect 8588 11744 8616 11775
rect 10594 11772 10600 11784
rect 10652 11772 10658 11824
rect 9769 11747 9827 11753
rect 9769 11744 9781 11747
rect 8588 11716 9781 11744
rect 9769 11713 9781 11716
rect 9815 11744 9827 11747
rect 10134 11744 10140 11756
rect 9815 11716 10140 11744
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11744 10287 11747
rect 10318 11744 10324 11756
rect 10275 11716 10324 11744
rect 10275 11713 10287 11716
rect 10229 11707 10287 11713
rect 1486 11676 1492 11688
rect 1447 11648 1492 11676
rect 1486 11636 1492 11648
rect 1544 11636 1550 11688
rect 2038 11676 2044 11688
rect 1999 11648 2044 11676
rect 2038 11636 2044 11648
rect 2096 11636 2102 11688
rect 2406 11636 2412 11688
rect 2464 11676 2470 11688
rect 3237 11679 3295 11685
rect 3237 11676 3249 11679
rect 2464 11648 3249 11676
rect 2464 11636 2470 11648
rect 3237 11645 3249 11648
rect 3283 11676 3295 11679
rect 4709 11679 4767 11685
rect 4709 11676 4721 11679
rect 3283 11648 4721 11676
rect 3283 11645 3295 11648
rect 3237 11639 3295 11645
rect 4709 11645 4721 11648
rect 4755 11676 4767 11679
rect 4798 11676 4804 11688
rect 4755 11648 4804 11676
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 4798 11636 4804 11648
rect 4856 11676 4862 11688
rect 5902 11676 5908 11688
rect 4856 11648 5908 11676
rect 4856 11636 4862 11648
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 7156 11648 7205 11676
rect 7156 11636 7162 11648
rect 7193 11645 7205 11648
rect 7239 11645 7251 11679
rect 7193 11639 7251 11645
rect 7282 11636 7288 11688
rect 7340 11676 7346 11688
rect 7449 11679 7507 11685
rect 7449 11676 7461 11679
rect 7340 11648 7461 11676
rect 7340 11636 7346 11648
rect 7449 11645 7461 11648
rect 7495 11645 7507 11679
rect 7449 11639 7507 11645
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 8938 11676 8944 11688
rect 8803 11648 8944 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 8938 11636 8944 11648
rect 8996 11636 9002 11688
rect 9033 11679 9091 11685
rect 9033 11645 9045 11679
rect 9079 11676 9091 11679
rect 9490 11676 9496 11688
rect 9079 11648 9496 11676
rect 9079 11645 9091 11648
rect 9033 11639 9091 11645
rect 9490 11636 9496 11648
rect 9548 11676 9554 11688
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 9548 11648 9597 11676
rect 9548 11636 9554 11648
rect 9585 11645 9597 11648
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 1762 11608 1768 11620
rect 1723 11580 1768 11608
rect 1762 11568 1768 11580
rect 1820 11568 1826 11620
rect 2317 11611 2375 11617
rect 2317 11577 2329 11611
rect 2363 11608 2375 11611
rect 2774 11608 2780 11620
rect 2363 11580 2780 11608
rect 2363 11577 2375 11580
rect 2317 11571 2375 11577
rect 2774 11568 2780 11580
rect 2832 11568 2838 11620
rect 3504 11611 3562 11617
rect 3504 11577 3516 11611
rect 3550 11608 3562 11611
rect 3786 11608 3792 11620
rect 3550 11580 3792 11608
rect 3550 11577 3562 11580
rect 3504 11571 3562 11577
rect 3786 11568 3792 11580
rect 3844 11568 3850 11620
rect 4982 11617 4988 11620
rect 4976 11608 4988 11617
rect 4632 11580 4988 11608
rect 3142 11540 3148 11552
rect 3103 11512 3148 11540
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 4632 11549 4660 11580
rect 4976 11571 4988 11580
rect 4982 11568 4988 11571
rect 5040 11568 5046 11620
rect 7006 11608 7012 11620
rect 5092 11580 7012 11608
rect 4617 11543 4675 11549
rect 4617 11509 4629 11543
rect 4663 11509 4675 11543
rect 4617 11503 4675 11509
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 5092 11540 5120 11580
rect 7006 11568 7012 11580
rect 7064 11568 7070 11620
rect 8294 11568 8300 11620
rect 8352 11608 8358 11620
rect 8352 11580 9076 11608
rect 8352 11568 8358 11580
rect 4948 11512 5120 11540
rect 6089 11543 6147 11549
rect 4948 11500 4954 11512
rect 6089 11509 6101 11543
rect 6135 11540 6147 11543
rect 6270 11540 6276 11552
rect 6135 11512 6276 11540
rect 6135 11509 6147 11512
rect 6089 11503 6147 11509
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 6641 11543 6699 11549
rect 6641 11509 6653 11543
rect 6687 11540 6699 11543
rect 6730 11540 6736 11552
rect 6687 11512 6736 11540
rect 6687 11509 6699 11512
rect 6641 11503 6699 11509
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 6825 11543 6883 11549
rect 6825 11509 6837 11543
rect 6871 11540 6883 11543
rect 7650 11540 7656 11552
rect 6871 11512 7656 11540
rect 6871 11509 6883 11512
rect 6825 11503 6883 11509
rect 7650 11500 7656 11512
rect 7708 11500 7714 11552
rect 9048 11540 9076 11580
rect 9122 11568 9128 11620
rect 9180 11608 9186 11620
rect 9766 11608 9772 11620
rect 9180 11580 9772 11608
rect 9180 11568 9186 11580
rect 9766 11568 9772 11580
rect 9824 11608 9830 11620
rect 9953 11611 10011 11617
rect 9953 11608 9965 11611
rect 9824 11580 9965 11608
rect 9824 11568 9830 11580
rect 9953 11577 9965 11580
rect 9999 11577 10011 11611
rect 9953 11571 10011 11577
rect 9493 11543 9551 11549
rect 9493 11540 9505 11543
rect 9048 11512 9505 11540
rect 9493 11509 9505 11512
rect 9539 11540 9551 11543
rect 10244 11540 10272 11707
rect 10318 11704 10324 11716
rect 10376 11704 10382 11756
rect 9539 11512 10272 11540
rect 9539 11509 9551 11512
rect 9493 11503 9551 11509
rect 1104 11450 16008 11472
rect 1104 11398 5979 11450
rect 6031 11398 6043 11450
rect 6095 11398 6107 11450
rect 6159 11398 6171 11450
rect 6223 11398 10976 11450
rect 11028 11398 11040 11450
rect 11092 11398 11104 11450
rect 11156 11398 11168 11450
rect 11220 11398 16008 11450
rect 1104 11376 16008 11398
rect 1489 11339 1547 11345
rect 1489 11305 1501 11339
rect 1535 11336 1547 11339
rect 2038 11336 2044 11348
rect 1535 11308 2044 11336
rect 1535 11305 1547 11308
rect 1489 11299 1547 11305
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 3786 11336 3792 11348
rect 3747 11308 3792 11336
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 4525 11339 4583 11345
rect 4525 11305 4537 11339
rect 4571 11336 4583 11339
rect 4614 11336 4620 11348
rect 4571 11308 4620 11336
rect 4571 11305 4583 11308
rect 4525 11299 4583 11305
rect 4614 11296 4620 11308
rect 4672 11336 4678 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 4672 11308 5181 11336
rect 4672 11296 4678 11308
rect 5169 11305 5181 11308
rect 5215 11336 5227 11339
rect 5626 11336 5632 11348
rect 5215 11308 5632 11336
rect 5215 11305 5227 11308
rect 5169 11299 5227 11305
rect 5626 11296 5632 11308
rect 5684 11296 5690 11348
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 5813 11339 5871 11345
rect 5813 11336 5825 11339
rect 5776 11308 5825 11336
rect 5776 11296 5782 11308
rect 5813 11305 5825 11308
rect 5859 11305 5871 11339
rect 5813 11299 5871 11305
rect 6365 11339 6423 11345
rect 6365 11305 6377 11339
rect 6411 11336 6423 11339
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 6411 11308 6837 11336
rect 6411 11305 6423 11308
rect 6365 11299 6423 11305
rect 6825 11305 6837 11308
rect 6871 11336 6883 11339
rect 7650 11336 7656 11348
rect 6871 11308 7420 11336
rect 7611 11308 7656 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 3804 11268 3832 11296
rect 6454 11268 6460 11280
rect 3804 11240 4660 11268
rect 1854 11200 1860 11212
rect 1815 11172 1860 11200
rect 1854 11160 1860 11172
rect 1912 11160 1918 11212
rect 2665 11203 2723 11209
rect 2665 11200 2677 11203
rect 2148 11172 2677 11200
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 2148 11141 2176 11172
rect 2665 11169 2677 11172
rect 2711 11200 2723 11203
rect 2958 11200 2964 11212
rect 2711 11172 2964 11200
rect 2711 11169 2723 11172
rect 2665 11163 2723 11169
rect 2958 11160 2964 11172
rect 3016 11160 3022 11212
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4479 11172 4568 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 1949 11135 2007 11141
rect 1949 11132 1961 11135
rect 1636 11104 1961 11132
rect 1636 11092 1642 11104
rect 1949 11101 1961 11104
rect 1995 11101 2007 11135
rect 1949 11095 2007 11101
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11101 2191 11135
rect 2406 11132 2412 11144
rect 2367 11104 2412 11132
rect 2133 11095 2191 11101
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11064 4123 11067
rect 4430 11064 4436 11076
rect 4111 11036 4436 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 4430 11024 4436 11036
rect 4488 11024 4494 11076
rect 4540 11064 4568 11172
rect 4632 11141 4660 11240
rect 4724 11240 6460 11268
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4724 11064 4752 11240
rect 6454 11228 6460 11240
rect 6512 11228 6518 11280
rect 7392 11268 7420 11308
rect 7650 11296 7656 11308
rect 7708 11296 7714 11348
rect 8849 11339 8907 11345
rect 8849 11336 8861 11339
rect 8312 11308 8861 11336
rect 8312 11280 8340 11308
rect 8849 11305 8861 11308
rect 8895 11305 8907 11339
rect 8849 11299 8907 11305
rect 9677 11339 9735 11345
rect 9677 11305 9689 11339
rect 9723 11336 9735 11339
rect 9858 11336 9864 11348
rect 9723 11308 9864 11336
rect 9723 11305 9735 11308
rect 9677 11299 9735 11305
rect 9858 11296 9864 11308
rect 9916 11296 9922 11348
rect 7834 11268 7840 11280
rect 7392 11240 7840 11268
rect 7834 11228 7840 11240
rect 7892 11268 7898 11280
rect 8110 11268 8116 11280
rect 7892 11240 8116 11268
rect 7892 11228 7898 11240
rect 8110 11228 8116 11240
rect 8168 11228 8174 11280
rect 8294 11228 8300 11280
rect 8352 11268 8358 11280
rect 8352 11240 8397 11268
rect 8680 11240 8984 11268
rect 8352 11228 8358 11240
rect 5074 11200 5080 11212
rect 5035 11172 5080 11200
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 5902 11200 5908 11212
rect 5592 11172 5908 11200
rect 5592 11160 5598 11172
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 7745 11203 7803 11209
rect 6104 11172 7144 11200
rect 4982 11092 4988 11144
rect 5040 11132 5046 11144
rect 6104 11141 6132 11172
rect 6089 11135 6147 11141
rect 6089 11132 6101 11135
rect 5040 11104 6101 11132
rect 5040 11092 5046 11104
rect 6089 11101 6101 11104
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 6730 11092 6736 11144
rect 6788 11132 6794 11144
rect 7116 11141 7144 11172
rect 7745 11169 7757 11203
rect 7791 11200 7803 11203
rect 8680 11200 8708 11240
rect 7791 11172 8708 11200
rect 8757 11203 8815 11209
rect 7791 11169 7803 11172
rect 7745 11163 7803 11169
rect 8757 11169 8769 11203
rect 8803 11200 8815 11203
rect 8956 11200 8984 11240
rect 9214 11228 9220 11280
rect 9272 11268 9278 11280
rect 9876 11268 9904 11296
rect 9272 11240 9628 11268
rect 9876 11240 11376 11268
rect 9272 11228 9278 11240
rect 9401 11203 9459 11209
rect 9401 11200 9413 11203
rect 8803 11172 8892 11200
rect 8803 11169 8815 11172
rect 8757 11163 8815 11169
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6788 11104 6929 11132
rect 6788 11092 6794 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7837 11135 7895 11141
rect 7837 11132 7849 11135
rect 7147 11104 7849 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 7837 11101 7849 11104
rect 7883 11101 7895 11135
rect 7837 11095 7895 11101
rect 4540 11036 4752 11064
rect 4798 11024 4804 11076
rect 4856 11064 4862 11076
rect 4893 11067 4951 11073
rect 4893 11064 4905 11067
rect 4856 11036 4905 11064
rect 4856 11024 4862 11036
rect 4893 11033 4905 11036
rect 4939 11033 4951 11067
rect 4893 11027 4951 11033
rect 5445 11067 5503 11073
rect 5445 11033 5457 11067
rect 5491 11064 5503 11067
rect 5534 11064 5540 11076
rect 5491 11036 5540 11064
rect 5491 11033 5503 11036
rect 5445 11027 5503 11033
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 6457 11067 6515 11073
rect 6457 11033 6469 11067
rect 6503 11064 6515 11067
rect 7190 11064 7196 11076
rect 6503 11036 7196 11064
rect 6503 11033 6515 11036
rect 6457 11027 6515 11033
rect 7190 11024 7196 11036
rect 7248 11024 7254 11076
rect 8864 11064 8892 11172
rect 8956 11172 9413 11200
rect 8956 11144 8984 11172
rect 9401 11169 9413 11172
rect 9447 11169 9459 11203
rect 9600 11200 9628 11240
rect 9861 11203 9919 11209
rect 9861 11200 9873 11203
rect 9600 11172 9873 11200
rect 9401 11163 9459 11169
rect 9861 11169 9873 11172
rect 9907 11169 9919 11203
rect 9861 11163 9919 11169
rect 8938 11092 8944 11144
rect 8996 11092 9002 11144
rect 9033 11135 9091 11141
rect 9033 11101 9045 11135
rect 9079 11132 9091 11135
rect 9122 11132 9128 11144
rect 9079 11104 9128 11132
rect 9079 11101 9091 11104
rect 9033 11095 9091 11101
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9416 11132 9444 11163
rect 10042 11160 10048 11212
rect 10100 11200 10106 11212
rect 11348 11209 11376 11240
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 10100 11172 10609 11200
rect 10100 11160 10106 11172
rect 10597 11169 10609 11172
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 11600 11203 11658 11209
rect 11600 11169 11612 11203
rect 11646 11200 11658 11203
rect 12986 11200 12992 11212
rect 11646 11172 12992 11200
rect 11646 11169 11658 11172
rect 11600 11163 11658 11169
rect 12986 11160 12992 11172
rect 13044 11160 13050 11212
rect 9950 11132 9956 11144
rect 9416 11104 9956 11132
rect 9950 11092 9956 11104
rect 10008 11092 10014 11144
rect 10134 11092 10140 11144
rect 10192 11132 10198 11144
rect 10689 11135 10747 11141
rect 10689 11132 10701 11135
rect 10192 11104 10701 11132
rect 10192 11092 10198 11104
rect 10689 11101 10701 11104
rect 10735 11101 10747 11135
rect 10689 11095 10747 11101
rect 10778 11092 10784 11144
rect 10836 11132 10842 11144
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 10836 11104 10885 11132
rect 10836 11092 10842 11104
rect 10873 11101 10885 11104
rect 10919 11132 10931 11135
rect 10919 11104 11192 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 10229 11067 10287 11073
rect 8864 11036 9260 11064
rect 9232 11008 9260 11036
rect 10229 11033 10241 11067
rect 10275 11064 10287 11067
rect 11054 11064 11060 11076
rect 10275 11036 11060 11064
rect 10275 11033 10287 11036
rect 10229 11027 10287 11033
rect 11054 11024 11060 11036
rect 11112 11024 11118 11076
rect 7282 10996 7288 11008
rect 7243 10968 7288 10996
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 8389 10999 8447 11005
rect 8389 10996 8401 10999
rect 8352 10968 8401 10996
rect 8352 10956 8358 10968
rect 8389 10965 8401 10968
rect 8435 10965 8447 10999
rect 8389 10959 8447 10965
rect 9030 10956 9036 11008
rect 9088 10996 9094 11008
rect 9214 10996 9220 11008
rect 9088 10968 9220 10996
rect 9088 10956 9094 10968
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 11164 10996 11192 11104
rect 12710 10996 12716 11008
rect 11164 10968 12716 10996
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 1104 10906 16008 10928
rect 1104 10854 3480 10906
rect 3532 10854 3544 10906
rect 3596 10854 3608 10906
rect 3660 10854 3672 10906
rect 3724 10854 8478 10906
rect 8530 10854 8542 10906
rect 8594 10854 8606 10906
rect 8658 10854 8670 10906
rect 8722 10854 13475 10906
rect 13527 10854 13539 10906
rect 13591 10854 13603 10906
rect 13655 10854 13667 10906
rect 13719 10854 16008 10906
rect 1104 10832 16008 10854
rect 1489 10795 1547 10801
rect 1489 10761 1501 10795
rect 1535 10792 1547 10795
rect 1854 10792 1860 10804
rect 1535 10764 1860 10792
rect 1535 10761 1547 10764
rect 1489 10755 1547 10761
rect 1854 10752 1860 10764
rect 1912 10752 1918 10804
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4614 10792 4620 10804
rect 4019 10764 4620 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 5166 10792 5172 10804
rect 5127 10764 5172 10792
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 5868 10764 6837 10792
rect 5868 10752 5874 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 6825 10755 6883 10761
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 9858 10792 9864 10804
rect 7156 10764 9864 10792
rect 7156 10752 7162 10764
rect 3142 10724 3148 10736
rect 2792 10696 3148 10724
rect 2130 10656 2136 10668
rect 2091 10628 2136 10656
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 2792 10665 2820 10696
rect 3142 10684 3148 10696
rect 3200 10724 3206 10736
rect 3200 10696 5212 10724
rect 3200 10684 3206 10696
rect 5184 10668 5212 10696
rect 5718 10684 5724 10736
rect 5776 10724 5782 10736
rect 6365 10727 6423 10733
rect 6365 10724 6377 10727
rect 5776 10696 6377 10724
rect 5776 10684 5782 10696
rect 6365 10693 6377 10696
rect 6411 10724 6423 10727
rect 6411 10696 8432 10724
rect 6411 10693 6423 10696
rect 6365 10687 6423 10693
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10625 2835 10659
rect 2777 10619 2835 10625
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 3694 10656 3700 10668
rect 3007 10628 3700 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 2590 10548 2596 10600
rect 2648 10588 2654 10600
rect 2976 10588 3004 10619
rect 3694 10616 3700 10628
rect 3752 10616 3758 10668
rect 4430 10656 4436 10668
rect 4391 10628 4436 10656
rect 4430 10616 4436 10628
rect 4488 10616 4494 10668
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10656 4675 10659
rect 4982 10656 4988 10668
rect 4663 10628 4988 10656
rect 4663 10625 4675 10628
rect 4617 10619 4675 10625
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 5166 10616 5172 10668
rect 5224 10616 5230 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 6270 10656 6276 10668
rect 5859 10628 6276 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 6270 10616 6276 10628
rect 6328 10656 6334 10668
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 6328 10628 7389 10656
rect 6328 10616 6334 10628
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 8202 10656 8208 10668
rect 8163 10628 8208 10656
rect 7377 10619 7435 10625
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 2648 10560 3004 10588
rect 3513 10591 3571 10597
rect 2648 10548 2654 10560
rect 3513 10557 3525 10591
rect 3559 10588 3571 10591
rect 5077 10591 5135 10597
rect 5077 10588 5089 10591
rect 3559 10560 5089 10588
rect 3559 10557 3571 10560
rect 3513 10551 3571 10557
rect 5077 10557 5089 10560
rect 5123 10588 5135 10591
rect 5350 10588 5356 10600
rect 5123 10560 5356 10588
rect 5123 10557 5135 10560
rect 5077 10551 5135 10557
rect 5350 10548 5356 10560
rect 5408 10548 5414 10600
rect 5534 10588 5540 10600
rect 5495 10560 5540 10588
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 6730 10588 6736 10600
rect 5960 10560 6736 10588
rect 5960 10548 5966 10560
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10588 7251 10591
rect 7282 10588 7288 10600
rect 7239 10560 7288 10588
rect 7239 10557 7251 10560
rect 7193 10551 7251 10557
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10588 8171 10591
rect 8294 10588 8300 10600
rect 8159 10560 8300 10588
rect 8159 10557 8171 10560
rect 8113 10551 8171 10557
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 8404 10588 8432 10696
rect 8496 10665 8524 10764
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 11330 10724 11336 10736
rect 11243 10696 11336 10724
rect 11330 10684 11336 10696
rect 11388 10724 11394 10736
rect 11388 10696 12020 10724
rect 11388 10684 11394 10696
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 9916 10628 9965 10656
rect 9916 10616 9922 10628
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11992 10665 12020 10696
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 11112 10628 11897 10656
rect 11112 10616 11118 10628
rect 11885 10625 11897 10628
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12710 10616 12716 10668
rect 12768 10656 12774 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12768 10628 13001 10656
rect 12768 10616 12774 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 9030 10588 9036 10600
rect 8404 10560 9036 10588
rect 9030 10548 9036 10560
rect 9088 10548 9094 10600
rect 10220 10591 10278 10597
rect 10220 10557 10232 10591
rect 10266 10588 10278 10591
rect 10778 10588 10784 10600
rect 10266 10560 10784 10588
rect 10266 10557 10278 10560
rect 10220 10551 10278 10557
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10520 1915 10523
rect 2685 10523 2743 10529
rect 1903 10492 2360 10520
rect 1903 10489 1915 10492
rect 1857 10483 1915 10489
rect 1949 10455 2007 10461
rect 1949 10421 1961 10455
rect 1995 10452 2007 10455
rect 2222 10452 2228 10464
rect 1995 10424 2228 10452
rect 1995 10421 2007 10424
rect 1949 10415 2007 10421
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 2332 10461 2360 10492
rect 2685 10489 2697 10523
rect 2731 10520 2743 10523
rect 3326 10520 3332 10532
rect 2731 10492 3332 10520
rect 2731 10489 2743 10492
rect 2685 10483 2743 10489
rect 3326 10480 3332 10492
rect 3384 10480 3390 10532
rect 3605 10523 3663 10529
rect 3605 10489 3617 10523
rect 3651 10520 3663 10523
rect 4246 10520 4252 10532
rect 3651 10492 4252 10520
rect 3651 10489 3663 10492
rect 3605 10483 3663 10489
rect 4246 10480 4252 10492
rect 4304 10480 4310 10532
rect 4614 10480 4620 10532
rect 4672 10520 4678 10532
rect 5629 10523 5687 10529
rect 5629 10520 5641 10523
rect 4672 10492 5641 10520
rect 4672 10480 4678 10492
rect 5629 10489 5641 10492
rect 5675 10489 5687 10523
rect 6914 10520 6920 10532
rect 5629 10483 5687 10489
rect 6012 10492 6920 10520
rect 2317 10455 2375 10461
rect 2317 10421 2329 10455
rect 2363 10421 2375 10455
rect 2317 10415 2375 10421
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 3145 10455 3203 10461
rect 3145 10452 3157 10455
rect 3108 10424 3157 10452
rect 3108 10412 3114 10424
rect 3145 10421 3157 10424
rect 3191 10421 3203 10455
rect 3145 10415 3203 10421
rect 4341 10455 4399 10461
rect 4341 10421 4353 10455
rect 4387 10452 4399 10455
rect 4893 10455 4951 10461
rect 4893 10452 4905 10455
rect 4387 10424 4905 10452
rect 4387 10421 4399 10424
rect 4341 10415 4399 10421
rect 4893 10421 4905 10424
rect 4939 10452 4951 10455
rect 6012 10452 6040 10492
rect 6914 10480 6920 10492
rect 6972 10520 6978 10532
rect 8748 10523 8806 10529
rect 6972 10492 8432 10520
rect 6972 10480 6978 10492
rect 4939 10424 6040 10452
rect 6089 10455 6147 10461
rect 4939 10421 4951 10424
rect 4893 10415 4951 10421
rect 6089 10421 6101 10455
rect 6135 10452 6147 10455
rect 6454 10452 6460 10464
rect 6135 10424 6460 10452
rect 6135 10421 6147 10424
rect 6089 10415 6147 10421
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10452 6607 10455
rect 6730 10452 6736 10464
rect 6595 10424 6736 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 7190 10412 7196 10464
rect 7248 10452 7254 10464
rect 7285 10455 7343 10461
rect 7285 10452 7297 10455
rect 7248 10424 7297 10452
rect 7248 10412 7254 10424
rect 7285 10421 7297 10424
rect 7331 10421 7343 10455
rect 7285 10415 7343 10421
rect 7374 10412 7380 10464
rect 7432 10452 7438 10464
rect 7653 10455 7711 10461
rect 7653 10452 7665 10455
rect 7432 10424 7665 10452
rect 7432 10412 7438 10424
rect 7653 10421 7665 10424
rect 7699 10421 7711 10455
rect 7653 10415 7711 10421
rect 8021 10455 8079 10461
rect 8021 10421 8033 10455
rect 8067 10452 8079 10455
rect 8294 10452 8300 10464
rect 8067 10424 8300 10452
rect 8067 10421 8079 10424
rect 8021 10415 8079 10421
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 8404 10452 8432 10492
rect 8748 10489 8760 10523
rect 8794 10520 8806 10523
rect 9122 10520 9128 10532
rect 8794 10492 9128 10520
rect 8794 10489 8806 10492
rect 8748 10483 8806 10489
rect 9122 10480 9128 10492
rect 9180 10480 9186 10532
rect 11793 10523 11851 10529
rect 11793 10489 11805 10523
rect 11839 10520 11851 10523
rect 11839 10492 12480 10520
rect 11839 10489 11851 10492
rect 11793 10483 11851 10489
rect 8846 10452 8852 10464
rect 8404 10424 8852 10452
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 9858 10452 9864 10464
rect 9819 10424 9864 10452
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 11422 10452 11428 10464
rect 11383 10424 11428 10452
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 12452 10461 12480 10492
rect 12618 10480 12624 10532
rect 12676 10520 12682 10532
rect 12897 10523 12955 10529
rect 12897 10520 12909 10523
rect 12676 10492 12909 10520
rect 12676 10480 12682 10492
rect 12897 10489 12909 10492
rect 12943 10489 12955 10523
rect 12897 10483 12955 10489
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10421 12495 10455
rect 12802 10452 12808 10464
rect 12763 10424 12808 10452
rect 12437 10415 12495 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13265 10455 13323 10461
rect 13265 10421 13277 10455
rect 13311 10452 13323 10455
rect 13354 10452 13360 10464
rect 13311 10424 13360 10452
rect 13311 10421 13323 10424
rect 13265 10415 13323 10421
rect 13354 10412 13360 10424
rect 13412 10412 13418 10464
rect 1104 10362 16008 10384
rect 1104 10310 5979 10362
rect 6031 10310 6043 10362
rect 6095 10310 6107 10362
rect 6159 10310 6171 10362
rect 6223 10310 10976 10362
rect 11028 10310 11040 10362
rect 11092 10310 11104 10362
rect 11156 10310 11168 10362
rect 11220 10310 16008 10362
rect 1104 10288 16008 10310
rect 2958 10248 2964 10260
rect 2919 10220 2964 10248
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 3605 10251 3663 10257
rect 3605 10217 3617 10251
rect 3651 10248 3663 10251
rect 4249 10251 4307 10257
rect 4249 10248 4261 10251
rect 3651 10220 4261 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 4249 10217 4261 10220
rect 4295 10217 4307 10251
rect 4249 10211 4307 10217
rect 4522 10208 4528 10260
rect 4580 10248 4586 10260
rect 4617 10251 4675 10257
rect 4617 10248 4629 10251
rect 4580 10220 4629 10248
rect 4580 10208 4586 10220
rect 4617 10217 4629 10220
rect 4663 10248 4675 10251
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 4663 10220 6837 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 6825 10217 6837 10220
rect 6871 10248 6883 10251
rect 6914 10248 6920 10260
rect 6871 10220 6920 10248
rect 6871 10217 6883 10220
rect 6825 10211 6883 10217
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7650 10208 7656 10260
rect 7708 10248 7714 10260
rect 8754 10248 8760 10260
rect 7708 10220 8760 10248
rect 7708 10208 7714 10220
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 12161 10251 12219 10257
rect 12161 10217 12173 10251
rect 12207 10248 12219 10251
rect 12618 10248 12624 10260
rect 12207 10220 12624 10248
rect 12207 10217 12219 10220
rect 12161 10211 12219 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 12989 10251 13047 10257
rect 12989 10248 13001 10251
rect 12860 10220 13001 10248
rect 12860 10208 12866 10220
rect 12989 10217 13001 10220
rect 13035 10217 13047 10251
rect 13354 10248 13360 10260
rect 13315 10220 13360 10248
rect 12989 10211 13047 10217
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 13449 10251 13507 10257
rect 13449 10217 13461 10251
rect 13495 10248 13507 10251
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 13495 10220 14289 10248
rect 13495 10217 13507 10220
rect 13449 10211 13507 10217
rect 14277 10217 14289 10220
rect 14323 10248 14335 10251
rect 16206 10248 16212 10260
rect 14323 10220 16212 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 2406 10180 2412 10192
rect 1596 10152 2412 10180
rect 1596 10121 1624 10152
rect 2406 10140 2412 10152
rect 2464 10140 2470 10192
rect 3513 10183 3571 10189
rect 3513 10149 3525 10183
rect 3559 10180 3571 10183
rect 3878 10180 3884 10192
rect 3559 10152 3884 10180
rect 3559 10149 3571 10152
rect 3513 10143 3571 10149
rect 3878 10140 3884 10152
rect 3936 10180 3942 10192
rect 4157 10183 4215 10189
rect 4157 10180 4169 10183
rect 3936 10152 4169 10180
rect 3936 10140 3942 10152
rect 4157 10149 4169 10152
rect 4203 10180 4215 10183
rect 4203 10152 5488 10180
rect 4203 10149 4215 10152
rect 4157 10143 4215 10149
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 1848 10115 1906 10121
rect 1848 10081 1860 10115
rect 1894 10112 1906 10115
rect 2130 10112 2136 10124
rect 1894 10084 2136 10112
rect 1894 10081 1906 10084
rect 1848 10075 1906 10081
rect 2130 10072 2136 10084
rect 2188 10072 2194 10124
rect 4338 10072 4344 10124
rect 4396 10112 4402 10124
rect 4709 10115 4767 10121
rect 4709 10112 4721 10115
rect 4396 10084 4721 10112
rect 4396 10072 4402 10084
rect 4709 10081 4721 10084
rect 4755 10081 4767 10115
rect 4709 10075 4767 10081
rect 3786 10044 3792 10056
rect 3747 10016 3792 10044
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 2958 9868 2964 9920
rect 3016 9908 3022 9920
rect 3145 9911 3203 9917
rect 3145 9908 3157 9911
rect 3016 9880 3157 9908
rect 3016 9868 3022 9880
rect 3145 9877 3157 9880
rect 3191 9877 3203 9911
rect 4724 9908 4752 10075
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 5353 10115 5411 10121
rect 5353 10112 5365 10115
rect 4856 10084 5365 10112
rect 4856 10072 4862 10084
rect 5353 10081 5365 10084
rect 5399 10081 5411 10115
rect 5460 10112 5488 10152
rect 5534 10140 5540 10192
rect 5592 10189 5598 10192
rect 5592 10183 5656 10189
rect 5592 10149 5610 10183
rect 5644 10149 5656 10183
rect 5592 10143 5656 10149
rect 5592 10140 5598 10143
rect 6730 10140 6736 10192
rect 6788 10180 6794 10192
rect 9398 10180 9404 10192
rect 6788 10152 9404 10180
rect 6788 10140 6794 10152
rect 9398 10140 9404 10152
rect 9456 10140 9462 10192
rect 10588 10183 10646 10189
rect 10588 10149 10600 10183
rect 10634 10180 10646 10183
rect 11330 10180 11336 10192
rect 10634 10152 11336 10180
rect 10634 10149 10646 10152
rect 10588 10143 10646 10149
rect 11330 10140 11336 10152
rect 11388 10140 11394 10192
rect 11974 10140 11980 10192
rect 12032 10180 12038 10192
rect 12434 10180 12440 10192
rect 12032 10152 12440 10180
rect 12032 10140 12038 10152
rect 12434 10140 12440 10152
rect 12492 10180 12498 10192
rect 14001 10183 14059 10189
rect 14001 10180 14013 10183
rect 12492 10152 14013 10180
rect 12492 10140 12498 10152
rect 7101 10115 7159 10121
rect 5460 10084 6408 10112
rect 5353 10075 5411 10081
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10013 4951 10047
rect 6380 10044 6408 10084
rect 7101 10081 7113 10115
rect 7147 10112 7159 10115
rect 7190 10112 7196 10124
rect 7147 10084 7196 10112
rect 7147 10081 7159 10084
rect 7101 10075 7159 10081
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 9490 10112 9496 10124
rect 7300 10084 9496 10112
rect 7300 10044 7328 10084
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 12636 10121 12664 10152
rect 14001 10149 14013 10152
rect 14047 10149 14059 10183
rect 14001 10143 14059 10149
rect 10321 10115 10379 10121
rect 10321 10112 10333 10115
rect 10008 10084 10333 10112
rect 10008 10072 10014 10084
rect 10321 10081 10333 10084
rect 10367 10081 10379 10115
rect 12529 10115 12587 10121
rect 12529 10112 12541 10115
rect 10321 10075 10379 10081
rect 10428 10084 12541 10112
rect 6380 10016 7328 10044
rect 4893 10007 4951 10013
rect 4908 9976 4936 10007
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 10428 10044 10456 10084
rect 12529 10081 12541 10084
rect 12575 10081 12587 10115
rect 12529 10075 12587 10081
rect 12621 10115 12679 10121
rect 12621 10081 12633 10115
rect 12667 10081 12679 10115
rect 12621 10075 12679 10081
rect 7524 10016 10456 10044
rect 7524 10004 7530 10016
rect 4908 9948 5396 9976
rect 5368 9920 5396 9948
rect 6914 9936 6920 9988
rect 6972 9976 6978 9988
rect 8110 9976 8116 9988
rect 6972 9948 8116 9976
rect 6972 9936 6978 9948
rect 8110 9936 8116 9948
rect 8168 9936 8174 9988
rect 8754 9936 8760 9988
rect 8812 9976 8818 9988
rect 9950 9976 9956 9988
rect 8812 9948 9956 9976
rect 8812 9936 8818 9948
rect 9950 9936 9956 9948
rect 10008 9936 10014 9988
rect 12544 9976 12572 10075
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10044 12771 10047
rect 12986 10044 12992 10056
rect 12759 10016 12992 10044
rect 12759 10013 12771 10016
rect 12713 10007 12771 10013
rect 12986 10004 12992 10016
rect 13044 10044 13050 10056
rect 13541 10047 13599 10053
rect 13541 10044 13553 10047
rect 13044 10016 13553 10044
rect 13044 10004 13050 10016
rect 13541 10013 13553 10016
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 12802 9976 12808 9988
rect 12544 9948 12808 9976
rect 12802 9936 12808 9948
rect 12860 9976 12866 9988
rect 13817 9979 13875 9985
rect 13817 9976 13829 9979
rect 12860 9948 13829 9976
rect 12860 9936 12866 9948
rect 13817 9945 13829 9948
rect 13863 9945 13875 9979
rect 13817 9939 13875 9945
rect 5074 9908 5080 9920
rect 4724 9880 5080 9908
rect 3145 9871 3203 9877
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5350 9868 5356 9920
rect 5408 9908 5414 9920
rect 6733 9911 6791 9917
rect 6733 9908 6745 9911
rect 5408 9880 6745 9908
rect 5408 9868 5414 9880
rect 6733 9877 6745 9880
rect 6779 9877 6791 9911
rect 6733 9871 6791 9877
rect 7006 9868 7012 9920
rect 7064 9908 7070 9920
rect 7558 9908 7564 9920
rect 7064 9880 7564 9908
rect 7064 9868 7070 9880
rect 7558 9868 7564 9880
rect 7616 9908 7622 9920
rect 8389 9911 8447 9917
rect 8389 9908 8401 9911
rect 7616 9880 8401 9908
rect 7616 9868 7622 9880
rect 8389 9877 8401 9880
rect 8435 9877 8447 9911
rect 8389 9871 8447 9877
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 11701 9911 11759 9917
rect 11701 9908 11713 9911
rect 9180 9880 11713 9908
rect 9180 9868 9186 9880
rect 11701 9877 11713 9880
rect 11747 9877 11759 9911
rect 11701 9871 11759 9877
rect 1104 9818 16008 9840
rect 1104 9766 3480 9818
rect 3532 9766 3544 9818
rect 3596 9766 3608 9818
rect 3660 9766 3672 9818
rect 3724 9766 8478 9818
rect 8530 9766 8542 9818
rect 8594 9766 8606 9818
rect 8658 9766 8670 9818
rect 8722 9766 13475 9818
rect 13527 9766 13539 9818
rect 13591 9766 13603 9818
rect 13655 9766 13667 9818
rect 13719 9766 16008 9818
rect 1104 9744 16008 9766
rect 5092 9676 6040 9704
rect 3786 9596 3792 9648
rect 3844 9636 3850 9648
rect 5092 9636 5120 9676
rect 3844 9608 5120 9636
rect 6012 9636 6040 9676
rect 6840 9676 7788 9704
rect 6457 9639 6515 9645
rect 6457 9636 6469 9639
rect 6012 9608 6469 9636
rect 3844 9596 3850 9608
rect 6457 9605 6469 9608
rect 6503 9605 6515 9639
rect 6457 9599 6515 9605
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6840 9636 6868 9676
rect 6604 9608 6868 9636
rect 7760 9636 7788 9676
rect 8110 9664 8116 9716
rect 8168 9704 8174 9716
rect 9766 9704 9772 9716
rect 8168 9676 9772 9704
rect 8168 9664 8174 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 11606 9664 11612 9716
rect 11664 9704 11670 9716
rect 11885 9707 11943 9713
rect 11885 9704 11897 9707
rect 11664 9676 11897 9704
rect 11664 9664 11670 9676
rect 11885 9673 11897 9676
rect 11931 9673 11943 9707
rect 11885 9667 11943 9673
rect 7760 9608 7880 9636
rect 6604 9596 6610 9608
rect 3694 9568 3700 9580
rect 3655 9540 3700 9568
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9537 4951 9571
rect 7852 9568 7880 9608
rect 8294 9596 8300 9648
rect 8352 9636 8358 9648
rect 8481 9639 8539 9645
rect 8481 9636 8493 9639
rect 8352 9608 8493 9636
rect 8352 9596 8358 9608
rect 8481 9605 8493 9608
rect 8527 9605 8539 9639
rect 8481 9599 8539 9605
rect 8754 9596 8760 9648
rect 8812 9636 8818 9648
rect 9214 9636 9220 9648
rect 8812 9608 9220 9636
rect 8812 9596 8818 9608
rect 9214 9596 9220 9608
rect 9272 9596 9278 9648
rect 10042 9636 10048 9648
rect 10003 9608 10048 9636
rect 10042 9596 10048 9608
rect 10100 9596 10106 9648
rect 10873 9639 10931 9645
rect 10873 9636 10885 9639
rect 10428 9608 10885 9636
rect 4893 9531 4951 9537
rect 6104 9540 6960 9568
rect 7852 9540 8432 9568
rect 1486 9500 1492 9512
rect 1447 9472 1492 9500
rect 1486 9460 1492 9472
rect 1544 9460 1550 9512
rect 2038 9500 2044 9512
rect 1999 9472 2044 9500
rect 2038 9460 2044 9472
rect 2096 9460 2102 9512
rect 3142 9460 3148 9512
rect 3200 9500 3206 9512
rect 3513 9503 3571 9509
rect 3513 9500 3525 9503
rect 3200 9472 3525 9500
rect 3200 9460 3206 9472
rect 3513 9469 3525 9472
rect 3559 9469 3571 9503
rect 3513 9463 3571 9469
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9500 4215 9503
rect 4246 9500 4252 9512
rect 4203 9472 4252 9500
rect 4203 9469 4215 9472
rect 4157 9463 4215 9469
rect 4246 9460 4252 9472
rect 4304 9500 4310 9512
rect 4798 9500 4804 9512
rect 4304 9472 4804 9500
rect 4304 9460 4310 9472
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 1762 9432 1768 9444
rect 1723 9404 1768 9432
rect 1762 9392 1768 9404
rect 1820 9392 1826 9444
rect 2308 9435 2366 9441
rect 2308 9401 2320 9435
rect 2354 9432 2366 9435
rect 2590 9432 2596 9444
rect 2354 9404 2596 9432
rect 2354 9401 2366 9404
rect 2308 9395 2366 9401
rect 2590 9392 2596 9404
rect 2648 9392 2654 9444
rect 4908 9432 4936 9531
rect 4982 9460 4988 9512
rect 5040 9500 5046 9512
rect 5350 9509 5356 9512
rect 5077 9503 5135 9509
rect 5077 9500 5089 9503
rect 5040 9472 5089 9500
rect 5040 9460 5046 9472
rect 5077 9469 5089 9472
rect 5123 9469 5135 9503
rect 5344 9500 5356 9509
rect 5311 9472 5356 9500
rect 5077 9463 5135 9469
rect 5344 9463 5356 9472
rect 5350 9460 5356 9463
rect 5408 9460 5414 9512
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 6104 9500 6132 9540
rect 5684 9472 6132 9500
rect 6641 9503 6699 9509
rect 5684 9460 5690 9472
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6687 9472 6837 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 6932 9500 6960 9540
rect 6932 9472 8248 9500
rect 6825 9463 6883 9469
rect 7098 9441 7104 9444
rect 7092 9432 7104 9441
rect 4908 9404 7104 9432
rect 7092 9395 7104 9404
rect 7098 9392 7104 9395
rect 7156 9392 7162 9444
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 3421 9367 3479 9373
rect 3421 9364 3433 9367
rect 2188 9336 3433 9364
rect 2188 9324 2194 9336
rect 3421 9333 3433 9336
rect 3467 9333 3479 9367
rect 4246 9364 4252 9376
rect 4207 9336 4252 9364
rect 3421 9327 3479 9333
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 4614 9364 4620 9376
rect 4575 9336 4620 9364
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 4709 9367 4767 9373
rect 4709 9333 4721 9367
rect 4755 9364 4767 9367
rect 6362 9364 6368 9376
rect 4755 9336 6368 9364
rect 4755 9333 4767 9336
rect 4709 9327 4767 9333
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 6641 9367 6699 9373
rect 6641 9333 6653 9367
rect 6687 9364 6699 9367
rect 7650 9364 7656 9376
rect 6687 9336 7656 9364
rect 6687 9333 6699 9336
rect 6641 9327 6699 9333
rect 7650 9324 7656 9336
rect 7708 9364 7714 9376
rect 8110 9364 8116 9376
rect 7708 9336 8116 9364
rect 7708 9324 7714 9336
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 8220 9373 8248 9472
rect 8404 9444 8432 9540
rect 8846 9528 8852 9580
rect 8904 9528 8910 9580
rect 9122 9568 9128 9580
rect 9083 9540 9128 9568
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 10318 9528 10324 9580
rect 10376 9568 10382 9580
rect 10428 9568 10456 9608
rect 10873 9605 10885 9608
rect 10919 9605 10931 9639
rect 10873 9599 10931 9605
rect 10686 9568 10692 9580
rect 10376 9540 10456 9568
rect 10647 9540 10692 9568
rect 10376 9528 10382 9540
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9568 11575 9571
rect 12710 9568 12716 9580
rect 11563 9540 12716 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 15286 9568 15292 9580
rect 15247 9540 15292 9568
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 8864 9500 8892 9528
rect 8941 9503 8999 9509
rect 8941 9500 8953 9503
rect 8864 9472 8953 9500
rect 8941 9469 8953 9472
rect 8987 9500 8999 9503
rect 9214 9500 9220 9512
rect 8987 9472 9220 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 9214 9460 9220 9472
rect 9272 9500 9278 9512
rect 9309 9503 9367 9509
rect 9309 9500 9321 9503
rect 9272 9472 9321 9500
rect 9272 9460 9278 9472
rect 9309 9469 9321 9472
rect 9355 9469 9367 9503
rect 9309 9463 9367 9469
rect 9490 9460 9496 9512
rect 9548 9500 9554 9512
rect 11241 9503 11299 9509
rect 9548 9472 9996 9500
rect 9548 9460 9554 9472
rect 8386 9432 8392 9444
rect 8299 9404 8392 9432
rect 8386 9392 8392 9404
rect 8444 9432 8450 9444
rect 9674 9432 9680 9444
rect 8444 9404 9680 9432
rect 8444 9392 8450 9404
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 8205 9367 8263 9373
rect 8205 9333 8217 9367
rect 8251 9333 8263 9367
rect 8205 9327 8263 9333
rect 8849 9367 8907 9373
rect 8849 9333 8861 9367
rect 8895 9364 8907 9367
rect 9398 9364 9404 9376
rect 8895 9336 9404 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9398 9324 9404 9336
rect 9456 9364 9462 9376
rect 9493 9367 9551 9373
rect 9493 9364 9505 9367
rect 9456 9336 9505 9364
rect 9456 9324 9462 9336
rect 9493 9333 9505 9336
rect 9539 9333 9551 9367
rect 9766 9364 9772 9376
rect 9727 9336 9772 9364
rect 9493 9327 9551 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 9968 9373 9996 9472
rect 11241 9469 11253 9503
rect 11287 9500 11299 9503
rect 11606 9500 11612 9512
rect 11287 9472 11612 9500
rect 11287 9469 11299 9472
rect 11241 9463 11299 9469
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 12066 9460 12072 9512
rect 12124 9500 12130 9512
rect 13078 9500 13084 9512
rect 12124 9472 13084 9500
rect 12124 9460 12130 9472
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 15010 9500 15016 9512
rect 14844 9472 15016 9500
rect 11330 9432 11336 9444
rect 11291 9404 11336 9432
rect 11330 9392 11336 9404
rect 11388 9392 11394 9444
rect 11422 9392 11428 9444
rect 11480 9432 11486 9444
rect 11701 9435 11759 9441
rect 11701 9432 11713 9435
rect 11480 9404 11713 9432
rect 11480 9392 11486 9404
rect 11701 9401 11713 9404
rect 11747 9401 11759 9435
rect 11701 9395 11759 9401
rect 9953 9367 10011 9373
rect 9953 9333 9965 9367
rect 9999 9364 10011 9367
rect 10042 9364 10048 9376
rect 9999 9336 10048 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 10226 9324 10232 9376
rect 10284 9364 10290 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 10284 9336 10425 9364
rect 10284 9324 10290 9336
rect 10413 9333 10425 9336
rect 10459 9333 10471 9367
rect 10413 9327 10471 9333
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 10560 9336 10605 9364
rect 10560 9324 10566 9336
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 14844 9373 14872 9472
rect 15010 9460 15016 9472
rect 15068 9460 15074 9512
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 13872 9336 14841 9364
rect 13872 9324 13878 9336
rect 14829 9333 14841 9336
rect 14875 9333 14887 9367
rect 14829 9327 14887 9333
rect 1104 9274 16008 9296
rect 1104 9222 5979 9274
rect 6031 9222 6043 9274
rect 6095 9222 6107 9274
rect 6159 9222 6171 9274
rect 6223 9222 10976 9274
rect 11028 9222 11040 9274
rect 11092 9222 11104 9274
rect 11156 9222 11168 9274
rect 11220 9222 16008 9274
rect 1104 9200 16008 9222
rect 1489 9163 1547 9169
rect 1489 9129 1501 9163
rect 1535 9160 1547 9163
rect 1578 9160 1584 9172
rect 1535 9132 1584 9160
rect 1535 9129 1547 9132
rect 1489 9123 1547 9129
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 2222 9120 2228 9172
rect 2280 9160 2286 9172
rect 2317 9163 2375 9169
rect 2317 9160 2329 9163
rect 2280 9132 2329 9160
rect 2280 9120 2286 9132
rect 2317 9129 2329 9132
rect 2363 9129 2375 9163
rect 3142 9160 3148 9172
rect 3103 9132 3148 9160
rect 2317 9123 2375 9129
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 4246 9160 4252 9172
rect 3559 9132 4252 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4709 9163 4767 9169
rect 4709 9160 4721 9163
rect 4396 9132 4721 9160
rect 4396 9120 4402 9132
rect 4709 9129 4721 9132
rect 4755 9129 4767 9163
rect 4709 9123 4767 9129
rect 5169 9163 5227 9169
rect 5169 9129 5181 9163
rect 5215 9160 5227 9163
rect 5537 9163 5595 9169
rect 5537 9160 5549 9163
rect 5215 9132 5549 9160
rect 5215 9129 5227 9132
rect 5169 9123 5227 9129
rect 5537 9129 5549 9132
rect 5583 9129 5595 9163
rect 5537 9123 5595 9129
rect 6825 9163 6883 9169
rect 6825 9129 6837 9163
rect 6871 9160 6883 9163
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 6871 9132 7297 9160
rect 6871 9129 6883 9132
rect 6825 9123 6883 9129
rect 7285 9129 7297 9132
rect 7331 9129 7343 9163
rect 7285 9123 7343 9129
rect 7653 9163 7711 9169
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 8386 9160 8392 9172
rect 7699 9132 8392 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 10045 9163 10103 9169
rect 10045 9129 10057 9163
rect 10091 9160 10103 9163
rect 10134 9160 10140 9172
rect 10091 9132 10140 9160
rect 10091 9129 10103 9132
rect 10045 9123 10103 9129
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10318 9120 10324 9172
rect 10376 9160 10382 9172
rect 10413 9163 10471 9169
rect 10413 9160 10425 9163
rect 10376 9132 10425 9160
rect 10376 9120 10382 9132
rect 10413 9129 10425 9132
rect 10459 9129 10471 9163
rect 11241 9163 11299 9169
rect 11241 9160 11253 9163
rect 10413 9123 10471 9129
rect 10520 9132 11253 9160
rect 1949 9095 2007 9101
rect 1949 9061 1961 9095
rect 1995 9092 2007 9095
rect 2866 9092 2872 9104
rect 1995 9064 2872 9092
rect 1995 9061 2007 9064
rect 1949 9055 2007 9061
rect 2866 9052 2872 9064
rect 2924 9052 2930 9104
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 4065 9095 4123 9101
rect 4065 9092 4077 9095
rect 3384 9064 4077 9092
rect 3384 9052 3390 9064
rect 4065 9061 4077 9064
rect 4111 9061 4123 9095
rect 4065 9055 4123 9061
rect 5077 9095 5135 9101
rect 5077 9061 5089 9095
rect 5123 9092 5135 9095
rect 6730 9092 6736 9104
rect 5123 9064 6736 9092
rect 5123 9061 5135 9064
rect 5077 9055 5135 9061
rect 6730 9052 6736 9064
rect 6788 9052 6794 9104
rect 6917 9095 6975 9101
rect 6917 9061 6929 9095
rect 6963 9092 6975 9095
rect 7374 9092 7380 9104
rect 6963 9064 7380 9092
rect 6963 9061 6975 9064
rect 6917 9055 6975 9061
rect 7374 9052 7380 9064
rect 7432 9052 7438 9104
rect 9490 9092 9496 9104
rect 7576 9064 9496 9092
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 8993 1915 9027
rect 2682 9024 2688 9036
rect 2643 8996 2688 9024
rect 1857 8987 1915 8993
rect 1872 8888 1900 8987
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 5442 9024 5448 9036
rect 2832 8996 2877 9024
rect 3712 8996 5448 9024
rect 2832 8984 2838 8996
rect 2130 8956 2136 8968
rect 2091 8928 2136 8956
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 3712 8965 3740 8996
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 5905 9027 5963 9033
rect 5905 9024 5917 9027
rect 5592 8996 5917 9024
rect 5592 8984 5598 8996
rect 5905 8993 5917 8996
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 6362 8984 6368 9036
rect 6420 9024 6426 9036
rect 7576 9024 7604 9064
rect 9490 9052 9496 9064
rect 9548 9052 9554 9104
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 10520 9092 10548 9132
rect 11241 9129 11253 9132
rect 11287 9160 11299 9163
rect 12250 9160 12256 9172
rect 11287 9132 12256 9160
rect 11287 9129 11299 9132
rect 11241 9123 11299 9129
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 12894 9160 12900 9172
rect 12584 9132 12900 9160
rect 12584 9120 12590 9132
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 13044 9132 13093 9160
rect 13044 9120 13050 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13081 9123 13139 9129
rect 9824 9064 10548 9092
rect 9824 9052 9830 9064
rect 10686 9052 10692 9104
rect 10744 9092 10750 9104
rect 13004 9092 13032 9120
rect 10744 9064 13032 9092
rect 10744 9052 10750 9064
rect 8202 9024 8208 9036
rect 6420 8996 7604 9024
rect 7944 8996 8208 9024
rect 6420 8984 6426 8996
rect 2915 8959 2973 8965
rect 2915 8956 2927 8959
rect 2648 8928 2927 8956
rect 2648 8916 2654 8928
rect 2915 8925 2927 8928
rect 2961 8925 2973 8959
rect 2915 8919 2973 8925
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8925 3663 8959
rect 3605 8919 3663 8925
rect 3697 8959 3755 8965
rect 3697 8925 3709 8959
rect 3743 8925 3755 8959
rect 3697 8919 3755 8925
rect 5353 8959 5411 8965
rect 5353 8925 5365 8959
rect 5399 8956 5411 8959
rect 5718 8956 5724 8968
rect 5399 8928 5724 8956
rect 5399 8925 5411 8928
rect 5353 8919 5411 8925
rect 3050 8888 3056 8900
rect 1872 8860 3056 8888
rect 3050 8848 3056 8860
rect 3108 8848 3114 8900
rect 3620 8888 3648 8919
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 5810 8916 5816 8968
rect 5868 8956 5874 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5868 8928 6009 8956
rect 5868 8916 5874 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 6178 8956 6184 8968
rect 6139 8928 6184 8956
rect 5997 8919 6055 8925
rect 6178 8916 6184 8928
rect 6236 8916 6242 8968
rect 7098 8956 7104 8968
rect 7011 8928 7104 8956
rect 7098 8916 7104 8928
rect 7156 8956 7162 8968
rect 7742 8956 7748 8968
rect 7156 8928 7236 8956
rect 7703 8928 7748 8956
rect 7156 8916 7162 8928
rect 6457 8891 6515 8897
rect 6457 8888 6469 8891
rect 3620 8860 6469 8888
rect 6457 8857 6469 8860
rect 6503 8857 6515 8891
rect 6457 8851 6515 8857
rect 2682 8780 2688 8832
rect 2740 8820 2746 8832
rect 4246 8820 4252 8832
rect 2740 8792 4252 8820
rect 2740 8780 2746 8792
rect 4246 8780 4252 8792
rect 4304 8820 4310 8832
rect 4341 8823 4399 8829
rect 4341 8820 4353 8823
rect 4304 8792 4353 8820
rect 4304 8780 4310 8792
rect 4341 8789 4353 8792
rect 4387 8789 4399 8823
rect 4522 8820 4528 8832
rect 4483 8792 4528 8820
rect 4341 8783 4399 8789
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 4614 8780 4620 8832
rect 4672 8820 4678 8832
rect 6546 8820 6552 8832
rect 4672 8792 6552 8820
rect 4672 8780 4678 8792
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 7208 8820 7236 8928
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 7944 8965 7972 8996
rect 8202 8984 8208 8996
rect 8260 9024 8266 9036
rect 8380 9027 8438 9033
rect 8380 9024 8392 9027
rect 8260 8996 8392 9024
rect 8260 8984 8266 8996
rect 8380 8993 8392 8996
rect 8426 9024 8438 9027
rect 9858 9024 9864 9036
rect 8426 8996 9864 9024
rect 8426 8993 8438 8996
rect 8380 8987 8438 8993
rect 9858 8984 9864 8996
rect 9916 9024 9922 9036
rect 10134 9024 10140 9036
rect 9916 8996 10140 9024
rect 9916 8984 9922 8996
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 10551 8996 10916 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 8110 8956 8116 8968
rect 8071 8928 8116 8956
rect 7929 8919 7987 8925
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8956 9735 8959
rect 10410 8956 10416 8968
rect 9723 8928 10416 8956
rect 9723 8925 9735 8928
rect 9677 8919 9735 8925
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10686 8956 10692 8968
rect 10647 8928 10692 8956
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 10888 8897 10916 8996
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 11296 8996 11345 9024
rect 11296 8984 11302 8996
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 11968 9027 12026 9033
rect 11968 9024 11980 9027
rect 11333 8987 11391 8993
rect 11532 8996 11980 9024
rect 11532 8965 11560 8996
rect 11968 8993 11980 8996
rect 12014 9024 12026 9027
rect 12710 9024 12716 9036
rect 12014 8996 12716 9024
rect 12014 8993 12026 8996
rect 11968 8987 12026 8993
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8925 11759 8959
rect 11701 8919 11759 8925
rect 10873 8891 10931 8897
rect 10873 8857 10885 8891
rect 10919 8857 10931 8891
rect 10873 8851 10931 8857
rect 11330 8848 11336 8900
rect 11388 8888 11394 8900
rect 11716 8888 11744 8919
rect 11388 8860 11744 8888
rect 11388 8848 11394 8860
rect 9493 8823 9551 8829
rect 9493 8820 9505 8823
rect 7208 8792 9505 8820
rect 9493 8789 9505 8792
rect 9539 8789 9551 8823
rect 9493 8783 9551 8789
rect 10134 8780 10140 8832
rect 10192 8820 10198 8832
rect 12986 8820 12992 8832
rect 10192 8792 12992 8820
rect 10192 8780 10198 8792
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 1104 8730 16008 8752
rect 1104 8678 3480 8730
rect 3532 8678 3544 8730
rect 3596 8678 3608 8730
rect 3660 8678 3672 8730
rect 3724 8678 8478 8730
rect 8530 8678 8542 8730
rect 8594 8678 8606 8730
rect 8658 8678 8670 8730
rect 8722 8678 13475 8730
rect 13527 8678 13539 8730
rect 13591 8678 13603 8730
rect 13655 8678 13667 8730
rect 13719 8678 16008 8730
rect 1104 8656 16008 8678
rect 7190 8616 7196 8628
rect 2148 8588 7196 8616
rect 2148 8489 2176 8588
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8665 8619 8723 8625
rect 8665 8616 8677 8619
rect 7800 8588 8677 8616
rect 7800 8576 7806 8588
rect 8665 8585 8677 8588
rect 8711 8585 8723 8619
rect 9490 8616 9496 8628
rect 9451 8588 9496 8616
rect 8665 8579 8723 8585
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 10008 8588 10456 8616
rect 10008 8576 10014 8588
rect 4433 8551 4491 8557
rect 4433 8517 4445 8551
rect 4479 8548 4491 8551
rect 4890 8548 4896 8560
rect 4479 8520 4896 8548
rect 4479 8517 4491 8520
rect 4433 8511 4491 8517
rect 4890 8508 4896 8520
rect 4948 8508 4954 8560
rect 6178 8508 6184 8560
rect 6236 8548 6242 8560
rect 6457 8551 6515 8557
rect 6457 8548 6469 8551
rect 6236 8520 6469 8548
rect 6236 8508 6242 8520
rect 6457 8517 6469 8520
rect 6503 8548 6515 8551
rect 6914 8548 6920 8560
rect 6503 8520 6920 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 7009 8551 7067 8557
rect 7009 8517 7021 8551
rect 7055 8548 7067 8551
rect 7837 8551 7895 8557
rect 7055 8520 7788 8548
rect 7055 8517 7067 8520
rect 7009 8511 7067 8517
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 4982 8480 4988 8492
rect 2133 8443 2191 8449
rect 4448 8452 4988 8480
rect 1578 8412 1584 8424
rect 1539 8384 1584 8412
rect 1578 8372 1584 8384
rect 1636 8372 1642 8424
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 3053 8415 3111 8421
rect 3053 8412 3065 8415
rect 2096 8384 3065 8412
rect 2096 8372 2102 8384
rect 3053 8381 3065 8384
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 3068 8288 3096 8375
rect 3326 8353 3332 8356
rect 3320 8344 3332 8353
rect 3287 8316 3332 8344
rect 3320 8307 3332 8316
rect 3326 8304 3332 8307
rect 3384 8304 3390 8356
rect 3050 8276 3056 8288
rect 2963 8248 3056 8276
rect 3050 8236 3056 8248
rect 3108 8276 3114 8288
rect 4448 8276 4476 8452
rect 4982 8440 4988 8452
rect 5040 8480 5046 8492
rect 5077 8483 5135 8489
rect 5077 8480 5089 8483
rect 5040 8452 5089 8480
rect 5040 8440 5046 8452
rect 5077 8449 5089 8452
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 6638 8480 6644 8492
rect 6328 8452 6644 8480
rect 6328 8440 6334 8452
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8449 7711 8483
rect 7760 8480 7788 8520
rect 7837 8517 7849 8551
rect 7883 8548 7895 8551
rect 8478 8548 8484 8560
rect 7883 8520 8484 8548
rect 7883 8517 7895 8520
rect 7837 8511 7895 8517
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 9766 8508 9772 8560
rect 9824 8548 9830 8560
rect 10321 8551 10379 8557
rect 10321 8548 10333 8551
rect 9824 8520 10333 8548
rect 9824 8508 9830 8520
rect 10321 8517 10333 8520
rect 10367 8517 10379 8551
rect 10428 8548 10456 8588
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10560 8588 10977 8616
rect 10560 8576 10566 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 12158 8576 12164 8628
rect 12216 8576 12222 8628
rect 10781 8551 10839 8557
rect 10781 8548 10793 8551
rect 10428 8520 10793 8548
rect 10321 8511 10379 8517
rect 10781 8517 10793 8520
rect 10827 8548 10839 8551
rect 11238 8548 11244 8560
rect 10827 8520 11244 8548
rect 10827 8517 10839 8520
rect 10781 8511 10839 8517
rect 11238 8508 11244 8520
rect 11296 8508 11302 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 11440 8520 11805 8548
rect 11440 8492 11468 8520
rect 11793 8517 11805 8520
rect 11839 8548 11851 8551
rect 12176 8548 12204 8576
rect 11839 8520 12204 8548
rect 11839 8517 11851 8520
rect 11793 8511 11851 8517
rect 12342 8508 12348 8560
rect 12400 8548 12406 8560
rect 12437 8551 12495 8557
rect 12437 8548 12449 8551
rect 12400 8520 12449 8548
rect 12400 8508 12406 8520
rect 12437 8517 12449 8520
rect 12483 8517 12495 8551
rect 12437 8511 12495 8517
rect 8294 8480 8300 8492
rect 7760 8452 8300 8480
rect 7653 8443 7711 8449
rect 4522 8372 4528 8424
rect 4580 8412 4586 8424
rect 4709 8415 4767 8421
rect 4709 8412 4721 8415
rect 4580 8384 4721 8412
rect 4580 8372 4586 8384
rect 4709 8381 4721 8384
rect 4755 8381 4767 8415
rect 4709 8375 4767 8381
rect 5344 8415 5402 8421
rect 5344 8381 5356 8415
rect 5390 8412 5402 8415
rect 6362 8412 6368 8424
rect 5390 8384 6368 8412
rect 5390 8381 5402 8384
rect 5344 8375 5402 8381
rect 6362 8372 6368 8384
rect 6420 8372 6426 8424
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8412 7527 8415
rect 7668 8412 7696 8443
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8449 8447 8483
rect 8389 8443 8447 8449
rect 8110 8412 8116 8424
rect 7515 8384 7604 8412
rect 7668 8384 8116 8412
rect 7515 8381 7527 8384
rect 7469 8375 7527 8381
rect 7576 8288 7604 8384
rect 8110 8372 8116 8384
rect 8168 8412 8174 8424
rect 8404 8412 8432 8443
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 9180 8452 9229 8480
rect 9180 8440 9186 8452
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 10134 8480 10140 8492
rect 10095 8452 10140 8480
rect 9217 8443 9275 8449
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 11422 8480 11428 8492
rect 11383 8452 11428 8480
rect 11422 8440 11428 8452
rect 11480 8440 11486 8492
rect 11609 8483 11667 8489
rect 11609 8449 11621 8483
rect 11655 8480 11667 8483
rect 12710 8480 12716 8492
rect 11655 8452 12716 8480
rect 11655 8449 11667 8452
rect 11609 8443 11667 8449
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12986 8480 12992 8492
rect 12947 8452 12992 8480
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 8168 8384 8432 8412
rect 8168 8372 8174 8384
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 9953 8415 10011 8421
rect 9953 8412 9965 8415
rect 8720 8384 9965 8412
rect 8720 8372 8726 8384
rect 9953 8381 9965 8384
rect 9999 8412 10011 8415
rect 10318 8412 10324 8424
rect 9999 8384 10324 8412
rect 9999 8381 10011 8384
rect 9953 8375 10011 8381
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 10502 8412 10508 8424
rect 10463 8384 10508 8412
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8412 10747 8415
rect 11790 8412 11796 8424
rect 10735 8384 11796 8412
rect 10735 8381 10747 8384
rect 10689 8375 10747 8381
rect 9125 8347 9183 8353
rect 9125 8313 9137 8347
rect 9171 8344 9183 8347
rect 9306 8344 9312 8356
rect 9171 8316 9312 8344
rect 9171 8313 9183 8316
rect 9125 8307 9183 8313
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 9861 8347 9919 8353
rect 9861 8313 9873 8347
rect 9907 8344 9919 8347
rect 10594 8344 10600 8356
rect 9907 8316 10600 8344
rect 9907 8313 9919 8316
rect 9861 8307 9919 8313
rect 10594 8304 10600 8316
rect 10652 8344 10658 8356
rect 10704 8344 10732 8375
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 12066 8412 12072 8424
rect 11979 8384 12072 8412
rect 12066 8372 12072 8384
rect 12124 8412 12130 8424
rect 12802 8412 12808 8424
rect 12124 8384 12388 8412
rect 12763 8384 12808 8412
rect 12124 8372 12130 8384
rect 10652 8316 10732 8344
rect 11333 8347 11391 8353
rect 10652 8304 10658 8316
rect 11333 8313 11345 8347
rect 11379 8344 11391 8347
rect 12161 8347 12219 8353
rect 12161 8344 12173 8347
rect 11379 8316 12173 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 12161 8313 12173 8316
rect 12207 8344 12219 8347
rect 12360 8344 12388 8384
rect 12802 8372 12808 8384
rect 12860 8372 12866 8424
rect 13906 8412 13912 8424
rect 12912 8384 13912 8412
rect 12912 8344 12940 8384
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 13170 8344 13176 8356
rect 12207 8316 12296 8344
rect 12360 8316 12940 8344
rect 13083 8316 13176 8344
rect 12207 8313 12219 8316
rect 12161 8307 12219 8313
rect 4525 8279 4583 8285
rect 4525 8276 4537 8279
rect 3108 8248 4537 8276
rect 3108 8236 3114 8248
rect 4525 8245 4537 8248
rect 4571 8245 4583 8279
rect 6638 8276 6644 8288
rect 6599 8248 6644 8276
rect 4525 8239 4583 8245
rect 6638 8236 6644 8248
rect 6696 8236 6702 8288
rect 6917 8279 6975 8285
rect 6917 8245 6929 8279
rect 6963 8276 6975 8279
rect 7377 8279 7435 8285
rect 7377 8276 7389 8279
rect 6963 8248 7389 8276
rect 6963 8245 6975 8248
rect 6917 8239 6975 8245
rect 7377 8245 7389 8248
rect 7423 8276 7435 8279
rect 7466 8276 7472 8288
rect 7423 8248 7472 8276
rect 7423 8245 7435 8248
rect 7377 8239 7435 8245
rect 7466 8236 7472 8248
rect 7524 8236 7530 8288
rect 7558 8236 7564 8288
rect 7616 8236 7622 8288
rect 7742 8236 7748 8288
rect 7800 8276 7806 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7800 8248 8217 8276
rect 7800 8236 7806 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 8205 8239 8263 8245
rect 8297 8279 8355 8285
rect 8297 8245 8309 8279
rect 8343 8276 8355 8279
rect 8386 8276 8392 8288
rect 8343 8248 8392 8276
rect 8343 8245 8355 8248
rect 8297 8239 8355 8245
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 9033 8279 9091 8285
rect 9033 8245 9045 8279
rect 9079 8276 9091 8279
rect 9950 8276 9956 8288
rect 9079 8248 9956 8276
rect 9079 8245 9091 8248
rect 9033 8239 9091 8245
rect 9950 8236 9956 8248
rect 10008 8236 10014 8288
rect 10318 8236 10324 8288
rect 10376 8276 10382 8288
rect 10410 8276 10416 8288
rect 10376 8248 10416 8276
rect 10376 8236 10382 8248
rect 10410 8236 10416 8248
rect 10468 8236 10474 8288
rect 12268 8276 12296 8316
rect 12434 8276 12440 8288
rect 12268 8248 12440 8276
rect 12434 8236 12440 8248
rect 12492 8276 12498 8288
rect 12802 8276 12808 8288
rect 12492 8248 12808 8276
rect 12492 8236 12498 8248
rect 12802 8236 12808 8248
rect 12860 8236 12866 8288
rect 12897 8279 12955 8285
rect 12897 8245 12909 8279
rect 12943 8276 12955 8279
rect 13096 8276 13124 8316
rect 13170 8304 13176 8316
rect 13228 8344 13234 8356
rect 13354 8344 13360 8356
rect 13228 8316 13360 8344
rect 13228 8304 13234 8316
rect 13354 8304 13360 8316
rect 13412 8304 13418 8356
rect 12943 8248 13124 8276
rect 12943 8245 12955 8248
rect 12897 8239 12955 8245
rect 1104 8186 16008 8208
rect 1104 8134 5979 8186
rect 6031 8134 6043 8186
rect 6095 8134 6107 8186
rect 6159 8134 6171 8186
rect 6223 8134 10976 8186
rect 11028 8134 11040 8186
rect 11092 8134 11104 8186
rect 11156 8134 11168 8186
rect 11220 8134 16008 8186
rect 1104 8112 16008 8134
rect 1489 8075 1547 8081
rect 1489 8041 1501 8075
rect 1535 8072 1547 8075
rect 1578 8072 1584 8084
rect 1535 8044 1584 8072
rect 1535 8041 1547 8044
rect 1489 8035 1547 8041
rect 1578 8032 1584 8044
rect 1636 8072 1642 8084
rect 5534 8072 5540 8084
rect 1636 8044 5304 8072
rect 5495 8044 5540 8072
rect 1636 8032 1642 8044
rect 5276 8004 5304 8044
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 7926 8072 7932 8084
rect 5776 8044 7932 8072
rect 5776 8032 5782 8044
rect 7926 8032 7932 8044
rect 7984 8072 7990 8084
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 7984 8044 8033 8072
rect 7984 8032 7990 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 8021 8035 8079 8041
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8041 8171 8075
rect 8478 8072 8484 8084
rect 8439 8044 8484 8072
rect 8113 8035 8171 8041
rect 5276 7976 6500 8004
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 2038 7936 2044 7948
rect 1995 7908 2044 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 2038 7896 2044 7908
rect 2096 7896 2102 7948
rect 2216 7939 2274 7945
rect 2216 7905 2228 7939
rect 2262 7936 2274 7939
rect 3234 7936 3240 7948
rect 2262 7908 3240 7936
rect 2262 7905 2274 7908
rect 2216 7899 2274 7905
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 4706 7936 4712 7948
rect 4479 7908 4712 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 5902 7936 5908 7948
rect 4856 7908 5488 7936
rect 5863 7908 5908 7936
rect 4856 7896 4862 7908
rect 5460 7880 5488 7908
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 3878 7828 3884 7880
rect 3936 7868 3942 7880
rect 4525 7871 4583 7877
rect 4525 7868 4537 7871
rect 3936 7840 4537 7868
rect 3936 7828 3942 7840
rect 4525 7837 4537 7840
rect 4571 7837 4583 7871
rect 4525 7831 4583 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4893 7871 4951 7877
rect 4893 7837 4905 7871
rect 4939 7868 4951 7871
rect 5074 7868 5080 7880
rect 4939 7840 5080 7868
rect 4939 7837 4951 7840
rect 4893 7831 4951 7837
rect 3326 7800 3332 7812
rect 3239 7772 3332 7800
rect 3326 7760 3332 7772
rect 3384 7800 3390 7812
rect 4632 7800 4660 7831
rect 5074 7828 5080 7840
rect 5132 7828 5138 7880
rect 5442 7868 5448 7880
rect 5355 7840 5448 7868
rect 5442 7828 5448 7840
rect 5500 7868 5506 7880
rect 5997 7871 6055 7877
rect 5997 7868 6009 7871
rect 5500 7840 6009 7868
rect 5500 7828 5506 7840
rect 5997 7837 6009 7840
rect 6043 7868 6055 7871
rect 6086 7868 6092 7880
rect 6043 7840 6092 7868
rect 6043 7837 6055 7840
rect 5997 7831 6055 7837
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7868 6239 7871
rect 6362 7868 6368 7880
rect 6227 7840 6368 7868
rect 6227 7837 6239 7840
rect 6181 7831 6239 7837
rect 6362 7828 6368 7840
rect 6420 7828 6426 7880
rect 3384 7772 4660 7800
rect 3384 7760 3390 7772
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 2924 7704 4077 7732
rect 2924 7692 2930 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4065 7695 4123 7701
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 5169 7735 5227 7741
rect 5169 7732 5181 7735
rect 4672 7704 5181 7732
rect 4672 7692 4678 7704
rect 5169 7701 5181 7704
rect 5215 7701 5227 7735
rect 6362 7732 6368 7744
rect 6323 7704 6368 7732
rect 5169 7695 5227 7701
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 6472 7732 6500 7976
rect 6730 7964 6736 8016
rect 6788 8004 6794 8016
rect 8128 8004 8156 8035
rect 8478 8032 8484 8044
rect 8536 8032 8542 8084
rect 8938 8072 8944 8084
rect 8899 8044 8944 8072
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 9306 8032 9312 8084
rect 9364 8072 9370 8084
rect 9582 8072 9588 8084
rect 9364 8044 9588 8072
rect 9364 8032 9370 8044
rect 9582 8032 9588 8044
rect 9640 8072 9646 8084
rect 9677 8075 9735 8081
rect 9677 8072 9689 8075
rect 9640 8044 9689 8072
rect 9640 8032 9646 8044
rect 9677 8041 9689 8044
rect 9723 8041 9735 8075
rect 9950 8072 9956 8084
rect 9863 8044 9956 8072
rect 9677 8035 9735 8041
rect 9950 8032 9956 8044
rect 10008 8072 10014 8084
rect 10778 8072 10784 8084
rect 10008 8044 10784 8072
rect 10008 8032 10014 8044
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 11330 8032 11336 8084
rect 11388 8032 11394 8084
rect 11422 8032 11428 8084
rect 11480 8072 11486 8084
rect 12158 8072 12164 8084
rect 11480 8044 12164 8072
rect 11480 8032 11486 8044
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 12710 8032 12716 8084
rect 12768 8072 12774 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 12768 8044 14105 8072
rect 12768 8032 12774 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 6788 7976 8156 8004
rect 6788 7964 6794 7976
rect 8294 7964 8300 8016
rect 8352 8004 8358 8016
rect 8573 8007 8631 8013
rect 8573 8004 8585 8007
rect 8352 7976 8585 8004
rect 8352 7964 8358 7976
rect 8573 7973 8585 7976
rect 8619 7973 8631 8007
rect 8573 7967 8631 7973
rect 8754 7964 8760 8016
rect 8812 8004 8818 8016
rect 9122 8004 9128 8016
rect 8812 7976 9128 8004
rect 8812 7964 8818 7976
rect 9122 7964 9128 7976
rect 9180 7964 9186 8016
rect 9766 7964 9772 8016
rect 9824 8004 9830 8016
rect 11348 8004 11376 8032
rect 9824 7976 12756 8004
rect 9824 7964 9830 7976
rect 6546 7896 6552 7948
rect 6604 7936 6610 7948
rect 6914 7945 6920 7948
rect 6908 7936 6920 7945
rect 6604 7908 6649 7936
rect 6827 7908 6920 7936
rect 6604 7896 6610 7908
rect 6908 7899 6920 7908
rect 6972 7936 6978 7948
rect 6972 7908 8800 7936
rect 6914 7896 6920 7899
rect 6972 7896 6978 7908
rect 8772 7877 8800 7908
rect 8938 7896 8944 7948
rect 8996 7936 9002 7948
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 8996 7908 9229 7936
rect 8996 7896 9002 7908
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 10686 7936 10692 7948
rect 10647 7908 10692 7936
rect 9217 7899 9275 7905
rect 10686 7896 10692 7908
rect 10744 7896 10750 7948
rect 11256 7945 11284 7976
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7905 11299 7939
rect 11241 7899 11299 7905
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 12728 7945 12756 7976
rect 11497 7939 11555 7945
rect 11497 7936 11509 7939
rect 11388 7908 11509 7936
rect 11388 7896 11394 7908
rect 11497 7905 11509 7908
rect 11543 7905 11555 7939
rect 11497 7899 11555 7905
rect 12713 7939 12771 7945
rect 12713 7905 12725 7939
rect 12759 7905 12771 7939
rect 12969 7939 13027 7945
rect 12969 7936 12981 7939
rect 12713 7899 12771 7905
rect 12820 7908 12981 7936
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7837 8815 7871
rect 8757 7831 8815 7837
rect 6546 7760 6552 7812
rect 6604 7800 6610 7812
rect 6656 7800 6684 7831
rect 9398 7828 9404 7880
rect 9456 7868 9462 7880
rect 10594 7868 10600 7880
rect 9456 7840 10600 7868
rect 9456 7828 9462 7840
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 10778 7868 10784 7880
rect 10739 7840 10784 7868
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7837 11023 7871
rect 12820 7868 12848 7908
rect 12969 7905 12981 7908
rect 13015 7905 13027 7939
rect 12969 7899 13027 7905
rect 10965 7831 11023 7837
rect 12636 7840 12848 7868
rect 10134 7800 10140 7812
rect 6604 7772 6684 7800
rect 7576 7772 10140 7800
rect 6604 7760 6610 7772
rect 7576 7732 7604 7772
rect 10134 7760 10140 7772
rect 10192 7760 10198 7812
rect 6472 7704 7604 7732
rect 7650 7692 7656 7744
rect 7708 7732 7714 7744
rect 9401 7735 9459 7741
rect 9401 7732 9413 7735
rect 7708 7704 9413 7732
rect 7708 7692 7714 7704
rect 9401 7701 9413 7704
rect 9447 7701 9459 7735
rect 10318 7732 10324 7744
rect 10279 7704 10324 7732
rect 9401 7695 9459 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 10980 7732 11008 7831
rect 12636 7741 12664 7840
rect 12621 7735 12679 7741
rect 12621 7732 12633 7735
rect 10980 7704 12633 7732
rect 12621 7701 12633 7704
rect 12667 7701 12679 7735
rect 12621 7695 12679 7701
rect 1104 7642 16008 7664
rect 1104 7590 3480 7642
rect 3532 7590 3544 7642
rect 3596 7590 3608 7642
rect 3660 7590 3672 7642
rect 3724 7590 8478 7642
rect 8530 7590 8542 7642
rect 8594 7590 8606 7642
rect 8658 7590 8670 7642
rect 8722 7590 13475 7642
rect 13527 7590 13539 7642
rect 13591 7590 13603 7642
rect 13655 7590 13667 7642
rect 13719 7590 16008 7642
rect 1104 7568 16008 7590
rect 3878 7528 3884 7540
rect 3839 7500 3884 7528
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 4706 7528 4712 7540
rect 4667 7500 4712 7528
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 5810 7528 5816 7540
rect 5771 7500 5816 7528
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 10318 7528 10324 7540
rect 6604 7500 10324 7528
rect 6604 7488 6610 7500
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 10686 7488 10692 7540
rect 10744 7528 10750 7540
rect 11425 7531 11483 7537
rect 11425 7528 11437 7531
rect 10744 7500 11437 7528
rect 10744 7488 10750 7500
rect 11425 7497 11437 7500
rect 11471 7497 11483 7531
rect 11425 7491 11483 7497
rect 10134 7420 10140 7472
rect 10192 7460 10198 7472
rect 14826 7460 14832 7472
rect 10192 7432 14832 7460
rect 10192 7420 10198 7432
rect 14826 7420 14832 7432
rect 14884 7420 14890 7472
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 3326 7392 3332 7404
rect 3287 7364 3332 7392
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 3712 7364 4445 7392
rect 1489 7327 1547 7333
rect 1489 7293 1501 7327
rect 1535 7324 1547 7327
rect 3142 7324 3148 7336
rect 1535 7296 3148 7324
rect 1535 7293 1547 7296
rect 1489 7287 1547 7293
rect 3142 7284 3148 7296
rect 3200 7284 3206 7336
rect 3234 7284 3240 7336
rect 3292 7324 3298 7336
rect 3712 7324 3740 7364
rect 4433 7361 4445 7364
rect 4479 7392 4491 7395
rect 5261 7395 5319 7401
rect 5261 7392 5273 7395
rect 4479 7364 5273 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 5261 7361 5273 7364
rect 5307 7361 5319 7395
rect 5810 7392 5816 7404
rect 5261 7355 5319 7361
rect 5552 7364 5816 7392
rect 3292 7296 3740 7324
rect 3292 7284 3298 7296
rect 3786 7284 3792 7336
rect 3844 7324 3850 7336
rect 5074 7324 5080 7336
rect 3844 7296 4752 7324
rect 5035 7296 5080 7324
rect 3844 7284 3850 7296
rect 3053 7259 3111 7265
rect 3053 7225 3065 7259
rect 3099 7256 3111 7259
rect 4062 7256 4068 7268
rect 3099 7228 4068 7256
rect 3099 7225 3111 7228
rect 3053 7219 3111 7225
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 4341 7259 4399 7265
rect 4341 7225 4353 7259
rect 4387 7256 4399 7259
rect 4614 7256 4620 7268
rect 4387 7228 4620 7256
rect 4387 7225 4399 7228
rect 4341 7219 4399 7225
rect 4614 7216 4620 7228
rect 4672 7216 4678 7268
rect 4724 7256 4752 7296
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 5166 7284 5172 7336
rect 5224 7324 5230 7336
rect 5552 7324 5580 7364
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 6914 7392 6920 7404
rect 6512 7364 6920 7392
rect 6512 7352 6518 7364
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7006 7352 7012 7404
rect 7064 7392 7070 7404
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 7064 7364 7389 7392
rect 7064 7352 7070 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 7377 7355 7435 7361
rect 10520 7364 11161 7392
rect 5224 7296 5580 7324
rect 5224 7284 5230 7296
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 5684 7296 5729 7324
rect 5684 7284 5690 7296
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 5960 7296 6684 7324
rect 5960 7284 5966 7296
rect 6656 7268 6684 7296
rect 7098 7284 7104 7336
rect 7156 7324 7162 7336
rect 7193 7327 7251 7333
rect 7193 7324 7205 7327
rect 7156 7296 7205 7324
rect 7156 7284 7162 7296
rect 7193 7293 7205 7296
rect 7239 7293 7251 7327
rect 7193 7287 7251 7293
rect 7282 7284 7288 7336
rect 7340 7324 7346 7336
rect 7653 7327 7711 7333
rect 7340 7296 7604 7324
rect 7340 7284 7346 7296
rect 6181 7259 6239 7265
rect 6181 7256 6193 7259
rect 4724 7228 6193 7256
rect 6181 7225 6193 7228
rect 6227 7256 6239 7259
rect 6546 7256 6552 7268
rect 6227 7228 6552 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 6546 7216 6552 7228
rect 6604 7216 6610 7268
rect 6638 7216 6644 7268
rect 6696 7256 6702 7268
rect 7374 7256 7380 7268
rect 6696 7228 7380 7256
rect 6696 7216 6702 7228
rect 7374 7216 7380 7228
rect 7432 7216 7438 7268
rect 2682 7188 2688 7200
rect 2643 7160 2688 7188
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 3142 7148 3148 7200
rect 3200 7188 3206 7200
rect 4246 7188 4252 7200
rect 3200 7160 3245 7188
rect 4159 7160 4252 7188
rect 3200 7148 3206 7160
rect 4246 7148 4252 7160
rect 4304 7188 4310 7200
rect 5626 7188 5632 7200
rect 4304 7160 5632 7188
rect 4304 7148 4310 7160
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6273 7191 6331 7197
rect 6273 7157 6285 7191
rect 6319 7188 6331 7191
rect 6825 7191 6883 7197
rect 6825 7188 6837 7191
rect 6319 7160 6837 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 6825 7157 6837 7160
rect 6871 7157 6883 7191
rect 7576 7188 7604 7296
rect 7653 7293 7665 7327
rect 7699 7324 7711 7327
rect 7742 7324 7748 7336
rect 7699 7296 7748 7324
rect 7699 7293 7711 7296
rect 7653 7287 7711 7293
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 7926 7333 7932 7336
rect 7920 7287 7932 7333
rect 7984 7324 7990 7336
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 7984 7296 8020 7324
rect 8128 7296 9137 7324
rect 7926 7284 7932 7287
rect 7984 7284 7990 7296
rect 7760 7256 7788 7284
rect 8128 7256 8156 7296
rect 9125 7293 9137 7296
rect 9171 7324 9183 7327
rect 9766 7324 9772 7336
rect 9171 7296 9772 7324
rect 9171 7293 9183 7296
rect 9125 7287 9183 7293
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 9306 7256 9312 7268
rect 7760 7228 8156 7256
rect 9048 7228 9312 7256
rect 7742 7188 7748 7200
rect 7576 7160 7748 7188
rect 6825 7151 6883 7157
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 9048 7197 9076 7228
rect 9306 7216 9312 7228
rect 9364 7265 9370 7268
rect 9364 7259 9428 7265
rect 9364 7225 9382 7259
rect 9416 7225 9428 7259
rect 9364 7219 9428 7225
rect 9364 7216 9370 7219
rect 9033 7191 9091 7197
rect 9033 7157 9045 7191
rect 9079 7157 9091 7191
rect 9033 7151 9091 7157
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10520 7197 10548 7364
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 11330 7352 11336 7404
rect 11388 7392 11394 7404
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11388 7364 11989 7392
rect 11388 7352 11394 7364
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 10594 7284 10600 7336
rect 10652 7324 10658 7336
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 10652 7296 11069 7324
rect 10652 7284 10658 7296
rect 11057 7293 11069 7296
rect 11103 7324 11115 7327
rect 11422 7324 11428 7336
rect 11103 7296 11428 7324
rect 11103 7293 11115 7296
rect 11057 7287 11115 7293
rect 11422 7284 11428 7296
rect 11480 7284 11486 7336
rect 11882 7284 11888 7336
rect 11940 7324 11946 7336
rect 12066 7324 12072 7336
rect 11940 7296 12072 7324
rect 11940 7284 11946 7296
rect 12066 7284 12072 7296
rect 12124 7284 12130 7336
rect 10686 7216 10692 7268
rect 10744 7256 10750 7268
rect 10870 7256 10876 7268
rect 10744 7228 10876 7256
rect 10744 7216 10750 7228
rect 10870 7216 10876 7228
rect 10928 7256 10934 7268
rect 10965 7259 11023 7265
rect 10965 7256 10977 7259
rect 10928 7228 10977 7256
rect 10928 7216 10934 7228
rect 10965 7225 10977 7228
rect 11011 7225 11023 7259
rect 10965 7219 11023 7225
rect 11793 7259 11851 7265
rect 11793 7225 11805 7259
rect 11839 7256 11851 7259
rect 12434 7256 12440 7268
rect 11839 7228 12440 7256
rect 11839 7225 11851 7228
rect 11793 7219 11851 7225
rect 12434 7216 12440 7228
rect 12492 7216 12498 7268
rect 10505 7191 10563 7197
rect 10505 7188 10517 7191
rect 9916 7160 10517 7188
rect 9916 7148 9922 7160
rect 10505 7157 10517 7160
rect 10551 7157 10563 7191
rect 10505 7151 10563 7157
rect 10594 7148 10600 7200
rect 10652 7188 10658 7200
rect 11882 7188 11888 7200
rect 10652 7160 10697 7188
rect 11843 7160 11888 7188
rect 10652 7148 10658 7160
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 1104 7098 16008 7120
rect 1104 7046 5979 7098
rect 6031 7046 6043 7098
rect 6095 7046 6107 7098
rect 6159 7046 6171 7098
rect 6223 7046 10976 7098
rect 11028 7046 11040 7098
rect 11092 7046 11104 7098
rect 11156 7046 11168 7098
rect 11220 7046 16008 7098
rect 1104 7024 16008 7046
rect 2593 6987 2651 6993
rect 2593 6953 2605 6987
rect 2639 6984 2651 6987
rect 2682 6984 2688 6996
rect 2639 6956 2688 6984
rect 2639 6953 2651 6956
rect 2593 6947 2651 6953
rect 2682 6944 2688 6956
rect 2740 6944 2746 6996
rect 2961 6987 3019 6993
rect 2961 6953 2973 6987
rect 3007 6984 3019 6987
rect 3142 6984 3148 6996
rect 3007 6956 3148 6984
rect 3007 6953 3019 6956
rect 2961 6947 3019 6953
rect 3142 6944 3148 6956
rect 3200 6944 3206 6996
rect 3329 6987 3387 6993
rect 3329 6953 3341 6987
rect 3375 6984 3387 6987
rect 3786 6984 3792 6996
rect 3375 6956 3792 6984
rect 3375 6953 3387 6956
rect 3329 6947 3387 6953
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 4062 6984 4068 6996
rect 4023 6956 4068 6984
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 5442 6984 5448 6996
rect 5403 6956 5448 6984
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 6546 6984 6552 6996
rect 6507 6956 6552 6984
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 8110 6984 8116 6996
rect 6972 6956 8116 6984
rect 6972 6944 6978 6956
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 8294 6984 8300 6996
rect 8255 6956 8300 6984
rect 8294 6944 8300 6956
rect 8352 6984 8358 6996
rect 9217 6987 9275 6993
rect 9217 6984 9229 6987
rect 8352 6956 9229 6984
rect 8352 6944 8358 6956
rect 9217 6953 9229 6956
rect 9263 6953 9275 6987
rect 11422 6984 11428 6996
rect 11383 6956 11428 6984
rect 9217 6947 9275 6953
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 11609 6987 11667 6993
rect 11609 6953 11621 6987
rect 11655 6984 11667 6987
rect 11882 6984 11888 6996
rect 11655 6956 11888 6984
rect 11655 6953 11667 6956
rect 11609 6947 11667 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 12492 6956 12537 6984
rect 12492 6944 12498 6956
rect 2501 6919 2559 6925
rect 2501 6885 2513 6919
rect 2547 6916 2559 6919
rect 2866 6916 2872 6928
rect 2547 6888 2872 6916
rect 2547 6885 2559 6888
rect 2501 6879 2559 6885
rect 2866 6876 2872 6888
rect 2924 6876 2930 6928
rect 3234 6876 3240 6928
rect 3292 6916 3298 6928
rect 4525 6919 4583 6925
rect 3292 6888 3556 6916
rect 3292 6876 3298 6888
rect 1489 6851 1547 6857
rect 1489 6817 1501 6851
rect 1535 6817 1547 6851
rect 1489 6811 1547 6817
rect 1504 6712 1532 6811
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 3421 6851 3479 6857
rect 3421 6848 3433 6851
rect 3384 6820 3433 6848
rect 3384 6808 3390 6820
rect 3421 6817 3433 6820
rect 3467 6817 3479 6851
rect 3421 6811 3479 6817
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 2774 6780 2780 6792
rect 2735 6752 2780 6780
rect 2774 6740 2780 6752
rect 2832 6740 2838 6792
rect 3528 6789 3556 6888
rect 4525 6885 4537 6919
rect 4571 6916 4583 6919
rect 4982 6916 4988 6928
rect 4571 6888 4988 6916
rect 4571 6885 4583 6888
rect 4525 6879 4583 6885
rect 4982 6876 4988 6888
rect 5040 6916 5046 6928
rect 5460 6916 5488 6944
rect 6362 6916 6368 6928
rect 5040 6888 5488 6916
rect 5736 6888 6368 6916
rect 5040 6876 5046 6888
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6848 4491 6851
rect 5077 6851 5135 6857
rect 4479 6820 5028 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 3513 6783 3571 6789
rect 3513 6749 3525 6783
rect 3559 6780 3571 6783
rect 4062 6780 4068 6792
rect 3559 6752 4068 6780
rect 3559 6749 3571 6752
rect 3513 6743 3571 6749
rect 4062 6740 4068 6752
rect 4120 6780 4126 6792
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 4120 6752 4629 6780
rect 4120 6740 4126 6752
rect 4617 6749 4629 6752
rect 4663 6749 4675 6783
rect 5000 6780 5028 6820
rect 5077 6817 5089 6851
rect 5123 6848 5135 6851
rect 5736 6848 5764 6888
rect 6362 6876 6368 6888
rect 6420 6916 6426 6928
rect 6420 6888 7144 6916
rect 6420 6876 6426 6888
rect 5902 6848 5908 6860
rect 5123 6820 5764 6848
rect 5863 6820 5908 6848
rect 5123 6817 5135 6820
rect 5077 6811 5135 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 5997 6851 6055 6857
rect 5997 6817 6009 6851
rect 6043 6848 6055 6851
rect 6822 6848 6828 6860
rect 6043 6820 6828 6848
rect 6043 6817 6055 6820
rect 5997 6811 6055 6817
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 7006 6857 7012 6860
rect 7000 6848 7012 6857
rect 6967 6820 7012 6848
rect 7000 6811 7012 6820
rect 7006 6808 7012 6811
rect 7064 6808 7070 6860
rect 7116 6848 7144 6888
rect 7374 6876 7380 6928
rect 7432 6916 7438 6928
rect 10134 6916 10140 6928
rect 7432 6888 10140 6916
rect 7432 6876 7438 6888
rect 10134 6876 10140 6888
rect 10192 6876 10198 6928
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 11241 6919 11299 6925
rect 11241 6916 11253 6919
rect 10744 6888 11253 6916
rect 10744 6876 10750 6888
rect 11241 6885 11253 6888
rect 11287 6885 11299 6919
rect 11241 6879 11299 6885
rect 11790 6876 11796 6928
rect 11848 6916 11854 6928
rect 11977 6919 12035 6925
rect 11977 6916 11989 6919
rect 11848 6888 11989 6916
rect 11848 6876 11854 6888
rect 11977 6885 11989 6888
rect 12023 6916 12035 6919
rect 13170 6916 13176 6928
rect 12023 6888 13176 6916
rect 12023 6885 12035 6888
rect 11977 6879 12035 6885
rect 13170 6876 13176 6888
rect 13228 6876 13234 6928
rect 8665 6851 8723 6857
rect 8665 6848 8677 6851
rect 7116 6820 8677 6848
rect 8665 6817 8677 6820
rect 8711 6817 8723 6851
rect 9122 6848 9128 6860
rect 9083 6820 9128 6848
rect 8665 6811 8723 6817
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 9766 6848 9772 6860
rect 9727 6820 9772 6848
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 10025 6851 10083 6857
rect 10025 6848 10037 6851
rect 9916 6820 10037 6848
rect 9916 6808 9922 6820
rect 10025 6817 10037 6820
rect 10071 6848 10083 6851
rect 12066 6848 12072 6860
rect 10071 6820 11008 6848
rect 12027 6820 12072 6848
rect 10071 6817 10083 6820
rect 10025 6811 10083 6817
rect 6089 6783 6147 6789
rect 5000 6752 5304 6780
rect 4617 6743 4675 6749
rect 4338 6712 4344 6724
rect 1504 6684 4344 6712
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 5276 6656 5304 6752
rect 6089 6749 6101 6783
rect 6135 6749 6147 6783
rect 6089 6743 6147 6749
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6749 6791 6783
rect 6733 6743 6791 6749
rect 5718 6672 5724 6724
rect 5776 6712 5782 6724
rect 6104 6712 6132 6743
rect 5776 6684 6132 6712
rect 5776 6672 5782 6684
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 2133 6647 2191 6653
rect 2133 6644 2145 6647
rect 1544 6616 2145 6644
rect 1544 6604 1550 6616
rect 2133 6613 2145 6616
rect 2179 6613 2191 6647
rect 2133 6607 2191 6613
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 4893 6647 4951 6653
rect 4893 6644 4905 6647
rect 4580 6616 4905 6644
rect 4580 6604 4586 6616
rect 4893 6613 4905 6616
rect 4939 6613 4951 6647
rect 5258 6644 5264 6656
rect 5219 6616 5264 6644
rect 4893 6607 4951 6613
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 5537 6647 5595 6653
rect 5537 6613 5549 6647
rect 5583 6644 5595 6647
rect 5626 6644 5632 6656
rect 5583 6616 5632 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 6362 6644 6368 6656
rect 5868 6616 6368 6644
rect 5868 6604 5874 6616
rect 6362 6604 6368 6616
rect 6420 6604 6426 6656
rect 6748 6644 6776 6743
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9364 6752 9409 6780
rect 9364 6740 9370 6752
rect 8481 6715 8539 6721
rect 8481 6681 8493 6715
rect 8527 6712 8539 6715
rect 10980 6712 11008 6820
rect 12066 6808 12072 6820
rect 12124 6808 12130 6860
rect 12802 6848 12808 6860
rect 12763 6820 12808 6848
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 13354 6848 13360 6860
rect 12912 6820 13360 6848
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6749 12219 6783
rect 12161 6743 12219 6749
rect 12176 6712 12204 6743
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 12912 6789 12940 6820
rect 13354 6808 13360 6820
rect 13412 6848 13418 6860
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 13412 6820 13645 6848
rect 13412 6808 13418 6820
rect 13633 6817 13645 6820
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12584 6752 12909 6780
rect 12584 6740 12590 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6749 13047 6783
rect 12989 6743 13047 6749
rect 13004 6712 13032 6743
rect 13449 6715 13507 6721
rect 13449 6712 13461 6715
rect 8527 6684 9812 6712
rect 10980 6684 13032 6712
rect 13096 6684 13461 6712
rect 8527 6681 8539 6684
rect 8481 6675 8539 6681
rect 7650 6644 7656 6656
rect 6748 6616 7656 6644
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6644 8815 6647
rect 9674 6644 9680 6656
rect 8803 6616 9680 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 9784 6644 9812 6684
rect 9950 6644 9956 6656
rect 9784 6616 9956 6644
rect 9950 6604 9956 6616
rect 10008 6644 10014 6656
rect 10502 6644 10508 6656
rect 10008 6616 10508 6644
rect 10008 6604 10014 6616
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 11146 6644 11152 6656
rect 11107 6616 11152 6644
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 12066 6604 12072 6656
rect 12124 6644 12130 6656
rect 13096 6644 13124 6684
rect 13449 6681 13461 6684
rect 13495 6681 13507 6715
rect 13449 6675 13507 6681
rect 12124 6616 13124 6644
rect 12124 6604 12130 6616
rect 13170 6604 13176 6656
rect 13228 6644 13234 6656
rect 13265 6647 13323 6653
rect 13265 6644 13277 6647
rect 13228 6616 13277 6644
rect 13228 6604 13234 6616
rect 13265 6613 13277 6616
rect 13311 6613 13323 6647
rect 13265 6607 13323 6613
rect 1104 6554 16008 6576
rect 1104 6502 3480 6554
rect 3532 6502 3544 6554
rect 3596 6502 3608 6554
rect 3660 6502 3672 6554
rect 3724 6502 8478 6554
rect 8530 6502 8542 6554
rect 8594 6502 8606 6554
rect 8658 6502 8670 6554
rect 8722 6502 13475 6554
rect 13527 6502 13539 6554
rect 13591 6502 13603 6554
rect 13655 6502 13667 6554
rect 13719 6502 16008 6554
rect 1104 6480 16008 6502
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 4525 6443 4583 6449
rect 4525 6440 4537 6443
rect 4120 6412 4537 6440
rect 4120 6400 4126 6412
rect 4525 6409 4537 6412
rect 4571 6409 4583 6443
rect 4525 6403 4583 6409
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 5960 6412 6837 6440
rect 5960 6400 5966 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 7098 6400 7104 6452
rect 7156 6440 7162 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 7156 6412 7849 6440
rect 7156 6400 7162 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 7837 6403 7895 6409
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8113 6443 8171 6449
rect 8113 6440 8125 6443
rect 8076 6412 8125 6440
rect 8076 6400 8082 6412
rect 8113 6409 8125 6412
rect 8159 6440 8171 6443
rect 8202 6440 8208 6452
rect 8159 6412 8208 6440
rect 8159 6409 8171 6412
rect 8113 6403 8171 6409
rect 8202 6400 8208 6412
rect 8260 6440 8266 6452
rect 10229 6443 10287 6449
rect 8260 6412 8892 6440
rect 8260 6400 8266 6412
rect 5997 6375 6055 6381
rect 5997 6341 6009 6375
rect 6043 6372 6055 6375
rect 6454 6372 6460 6384
rect 6043 6344 6460 6372
rect 6043 6341 6055 6344
rect 5997 6335 6055 6341
rect 6454 6332 6460 6344
rect 6512 6332 6518 6384
rect 8294 6332 8300 6384
rect 8352 6372 8358 6384
rect 8754 6372 8760 6384
rect 8352 6344 8760 6372
rect 8352 6332 8358 6344
rect 8754 6332 8760 6344
rect 8812 6332 8818 6384
rect 3050 6264 3056 6316
rect 3108 6304 3114 6316
rect 3145 6307 3203 6313
rect 3145 6304 3157 6307
rect 3108 6276 3157 6304
rect 3108 6264 3114 6276
rect 3145 6273 3157 6276
rect 3191 6273 3203 6307
rect 3145 6267 3203 6273
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6304 6239 6307
rect 6270 6304 6276 6316
rect 6227 6276 6276 6304
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 7466 6304 7472 6316
rect 7427 6276 7472 6304
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 8864 6313 8892 6412
rect 10229 6409 10241 6443
rect 10275 6440 10287 6443
rect 10778 6440 10784 6452
rect 10275 6412 10784 6440
rect 10275 6409 10287 6412
rect 10229 6403 10287 6409
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6304 9091 6307
rect 9306 6304 9312 6316
rect 9079 6276 9312 6304
rect 9079 6273 9091 6276
rect 9033 6267 9091 6273
rect 9306 6264 9312 6276
rect 9364 6264 9370 6316
rect 9674 6304 9680 6316
rect 9635 6276 9680 6304
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 9858 6304 9864 6316
rect 9819 6276 9864 6304
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6304 10931 6307
rect 11146 6304 11152 6316
rect 10919 6276 11152 6304
rect 10919 6273 10931 6276
rect 10873 6267 10931 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6304 12127 6307
rect 12802 6304 12808 6316
rect 12115 6276 12808 6304
rect 12115 6273 12127 6276
rect 12069 6267 12127 6273
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 1486 6236 1492 6248
rect 1447 6208 1492 6236
rect 1486 6196 1492 6208
rect 1544 6196 1550 6248
rect 4890 6245 4896 6248
rect 4617 6239 4675 6245
rect 4617 6205 4629 6239
rect 4663 6205 4675 6239
rect 4884 6236 4896 6245
rect 4851 6208 4896 6236
rect 4617 6199 4675 6205
rect 4884 6199 4896 6208
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 2958 6168 2964 6180
rect 1811 6140 2964 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 3418 6177 3424 6180
rect 3412 6168 3424 6177
rect 3379 6140 3424 6168
rect 3412 6131 3424 6140
rect 3418 6128 3424 6131
rect 3476 6128 3482 6180
rect 4632 6168 4660 6199
rect 4890 6196 4896 6199
rect 4948 6196 4954 6248
rect 7098 6236 7104 6248
rect 6840 6208 7104 6236
rect 5442 6168 5448 6180
rect 4632 6140 5448 6168
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 6549 6171 6607 6177
rect 6549 6137 6561 6171
rect 6595 6168 6607 6171
rect 6638 6168 6644 6180
rect 6595 6140 6644 6168
rect 6595 6137 6607 6140
rect 6549 6131 6607 6137
rect 6638 6128 6644 6140
rect 6696 6128 6702 6180
rect 5166 6060 5172 6112
rect 5224 6100 5230 6112
rect 6840 6100 6868 6208
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 8757 6239 8815 6245
rect 8757 6205 8769 6239
rect 8803 6236 8815 6239
rect 8938 6236 8944 6248
rect 8803 6208 8944 6236
rect 8803 6205 8815 6208
rect 8757 6199 8815 6205
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 9214 6236 9220 6248
rect 9048 6208 9220 6236
rect 8205 6171 8263 6177
rect 8205 6137 8217 6171
rect 8251 6168 8263 6171
rect 9048 6168 9076 6208
rect 9214 6196 9220 6208
rect 9272 6236 9278 6248
rect 9585 6239 9643 6245
rect 9585 6236 9597 6239
rect 9272 6208 9597 6236
rect 9272 6196 9278 6208
rect 9585 6205 9597 6208
rect 9631 6205 9643 6239
rect 10594 6236 10600 6248
rect 10555 6208 10600 6236
rect 9585 6199 9643 6205
rect 10594 6196 10600 6208
rect 10652 6196 10658 6248
rect 10689 6171 10747 6177
rect 10689 6168 10701 6171
rect 8251 6140 9076 6168
rect 9232 6140 10701 6168
rect 8251 6137 8263 6140
rect 8205 6131 8263 6137
rect 7190 6100 7196 6112
rect 5224 6072 6868 6100
rect 7151 6072 7196 6100
rect 5224 6060 5230 6072
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 7742 6100 7748 6112
rect 7340 6072 7385 6100
rect 7703 6072 7748 6100
rect 7340 6060 7346 6072
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 9232 6109 9260 6140
rect 10689 6137 10701 6140
rect 10735 6137 10747 6171
rect 10689 6131 10747 6137
rect 8389 6103 8447 6109
rect 8389 6100 8401 6103
rect 8352 6072 8401 6100
rect 8352 6060 8358 6072
rect 8389 6069 8401 6072
rect 8435 6069 8447 6103
rect 8389 6063 8447 6069
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6069 9275 6103
rect 9217 6063 9275 6069
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 9548 6072 10057 6100
rect 9548 6060 9554 6072
rect 10045 6069 10057 6072
rect 10091 6069 10103 6103
rect 10045 6063 10103 6069
rect 1104 6010 16008 6032
rect 1104 5958 5979 6010
rect 6031 5958 6043 6010
rect 6095 5958 6107 6010
rect 6159 5958 6171 6010
rect 6223 5958 10976 6010
rect 11028 5958 11040 6010
rect 11092 5958 11104 6010
rect 11156 5958 11168 6010
rect 11220 5958 16008 6010
rect 1104 5936 16008 5958
rect 3326 5856 3332 5908
rect 3384 5896 3390 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3384 5868 4077 5896
rect 3384 5856 3390 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4525 5899 4583 5905
rect 4525 5865 4537 5899
rect 4571 5896 4583 5899
rect 4706 5896 4712 5908
rect 4571 5868 4712 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 6880 5868 7021 5896
rect 6880 5856 6886 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 7009 5859 7067 5865
rect 7469 5899 7527 5905
rect 7469 5865 7481 5899
rect 7515 5896 7527 5899
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7515 5868 7849 5896
rect 7515 5865 7527 5868
rect 7469 5859 7527 5865
rect 7837 5865 7849 5868
rect 7883 5865 7895 5899
rect 7837 5859 7895 5865
rect 8297 5899 8355 5905
rect 8297 5865 8309 5899
rect 8343 5896 8355 5899
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 8343 5868 8677 5896
rect 8343 5865 8355 5868
rect 8297 5859 8355 5865
rect 8665 5865 8677 5868
rect 8711 5865 8723 5899
rect 8665 5859 8723 5865
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 8812 5868 9137 5896
rect 8812 5856 8818 5868
rect 9125 5865 9137 5868
rect 9171 5896 9183 5899
rect 9677 5899 9735 5905
rect 9677 5896 9689 5899
rect 9171 5868 9689 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 9677 5865 9689 5868
rect 9723 5865 9735 5899
rect 9677 5859 9735 5865
rect 10042 5856 10048 5908
rect 10100 5896 10106 5908
rect 10229 5899 10287 5905
rect 10229 5896 10241 5899
rect 10100 5868 10241 5896
rect 10100 5856 10106 5868
rect 10229 5865 10241 5868
rect 10275 5865 10287 5899
rect 10229 5859 10287 5865
rect 3050 5788 3056 5840
rect 3108 5828 3114 5840
rect 5718 5837 5724 5840
rect 3605 5831 3663 5837
rect 3605 5828 3617 5831
rect 3108 5800 3617 5828
rect 3108 5788 3114 5800
rect 3605 5797 3617 5800
rect 3651 5828 3663 5831
rect 5712 5828 5724 5837
rect 3651 5800 5580 5828
rect 5679 5800 5724 5828
rect 3651 5797 3663 5800
rect 3605 5791 3663 5797
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5760 2099 5763
rect 2130 5760 2136 5772
rect 2087 5732 2136 5760
rect 2087 5729 2099 5732
rect 2041 5723 2099 5729
rect 2130 5720 2136 5732
rect 2188 5720 2194 5772
rect 2308 5763 2366 5769
rect 2308 5729 2320 5763
rect 2354 5760 2366 5763
rect 2774 5760 2780 5772
rect 2354 5732 2780 5760
rect 2354 5729 2366 5732
rect 2308 5723 2366 5729
rect 2774 5720 2780 5732
rect 2832 5720 2838 5772
rect 3234 5720 3240 5772
rect 3292 5760 3298 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 3292 5732 4445 5760
rect 3292 5720 3298 5732
rect 4433 5729 4445 5732
rect 4479 5760 4491 5763
rect 5166 5760 5172 5772
rect 4479 5732 5172 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 5552 5760 5580 5800
rect 5712 5791 5724 5800
rect 5718 5788 5724 5791
rect 5776 5788 5782 5840
rect 7926 5828 7932 5840
rect 5828 5800 7932 5828
rect 5828 5760 5856 5800
rect 7926 5788 7932 5800
rect 7984 5828 7990 5840
rect 10060 5828 10088 5856
rect 7984 5800 10088 5828
rect 10137 5831 10195 5837
rect 7984 5788 7990 5800
rect 10137 5797 10149 5831
rect 10183 5828 10195 5831
rect 10318 5828 10324 5840
rect 10183 5800 10324 5828
rect 10183 5797 10195 5800
rect 10137 5791 10195 5797
rect 10318 5788 10324 5800
rect 10376 5788 10382 5840
rect 10686 5788 10692 5840
rect 10744 5837 10750 5840
rect 10744 5831 10808 5837
rect 10744 5797 10762 5831
rect 10796 5797 10808 5831
rect 10744 5791 10808 5797
rect 10744 5788 10750 5791
rect 7374 5760 7380 5772
rect 5552 5732 5856 5760
rect 7335 5732 7380 5760
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 8205 5763 8263 5769
rect 8205 5729 8217 5763
rect 8251 5760 8263 5763
rect 8846 5760 8852 5772
rect 8251 5732 8852 5760
rect 8251 5729 8263 5732
rect 8205 5723 8263 5729
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 9033 5763 9091 5769
rect 9033 5729 9045 5763
rect 9079 5760 9091 5763
rect 9122 5760 9128 5772
rect 9079 5732 9128 5760
rect 9079 5729 9091 5732
rect 9033 5723 9091 5729
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 9398 5720 9404 5772
rect 9456 5760 9462 5772
rect 9858 5760 9864 5772
rect 9456 5732 9864 5760
rect 9456 5720 9462 5732
rect 9858 5720 9864 5732
rect 9916 5720 9922 5772
rect 10042 5720 10048 5772
rect 10100 5760 10106 5772
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 10100 5732 10517 5760
rect 10100 5720 10106 5732
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 5442 5692 5448 5704
rect 5403 5664 5448 5692
rect 4617 5655 4675 5661
rect 3418 5624 3424 5636
rect 3331 5596 3424 5624
rect 3418 5584 3424 5596
rect 3476 5624 3482 5636
rect 4632 5624 4660 5655
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7466 5692 7472 5704
rect 6972 5664 7472 5692
rect 6972 5652 6978 5664
rect 7466 5652 7472 5664
rect 7524 5692 7530 5704
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 7524 5664 7573 5692
rect 7524 5652 7530 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 8389 5695 8447 5701
rect 8389 5692 8401 5695
rect 7561 5655 7619 5661
rect 8220 5664 8401 5692
rect 8220 5636 8248 5664
rect 8389 5661 8401 5664
rect 8435 5661 8447 5695
rect 9306 5692 9312 5704
rect 9267 5664 9312 5692
rect 8389 5655 8447 5661
rect 9306 5652 9312 5664
rect 9364 5692 9370 5704
rect 9364 5664 9996 5692
rect 9364 5652 9370 5664
rect 3476 5596 4660 5624
rect 6825 5627 6883 5633
rect 3476 5584 3482 5596
rect 6825 5593 6837 5627
rect 6871 5624 6883 5627
rect 7006 5624 7012 5636
rect 6871 5596 7012 5624
rect 6871 5593 6883 5596
rect 6825 5587 6883 5593
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 8202 5584 8208 5636
rect 8260 5584 8266 5636
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 4985 5559 5043 5565
rect 4985 5556 4997 5559
rect 4764 5528 4997 5556
rect 4764 5516 4770 5528
rect 4985 5525 4997 5528
rect 5031 5556 5043 5559
rect 7742 5556 7748 5568
rect 5031 5528 7748 5556
rect 5031 5525 5043 5528
rect 4985 5519 5043 5525
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 9490 5556 9496 5568
rect 9180 5528 9496 5556
rect 9180 5516 9186 5528
rect 9490 5516 9496 5528
rect 9548 5556 9554 5568
rect 9861 5559 9919 5565
rect 9861 5556 9873 5559
rect 9548 5528 9873 5556
rect 9548 5516 9554 5528
rect 9861 5525 9873 5528
rect 9907 5525 9919 5559
rect 9968 5556 9996 5664
rect 11885 5559 11943 5565
rect 11885 5556 11897 5559
rect 9968 5528 11897 5556
rect 9861 5519 9919 5525
rect 11885 5525 11897 5528
rect 11931 5525 11943 5559
rect 11885 5519 11943 5525
rect 1104 5466 16008 5488
rect 1104 5414 3480 5466
rect 3532 5414 3544 5466
rect 3596 5414 3608 5466
rect 3660 5414 3672 5466
rect 3724 5414 8478 5466
rect 8530 5414 8542 5466
rect 8594 5414 8606 5466
rect 8658 5414 8670 5466
rect 8722 5414 13475 5466
rect 13527 5414 13539 5466
rect 13591 5414 13603 5466
rect 13655 5414 13667 5466
rect 13719 5414 16008 5466
rect 1104 5392 16008 5414
rect 5626 5352 5632 5364
rect 2056 5324 5632 5352
rect 2056 5157 2084 5324
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 5718 5312 5724 5364
rect 5776 5352 5782 5364
rect 6089 5355 6147 5361
rect 6089 5352 6101 5355
rect 5776 5324 6101 5352
rect 5776 5312 5782 5324
rect 6089 5321 6101 5324
rect 6135 5321 6147 5355
rect 6362 5352 6368 5364
rect 6323 5324 6368 5352
rect 6089 5315 6147 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 7524 5324 8217 5352
rect 7524 5312 7530 5324
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 8205 5315 8263 5321
rect 8389 5355 8447 5361
rect 8389 5321 8401 5355
rect 8435 5352 8447 5355
rect 8938 5352 8944 5364
rect 8435 5324 8944 5352
rect 8435 5321 8447 5324
rect 8389 5315 8447 5321
rect 6273 5287 6331 5293
rect 6273 5253 6285 5287
rect 6319 5284 6331 5287
rect 6822 5284 6828 5296
rect 6319 5256 6828 5284
rect 6319 5253 6331 5256
rect 6273 5247 6331 5253
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 2222 5216 2228 5228
rect 2183 5188 2228 5216
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 6730 5216 6736 5228
rect 6687 5188 6736 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 6730 5176 6736 5188
rect 6788 5216 6794 5228
rect 6788 5188 6960 5216
rect 6788 5176 6794 5188
rect 1489 5151 1547 5157
rect 1489 5117 1501 5151
rect 1535 5117 1547 5151
rect 1489 5111 1547 5117
rect 2041 5151 2099 5157
rect 2041 5117 2053 5151
rect 2087 5117 2099 5151
rect 2041 5111 2099 5117
rect 1504 5012 1532 5111
rect 2130 5108 2136 5160
rect 2188 5148 2194 5160
rect 2869 5151 2927 5157
rect 2869 5148 2881 5151
rect 2188 5120 2881 5148
rect 2188 5108 2194 5120
rect 2869 5117 2881 5120
rect 2915 5148 2927 5151
rect 4522 5148 4528 5160
rect 2915 5120 4384 5148
rect 4483 5120 4528 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 1762 5080 1768 5092
rect 1723 5052 1768 5080
rect 1762 5040 1768 5052
rect 1820 5040 1826 5092
rect 3136 5083 3194 5089
rect 3136 5049 3148 5083
rect 3182 5080 3194 5083
rect 4154 5080 4160 5092
rect 3182 5052 4160 5080
rect 3182 5049 3194 5052
rect 3136 5043 3194 5049
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 3326 5012 3332 5024
rect 1504 4984 3332 5012
rect 3326 4972 3332 4984
rect 3384 4972 3390 5024
rect 3970 4972 3976 5024
rect 4028 5012 4034 5024
rect 4356 5021 4384 5120
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 5442 5148 5448 5160
rect 4755 5120 5448 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 4249 5015 4307 5021
rect 4249 5012 4261 5015
rect 4028 4984 4261 5012
rect 4028 4972 4034 4984
rect 4249 4981 4261 4984
rect 4295 4981 4307 5015
rect 4249 4975 4307 4981
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 4724 5012 4752 5111
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 6822 5148 6828 5160
rect 6196 5120 6684 5148
rect 6783 5120 6828 5148
rect 4976 5083 5034 5089
rect 4976 5049 4988 5083
rect 5022 5080 5034 5083
rect 6196 5080 6224 5120
rect 5022 5052 6224 5080
rect 6656 5080 6684 5120
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 6932 5148 6960 5188
rect 8404 5148 8432 5315
rect 8938 5312 8944 5324
rect 8996 5352 9002 5364
rect 9490 5352 9496 5364
rect 8996 5324 9496 5352
rect 8996 5312 9002 5324
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 12066 5352 12072 5364
rect 9732 5324 12072 5352
rect 9732 5312 9738 5324
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 14826 5352 14832 5364
rect 14787 5324 14832 5352
rect 14826 5312 14832 5324
rect 14884 5312 14890 5364
rect 12342 5176 12348 5228
rect 12400 5216 12406 5228
rect 13081 5219 13139 5225
rect 13081 5216 13093 5219
rect 12400 5188 13093 5216
rect 12400 5176 12406 5188
rect 13081 5185 13093 5188
rect 13127 5216 13139 5219
rect 13354 5216 13360 5228
rect 13127 5188 13360 5216
rect 13127 5185 13139 5188
rect 13081 5179 13139 5185
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 6932 5120 8432 5148
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5148 8631 5151
rect 8840 5151 8898 5157
rect 8619 5120 8708 5148
rect 8619 5117 8631 5120
rect 8573 5111 8631 5117
rect 6914 5080 6920 5092
rect 6656 5052 6920 5080
rect 5022 5049 5034 5052
rect 4976 5043 5034 5049
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 7092 5083 7150 5089
rect 7092 5049 7104 5083
rect 7138 5080 7150 5083
rect 8202 5080 8208 5092
rect 7138 5052 8208 5080
rect 7138 5049 7150 5052
rect 7092 5043 7150 5049
rect 8202 5040 8208 5052
rect 8260 5080 8266 5092
rect 8680 5080 8708 5120
rect 8840 5117 8852 5151
rect 8886 5148 8898 5151
rect 9306 5148 9312 5160
rect 8886 5120 9312 5148
rect 8886 5117 8898 5120
rect 8840 5111 8898 5117
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 10042 5148 10048 5160
rect 9955 5120 10048 5148
rect 10042 5108 10048 5120
rect 10100 5148 10106 5160
rect 11330 5148 11336 5160
rect 10100 5120 11336 5148
rect 10100 5108 10106 5120
rect 11330 5108 11336 5120
rect 11388 5108 11394 5160
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12894 5148 12900 5160
rect 12492 5120 12900 5148
rect 12492 5108 12498 5120
rect 12894 5108 12900 5120
rect 12952 5148 12958 5160
rect 13541 5151 13599 5157
rect 13541 5148 13553 5151
rect 12952 5120 13553 5148
rect 12952 5108 12958 5120
rect 13541 5117 13553 5120
rect 13587 5117 13599 5151
rect 13541 5111 13599 5117
rect 14826 5108 14832 5160
rect 14884 5148 14890 5160
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 14884 5120 15025 5148
rect 14884 5108 14890 5120
rect 15013 5117 15025 5120
rect 15059 5117 15071 5151
rect 15013 5111 15071 5117
rect 9398 5080 9404 5092
rect 8260 5052 8616 5080
rect 8680 5052 9404 5080
rect 8260 5040 8266 5052
rect 8588 5024 8616 5052
rect 9398 5040 9404 5052
rect 9456 5080 9462 5092
rect 10060 5080 10088 5108
rect 10318 5089 10324 5092
rect 10312 5080 10324 5089
rect 9456 5052 10088 5080
rect 10279 5052 10324 5080
rect 9456 5040 9462 5052
rect 10312 5043 10324 5052
rect 10318 5040 10324 5043
rect 10376 5040 10382 5092
rect 12805 5083 12863 5089
rect 12805 5049 12817 5083
rect 12851 5080 12863 5083
rect 13265 5083 13323 5089
rect 13265 5080 13277 5083
rect 12851 5052 13277 5080
rect 12851 5049 12863 5052
rect 12805 5043 12863 5049
rect 13265 5049 13277 5052
rect 13311 5049 13323 5083
rect 13265 5043 13323 5049
rect 15289 5083 15347 5089
rect 15289 5049 15301 5083
rect 15335 5080 15347 5083
rect 16206 5080 16212 5092
rect 15335 5052 16212 5080
rect 15335 5049 15347 5052
rect 15289 5043 15347 5049
rect 16206 5040 16212 5052
rect 16264 5040 16270 5092
rect 4387 4984 4752 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 5258 4972 5264 5024
rect 5316 5012 5322 5024
rect 7006 5012 7012 5024
rect 5316 4984 7012 5012
rect 5316 4972 5322 4984
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 9953 5015 10011 5021
rect 9953 5012 9965 5015
rect 8628 4984 9965 5012
rect 8628 4972 8634 4984
rect 9953 4981 9965 4984
rect 9999 4981 10011 5015
rect 9953 4975 10011 4981
rect 10686 4972 10692 5024
rect 10744 5012 10750 5024
rect 11425 5015 11483 5021
rect 11425 5012 11437 5015
rect 10744 4984 11437 5012
rect 10744 4972 10750 4984
rect 11425 4981 11437 4984
rect 11471 4981 11483 5015
rect 11425 4975 11483 4981
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 12618 5012 12624 5024
rect 12483 4984 12624 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 1104 4922 16008 4944
rect 1104 4870 5979 4922
rect 6031 4870 6043 4922
rect 6095 4870 6107 4922
rect 6159 4870 6171 4922
rect 6223 4870 10976 4922
rect 11028 4870 11040 4922
rect 11092 4870 11104 4922
rect 11156 4870 11168 4922
rect 11220 4870 16008 4922
rect 1104 4848 16008 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3605 4811 3663 4817
rect 2832 4780 2877 4808
rect 2832 4768 2838 4780
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 4341 4811 4399 4817
rect 4341 4808 4353 4811
rect 3651 4780 4353 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 4341 4777 4353 4780
rect 4387 4777 4399 4811
rect 4798 4808 4804 4820
rect 4759 4780 4804 4808
rect 4341 4771 4399 4777
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 5169 4811 5227 4817
rect 5169 4777 5181 4811
rect 5215 4777 5227 4811
rect 5169 4771 5227 4777
rect 2130 4740 2136 4752
rect 1504 4712 2136 4740
rect 1504 4684 1532 4712
rect 2130 4700 2136 4712
rect 2188 4700 2194 4752
rect 3513 4743 3571 4749
rect 3513 4709 3525 4743
rect 3559 4740 3571 4743
rect 5184 4740 5212 4771
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 5629 4811 5687 4817
rect 5629 4808 5641 4811
rect 5316 4780 5641 4808
rect 5316 4768 5322 4780
rect 5629 4777 5641 4780
rect 5675 4808 5687 4811
rect 6270 4808 6276 4820
rect 5675 4780 6276 4808
rect 5675 4777 5687 4780
rect 5629 4771 5687 4777
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 6546 4808 6552 4820
rect 6507 4780 6552 4808
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 6641 4811 6699 4817
rect 6641 4777 6653 4811
rect 6687 4808 6699 4811
rect 7282 4808 7288 4820
rect 6687 4780 7288 4808
rect 6687 4777 6699 4780
rect 6641 4771 6699 4777
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 7374 4768 7380 4820
rect 7432 4808 7438 4820
rect 7929 4811 7987 4817
rect 7929 4808 7941 4811
rect 7432 4780 7941 4808
rect 7432 4768 7438 4780
rect 7929 4777 7941 4780
rect 7975 4777 7987 4811
rect 7929 4771 7987 4777
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 8389 4811 8447 4817
rect 8389 4808 8401 4811
rect 8352 4780 8401 4808
rect 8352 4768 8358 4780
rect 8389 4777 8401 4780
rect 8435 4777 8447 4811
rect 8389 4771 8447 4777
rect 8757 4811 8815 4817
rect 8757 4777 8769 4811
rect 8803 4808 8815 4811
rect 8846 4808 8852 4820
rect 8803 4780 8852 4808
rect 8803 4777 8815 4780
rect 8757 4771 8815 4777
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 9214 4808 9220 4820
rect 9175 4780 9220 4808
rect 9214 4768 9220 4780
rect 9272 4768 9278 4820
rect 9582 4768 9588 4820
rect 9640 4808 9646 4820
rect 9953 4811 10011 4817
rect 9953 4808 9965 4811
rect 9640 4780 9965 4808
rect 9640 4768 9646 4780
rect 9953 4777 9965 4780
rect 9999 4777 10011 4811
rect 9953 4771 10011 4777
rect 10229 4811 10287 4817
rect 10229 4777 10241 4811
rect 10275 4808 10287 4811
rect 11422 4808 11428 4820
rect 10275 4780 11428 4808
rect 10275 4777 10287 4780
rect 10229 4771 10287 4777
rect 9600 4740 9628 4768
rect 10134 4740 10140 4752
rect 3559 4712 5212 4740
rect 5368 4712 8248 4740
rect 3559 4709 3571 4712
rect 3513 4703 3571 4709
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1486 4672 1492 4684
rect 1443 4644 1492 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 1486 4632 1492 4644
rect 1544 4632 1550 4684
rect 1664 4675 1722 4681
rect 1664 4641 1676 4675
rect 1710 4672 1722 4675
rect 4246 4672 4252 4684
rect 1710 4644 3740 4672
rect 4207 4644 4252 4672
rect 1710 4641 1722 4644
rect 1664 4635 1722 4641
rect 3712 4613 3740 4644
rect 4246 4632 4252 4644
rect 4304 4672 4310 4684
rect 4709 4675 4767 4681
rect 4709 4672 4721 4675
rect 4304 4644 4721 4672
rect 4304 4632 4310 4644
rect 4709 4641 4721 4644
rect 4755 4672 4767 4675
rect 5368 4672 5396 4712
rect 5534 4672 5540 4684
rect 4755 4644 5396 4672
rect 5495 4644 5540 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 6089 4675 6147 4681
rect 6089 4641 6101 4675
rect 6135 4672 6147 4675
rect 6638 4672 6644 4684
rect 6135 4644 6644 4672
rect 6135 4641 6147 4644
rect 6089 4635 6147 4641
rect 6638 4632 6644 4644
rect 6696 4632 6702 4684
rect 7009 4675 7067 4681
rect 7009 4641 7021 4675
rect 7055 4672 7067 4675
rect 7834 4672 7840 4684
rect 7055 4644 7840 4672
rect 7055 4641 7067 4644
rect 7009 4635 7067 4641
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 3697 4607 3755 4613
rect 3697 4573 3709 4607
rect 3743 4604 3755 4607
rect 3970 4604 3976 4616
rect 3743 4576 3976 4604
rect 3743 4573 3755 4576
rect 3697 4567 3755 4573
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4154 4564 4160 4616
rect 4212 4564 4218 4616
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4573 7343 4607
rect 7466 4604 7472 4616
rect 7427 4576 7472 4604
rect 7285 4567 7343 4573
rect 4172 4536 4200 4564
rect 4908 4536 4936 4567
rect 4982 4536 4988 4548
rect 2976 4508 4016 4536
rect 4172 4508 4988 4536
rect 2682 4428 2688 4480
rect 2740 4468 2746 4480
rect 2976 4477 3004 4508
rect 2961 4471 3019 4477
rect 2961 4468 2973 4471
rect 2740 4440 2973 4468
rect 2740 4428 2746 4440
rect 2961 4437 2973 4440
rect 3007 4437 3019 4471
rect 3142 4468 3148 4480
rect 3103 4440 3148 4468
rect 2961 4431 3019 4437
rect 3142 4428 3148 4440
rect 3200 4428 3206 4480
rect 3988 4468 4016 4508
rect 4982 4496 4988 4508
rect 5040 4536 5046 4548
rect 5736 4536 5764 4567
rect 5040 4508 5764 4536
rect 5040 4496 5046 4508
rect 4614 4468 4620 4480
rect 3988 4440 4620 4468
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 6270 4468 6276 4480
rect 6231 4440 6276 4468
rect 6270 4428 6276 4440
rect 6328 4428 6334 4480
rect 7107 4468 7135 4567
rect 7300 4536 7328 4567
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 8220 4604 8248 4712
rect 8312 4712 9628 4740
rect 9784 4712 10140 4740
rect 8312 4681 8340 4712
rect 8297 4675 8355 4681
rect 8297 4641 8309 4675
rect 8343 4641 8355 4675
rect 9125 4675 9183 4681
rect 8297 4635 8355 4641
rect 8404 4644 8708 4672
rect 8404 4604 8432 4644
rect 8570 4604 8576 4616
rect 8220 4576 8432 4604
rect 8531 4576 8576 4604
rect 8570 4564 8576 4576
rect 8628 4564 8634 4616
rect 7650 4536 7656 4548
rect 7300 4508 7656 4536
rect 7650 4496 7656 4508
rect 7708 4536 7714 4548
rect 8588 4536 8616 4564
rect 7708 4508 8616 4536
rect 8680 4536 8708 4644
rect 9125 4641 9137 4675
rect 9171 4672 9183 4675
rect 9784 4672 9812 4712
rect 10134 4700 10140 4712
rect 10192 4740 10198 4752
rect 10244 4740 10272 4771
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 13173 4811 13231 4817
rect 13173 4808 13185 4811
rect 12768 4780 13185 4808
rect 12768 4768 12774 4780
rect 13173 4777 13185 4780
rect 13219 4808 13231 4811
rect 13446 4808 13452 4820
rect 13219 4780 13452 4808
rect 13219 4777 13231 4780
rect 13173 4771 13231 4777
rect 13446 4768 13452 4780
rect 13504 4808 13510 4820
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13504 4780 13645 4808
rect 13504 4768 13510 4780
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13633 4771 13691 4777
rect 13909 4811 13967 4817
rect 13909 4777 13921 4811
rect 13955 4808 13967 4811
rect 14734 4808 14740 4820
rect 13955 4780 14740 4808
rect 13955 4777 13967 4780
rect 13909 4771 13967 4777
rect 10192 4712 10272 4740
rect 10192 4700 10198 4712
rect 10318 4700 10324 4752
rect 10376 4740 10382 4752
rect 10376 4712 12756 4740
rect 10376 4700 10382 4712
rect 9171 4644 9812 4672
rect 9861 4675 9919 4681
rect 9171 4641 9183 4644
rect 9125 4635 9183 4641
rect 9861 4641 9873 4675
rect 9907 4672 9919 4675
rect 9950 4672 9956 4684
rect 9907 4644 9956 4672
rect 9907 4641 9919 4644
rect 9861 4635 9919 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10778 4672 10784 4684
rect 10739 4644 10784 4672
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 9306 4604 9312 4616
rect 9267 4576 9312 4604
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 10410 4604 10416 4616
rect 9640 4576 10416 4604
rect 9640 4564 9646 4576
rect 10410 4564 10416 4576
rect 10468 4564 10474 4616
rect 10870 4604 10876 4616
rect 10831 4576 10876 4604
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 10980 4613 11008 4712
rect 12728 4684 12756 4712
rect 12802 4700 12808 4752
rect 12860 4740 12866 4752
rect 13265 4743 13323 4749
rect 13265 4740 13277 4743
rect 12860 4712 13277 4740
rect 12860 4700 12866 4712
rect 13265 4709 13277 4712
rect 13311 4740 13323 4743
rect 13924 4740 13952 4771
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 13311 4712 13952 4740
rect 13311 4709 13323 4712
rect 13265 4703 13323 4709
rect 11330 4672 11336 4684
rect 11291 4644 11336 4672
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 11600 4675 11658 4681
rect 11600 4641 11612 4675
rect 11646 4672 11658 4675
rect 12342 4672 12348 4684
rect 11646 4644 12348 4672
rect 11646 4641 11658 4644
rect 11600 4635 11658 4641
rect 12342 4632 12348 4644
rect 12400 4632 12406 4684
rect 12710 4632 12716 4684
rect 12768 4632 12774 4684
rect 10965 4607 11023 4613
rect 10965 4573 10977 4607
rect 11011 4573 11023 4607
rect 10965 4567 11023 4573
rect 13354 4564 13360 4616
rect 13412 4604 13418 4616
rect 13412 4576 13457 4604
rect 13412 4564 13418 4576
rect 10318 4536 10324 4548
rect 8680 4508 10324 4536
rect 7708 4496 7714 4508
rect 10318 4496 10324 4508
rect 10376 4496 10382 4548
rect 13446 4496 13452 4548
rect 13504 4496 13510 4548
rect 7926 4468 7932 4480
rect 7107 4440 7932 4468
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 9398 4428 9404 4480
rect 9456 4468 9462 4480
rect 9677 4471 9735 4477
rect 9677 4468 9689 4471
rect 9456 4440 9689 4468
rect 9456 4428 9462 4440
rect 9677 4437 9689 4440
rect 9723 4437 9735 4471
rect 10410 4468 10416 4480
rect 10371 4440 10416 4468
rect 9677 4431 9735 4437
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 12710 4468 12716 4480
rect 12671 4440 12716 4468
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 12802 4428 12808 4480
rect 12860 4468 12866 4480
rect 12860 4440 12905 4468
rect 12860 4428 12866 4440
rect 13354 4428 13360 4480
rect 13412 4468 13418 4480
rect 13464 4468 13492 4496
rect 13412 4440 13492 4468
rect 13412 4428 13418 4440
rect 1104 4378 16008 4400
rect 1104 4326 3480 4378
rect 3532 4326 3544 4378
rect 3596 4326 3608 4378
rect 3660 4326 3672 4378
rect 3724 4326 8478 4378
rect 8530 4326 8542 4378
rect 8594 4326 8606 4378
rect 8658 4326 8670 4378
rect 8722 4326 13475 4378
rect 13527 4326 13539 4378
rect 13591 4326 13603 4378
rect 13655 4326 13667 4378
rect 13719 4326 16008 4378
rect 1104 4304 16008 4326
rect 2133 4267 2191 4273
rect 2133 4233 2145 4267
rect 2179 4264 2191 4267
rect 2498 4264 2504 4276
rect 2179 4236 2504 4264
rect 2179 4233 2191 4236
rect 2133 4227 2191 4233
rect 2498 4224 2504 4236
rect 2556 4224 2562 4276
rect 3326 4224 3332 4276
rect 3384 4264 3390 4276
rect 9953 4267 10011 4273
rect 9953 4264 9965 4267
rect 3384 4236 9965 4264
rect 3384 4224 3390 4236
rect 9953 4233 9965 4236
rect 9999 4233 10011 4267
rect 10778 4264 10784 4276
rect 10739 4236 10784 4264
rect 9953 4227 10011 4233
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 2409 4199 2467 4205
rect 2409 4165 2421 4199
rect 2455 4165 2467 4199
rect 2409 4159 2467 4165
rect 2424 4128 2452 4159
rect 2774 4156 2780 4208
rect 2832 4196 2838 4208
rect 2832 4168 3004 4196
rect 2832 4156 2838 4168
rect 2976 4137 3004 4168
rect 5534 4156 5540 4208
rect 5592 4156 5598 4208
rect 6362 4196 6368 4208
rect 5644 4168 6368 4196
rect 1504 4100 2452 4128
rect 2961 4131 3019 4137
rect 1504 4069 1532 4100
rect 2961 4097 2973 4131
rect 3007 4097 3019 4131
rect 3970 4128 3976 4140
rect 3931 4100 3976 4128
rect 2961 4091 3019 4097
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4982 4128 4988 4140
rect 4943 4100 4988 4128
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4128 5319 4131
rect 5552 4128 5580 4156
rect 5307 4100 5580 4128
rect 5307 4097 5319 4100
rect 5261 4091 5319 4097
rect 1489 4063 1547 4069
rect 1489 4029 1501 4063
rect 1535 4029 1547 4063
rect 1489 4023 1547 4029
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 3142 4060 3148 4072
rect 2823 4032 3148 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 3326 4060 3332 4072
rect 3287 4032 3332 4060
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4060 4399 4063
rect 5534 4060 5540 4072
rect 4387 4032 4844 4060
rect 5495 4032 5540 4060
rect 4387 4029 4399 4032
rect 4341 4023 4399 4029
rect 1765 3995 1823 4001
rect 1765 3961 1777 3995
rect 1811 3992 1823 3995
rect 2869 3995 2927 4001
rect 1811 3964 2820 3992
rect 1811 3961 1823 3964
rect 1765 3955 1823 3961
rect 2792 3936 2820 3964
rect 2869 3961 2881 3995
rect 2915 3992 2927 3995
rect 3789 3995 3847 4001
rect 2915 3964 3464 3992
rect 2915 3961 2927 3964
rect 2869 3955 2927 3961
rect 2317 3927 2375 3933
rect 2317 3893 2329 3927
rect 2363 3924 2375 3927
rect 2406 3924 2412 3936
rect 2363 3896 2412 3924
rect 2363 3893 2375 3896
rect 2317 3887 2375 3893
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 2774 3884 2780 3936
rect 2832 3884 2838 3936
rect 3436 3933 3464 3964
rect 3789 3961 3801 3995
rect 3835 3992 3847 3995
rect 3835 3964 4476 3992
rect 3835 3961 3847 3964
rect 3789 3955 3847 3961
rect 3421 3927 3479 3933
rect 3421 3893 3433 3927
rect 3467 3893 3479 3927
rect 3878 3924 3884 3936
rect 3839 3896 3884 3924
rect 3421 3887 3479 3893
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 4448 3933 4476 3964
rect 4816 3936 4844 4032
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 4433 3927 4491 3933
rect 4433 3893 4445 3927
rect 4479 3893 4491 3927
rect 4798 3924 4804 3936
rect 4759 3896 4804 3924
rect 4433 3887 4491 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 4893 3927 4951 3933
rect 4893 3893 4905 3927
rect 4939 3924 4951 3927
rect 5350 3924 5356 3936
rect 4939 3896 5356 3924
rect 4939 3893 4951 3896
rect 4893 3887 4951 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 5644 3924 5672 4168
rect 6362 4156 6368 4168
rect 6420 4156 6426 4208
rect 7650 4196 7656 4208
rect 7484 4168 7656 4196
rect 6454 4128 6460 4140
rect 6415 4100 6460 4128
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 7484 4137 7512 4168
rect 7650 4156 7656 4168
rect 7708 4156 7714 4208
rect 8754 4156 8760 4208
rect 8812 4196 8818 4208
rect 9861 4199 9919 4205
rect 9861 4196 9873 4199
rect 8812 4168 9873 4196
rect 8812 4156 8818 4168
rect 9861 4165 9873 4168
rect 9907 4196 9919 4199
rect 10226 4196 10232 4208
rect 9907 4168 10232 4196
rect 9907 4165 9919 4168
rect 9861 4159 9919 4165
rect 10226 4156 10232 4168
rect 10284 4156 10290 4208
rect 10686 4196 10692 4208
rect 10612 4168 10692 4196
rect 7285 4131 7343 4137
rect 7285 4128 7297 4131
rect 6788 4100 7297 4128
rect 6788 4088 6794 4100
rect 7285 4097 7297 4100
rect 7331 4097 7343 4131
rect 7285 4091 7343 4097
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 8260 4100 8401 4128
rect 8260 4088 8266 4100
rect 8389 4097 8401 4100
rect 8435 4128 8447 4131
rect 9125 4131 9183 4137
rect 9125 4128 9137 4131
rect 8435 4100 9137 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 9125 4097 9137 4100
rect 9171 4097 9183 4131
rect 10410 4128 10416 4140
rect 10371 4100 10416 4128
rect 9125 4091 9183 4097
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 10612 4137 10640 4168
rect 10686 4156 10692 4168
rect 10744 4156 10750 4208
rect 12710 4156 12716 4208
rect 12768 4196 12774 4208
rect 12768 4168 13032 4196
rect 12768 4156 12774 4168
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4097 10655 4131
rect 11422 4128 11428 4140
rect 11335 4100 11428 4128
rect 10597 4091 10655 4097
rect 11422 4088 11428 4100
rect 11480 4128 11486 4140
rect 12342 4128 12348 4140
rect 11480 4100 12348 4128
rect 11480 4088 11486 4100
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 12802 4088 12808 4140
rect 12860 4128 12866 4140
rect 13004 4137 13032 4168
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12860 4100 12909 4128
rect 12860 4088 12866 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 12989 4091 13047 4097
rect 6362 4060 6368 4072
rect 5736 4032 6368 4060
rect 5736 3933 5764 4032
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4060 7251 4063
rect 7374 4060 7380 4072
rect 7239 4032 7380 4060
rect 7239 4029 7251 4032
rect 7193 4023 7251 4029
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 9030 4060 9036 4072
rect 7484 4032 9036 4060
rect 5994 3952 6000 4004
rect 6052 3992 6058 4004
rect 6273 3995 6331 4001
rect 6273 3992 6285 3995
rect 6052 3964 6285 3992
rect 6052 3952 6058 3964
rect 6273 3961 6285 3964
rect 6319 3992 6331 3995
rect 7484 3992 7512 4032
rect 9030 4020 9036 4032
rect 9088 4060 9094 4072
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9088 4032 9689 4060
rect 9088 4020 9094 4032
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 11149 4063 11207 4069
rect 11149 4060 11161 4063
rect 10008 4032 11161 4060
rect 10008 4020 10014 4032
rect 11149 4029 11161 4032
rect 11195 4060 11207 4063
rect 12066 4060 12072 4072
rect 11195 4032 12072 4060
rect 11195 4029 11207 4032
rect 11149 4023 11207 4029
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 8205 3995 8263 4001
rect 8205 3992 8217 3995
rect 6319 3964 7512 3992
rect 7576 3964 8217 3992
rect 6319 3961 6331 3964
rect 6273 3955 6331 3961
rect 5592 3896 5672 3924
rect 5721 3927 5779 3933
rect 5592 3884 5598 3896
rect 5721 3893 5733 3927
rect 5767 3893 5779 3927
rect 5721 3887 5779 3893
rect 5810 3884 5816 3936
rect 5868 3924 5874 3936
rect 5905 3927 5963 3933
rect 5905 3924 5917 3927
rect 5868 3896 5917 3924
rect 5868 3884 5874 3896
rect 5905 3893 5917 3896
rect 5951 3893 5963 3927
rect 5905 3887 5963 3893
rect 6365 3927 6423 3933
rect 6365 3893 6377 3927
rect 6411 3924 6423 3927
rect 6546 3924 6552 3936
rect 6411 3896 6552 3924
rect 6411 3893 6423 3896
rect 6365 3887 6423 3893
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 6825 3927 6883 3933
rect 6825 3893 6837 3927
rect 6871 3924 6883 3927
rect 7190 3924 7196 3936
rect 6871 3896 7196 3924
rect 6871 3893 6883 3896
rect 6825 3887 6883 3893
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7576 3924 7604 3964
rect 8205 3961 8217 3964
rect 8251 3961 8263 3995
rect 8205 3955 8263 3961
rect 10321 3995 10379 4001
rect 10321 3961 10333 3995
rect 10367 3992 10379 3995
rect 10367 3964 12480 3992
rect 10367 3961 10379 3964
rect 10321 3955 10379 3961
rect 7742 3924 7748 3936
rect 7340 3896 7604 3924
rect 7703 3896 7748 3924
rect 7340 3884 7346 3896
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 8573 3927 8631 3933
rect 8573 3924 8585 3927
rect 8352 3896 8585 3924
rect 8352 3884 8358 3896
rect 8573 3893 8585 3896
rect 8619 3893 8631 3927
rect 8938 3924 8944 3936
rect 8899 3896 8944 3924
rect 8573 3887 8631 3893
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9030 3884 9036 3936
rect 9088 3924 9094 3936
rect 9088 3896 9133 3924
rect 9088 3884 9094 3896
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9401 3927 9459 3933
rect 9401 3924 9413 3927
rect 9272 3896 9413 3924
rect 9272 3884 9278 3896
rect 9401 3893 9413 3896
rect 9447 3893 9459 3927
rect 9401 3887 9459 3893
rect 10502 3884 10508 3936
rect 10560 3924 10566 3936
rect 10686 3924 10692 3936
rect 10560 3896 10692 3924
rect 10560 3884 10566 3896
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 11241 3927 11299 3933
rect 11241 3893 11253 3927
rect 11287 3924 11299 3927
rect 11514 3924 11520 3936
rect 11287 3896 11520 3924
rect 11287 3893 11299 3896
rect 11241 3887 11299 3893
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 11701 3927 11759 3933
rect 11701 3893 11713 3927
rect 11747 3924 11759 3927
rect 12066 3924 12072 3936
rect 11747 3896 12072 3924
rect 11747 3893 11759 3896
rect 11701 3887 11759 3893
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 12452 3933 12480 3964
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 12805 3995 12863 4001
rect 12805 3992 12817 3995
rect 12676 3964 12817 3992
rect 12676 3952 12682 3964
rect 12805 3961 12817 3964
rect 12851 3961 12863 3995
rect 12805 3955 12863 3961
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3893 12495 3927
rect 12437 3887 12495 3893
rect 1104 3834 16008 3856
rect 1104 3782 5979 3834
rect 6031 3782 6043 3834
rect 6095 3782 6107 3834
rect 6159 3782 6171 3834
rect 6223 3782 10976 3834
rect 11028 3782 11040 3834
rect 11092 3782 11104 3834
rect 11156 3782 11168 3834
rect 11220 3782 16008 3834
rect 1104 3760 16008 3782
rect 2593 3723 2651 3729
rect 2593 3689 2605 3723
rect 2639 3720 2651 3723
rect 3234 3720 3240 3732
rect 2639 3692 3240 3720
rect 2639 3689 2651 3692
rect 2593 3683 2651 3689
rect 3234 3680 3240 3692
rect 3292 3680 3298 3732
rect 3697 3723 3755 3729
rect 3697 3689 3709 3723
rect 3743 3720 3755 3723
rect 5258 3720 5264 3732
rect 3743 3692 5264 3720
rect 3743 3689 3755 3692
rect 3697 3683 3755 3689
rect 5258 3680 5264 3692
rect 5316 3720 5322 3732
rect 5316 3692 5387 3720
rect 5316 3680 5322 3692
rect 3881 3655 3939 3661
rect 3881 3621 3893 3655
rect 3927 3652 3939 3655
rect 4430 3652 4436 3664
rect 3927 3624 4436 3652
rect 3927 3621 3939 3624
rect 3881 3615 3939 3621
rect 4430 3612 4436 3624
rect 4488 3612 4494 3664
rect 1489 3587 1547 3593
rect 1489 3553 1501 3587
rect 1535 3584 1547 3587
rect 1854 3584 1860 3596
rect 1535 3556 1860 3584
rect 1535 3553 1547 3556
rect 1489 3547 1547 3553
rect 1854 3544 1860 3556
rect 1912 3544 1918 3596
rect 2041 3587 2099 3593
rect 2041 3553 2053 3587
rect 2087 3584 2099 3587
rect 2406 3584 2412 3596
rect 2087 3556 2412 3584
rect 2087 3553 2099 3556
rect 2041 3547 2099 3553
rect 2406 3544 2412 3556
rect 2464 3544 2470 3596
rect 3050 3584 3056 3596
rect 3011 3556 3056 3584
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4522 3584 4528 3596
rect 4387 3556 4528 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3553 4859 3587
rect 4801 3547 4859 3553
rect 4893 3587 4951 3593
rect 4893 3553 4905 3587
rect 4939 3584 4951 3587
rect 5267 3587 5325 3593
rect 4939 3556 5212 3584
rect 4939 3553 4951 3556
rect 4893 3547 4951 3553
rect 1670 3516 1676 3528
rect 1631 3488 1676 3516
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 2774 3476 2780 3528
rect 2832 3476 2838 3528
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3516 3019 3519
rect 3142 3516 3148 3528
rect 3007 3488 3148 3516
rect 3007 3485 3019 3488
rect 2961 3479 3019 3485
rect 3142 3476 3148 3488
rect 3200 3476 3206 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3516 4215 3519
rect 4706 3516 4712 3528
rect 4203 3488 4712 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 2409 3451 2467 3457
rect 2409 3448 2421 3451
rect 2004 3420 2421 3448
rect 2004 3408 2010 3420
rect 2409 3417 2421 3420
rect 2455 3448 2467 3451
rect 2593 3451 2651 3457
rect 2593 3448 2605 3451
rect 2455 3420 2605 3448
rect 2455 3417 2467 3420
rect 2409 3411 2467 3417
rect 2593 3417 2605 3420
rect 2639 3417 2651 3451
rect 2792 3448 2820 3476
rect 3237 3451 3295 3457
rect 3237 3448 3249 3451
rect 2792 3420 3249 3448
rect 2593 3411 2651 3417
rect 3237 3417 3249 3420
rect 3283 3417 3295 3451
rect 3237 3411 3295 3417
rect 3513 3451 3571 3457
rect 3513 3417 3525 3451
rect 3559 3448 3571 3451
rect 4816 3448 4844 3547
rect 5184 3528 5212 3556
rect 5267 3553 5279 3587
rect 5313 3584 5325 3587
rect 5359 3584 5387 3692
rect 5810 3680 5816 3732
rect 5868 3720 5874 3732
rect 7561 3723 7619 3729
rect 7561 3720 7573 3723
rect 5868 3692 7573 3720
rect 5868 3680 5874 3692
rect 7561 3689 7573 3692
rect 7607 3689 7619 3723
rect 7561 3683 7619 3689
rect 7926 3680 7932 3732
rect 7984 3720 7990 3732
rect 8754 3720 8760 3732
rect 7984 3692 8760 3720
rect 7984 3680 7990 3692
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 9677 3723 9735 3729
rect 9677 3720 9689 3723
rect 8904 3692 9689 3720
rect 8904 3680 8910 3692
rect 9677 3689 9689 3692
rect 9723 3689 9735 3723
rect 10134 3720 10140 3732
rect 10095 3692 10140 3720
rect 9677 3683 9735 3689
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10689 3723 10747 3729
rect 10689 3689 10701 3723
rect 10735 3720 10747 3723
rect 10870 3720 10876 3732
rect 10735 3692 10876 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 11330 3680 11336 3732
rect 11388 3680 11394 3732
rect 11606 3680 11612 3732
rect 11664 3720 11670 3732
rect 11790 3720 11796 3732
rect 11664 3692 11796 3720
rect 11664 3680 11670 3692
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12342 3680 12348 3732
rect 12400 3720 12406 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 12400 3692 12909 3720
rect 12400 3680 12406 3692
rect 12897 3689 12909 3692
rect 12943 3689 12955 3723
rect 12897 3683 12955 3689
rect 5896 3655 5954 3661
rect 5896 3621 5908 3655
rect 5942 3652 5954 3655
rect 6454 3652 6460 3664
rect 5942 3624 6460 3652
rect 5942 3621 5954 3624
rect 5896 3615 5954 3621
rect 6454 3612 6460 3624
rect 6512 3612 6518 3664
rect 7466 3652 7472 3664
rect 7427 3624 7472 3652
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 7650 3652 7656 3664
rect 7576 3624 7656 3652
rect 5313 3556 5387 3584
rect 5313 3553 5325 3556
rect 5267 3547 5325 3553
rect 7190 3544 7196 3596
rect 7248 3584 7254 3596
rect 7576 3584 7604 3624
rect 7650 3612 7656 3624
rect 7708 3612 7714 3664
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 8358 3655 8416 3661
rect 8358 3652 8370 3655
rect 8260 3624 8370 3652
rect 8260 3612 8266 3624
rect 8358 3621 8370 3624
rect 8404 3621 8416 3655
rect 8358 3615 8416 3621
rect 9490 3612 9496 3664
rect 9548 3652 9554 3664
rect 9861 3655 9919 3661
rect 9861 3652 9873 3655
rect 9548 3624 9873 3652
rect 9548 3612 9554 3624
rect 9861 3621 9873 3624
rect 9907 3621 9919 3655
rect 11348 3652 11376 3680
rect 11348 3624 11560 3652
rect 9861 3615 9919 3621
rect 8113 3587 8171 3593
rect 8113 3584 8125 3587
rect 7248 3556 7604 3584
rect 7668 3556 8125 3584
rect 7248 3544 7254 3556
rect 5074 3516 5080 3528
rect 5035 3488 5080 3516
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 5166 3476 5172 3528
rect 5224 3476 5230 3528
rect 5442 3476 5448 3528
rect 5500 3516 5506 3528
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 5500 3488 5641 3516
rect 5500 3476 5506 3488
rect 5629 3485 5641 3488
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 7668 3516 7696 3556
rect 8113 3553 8125 3556
rect 8159 3584 8171 3587
rect 9398 3584 9404 3596
rect 8159 3556 9404 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 10870 3584 10876 3596
rect 9824 3556 10876 3584
rect 9824 3544 9830 3556
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 11330 3584 11336 3596
rect 11103 3556 11336 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 11330 3544 11336 3556
rect 11388 3544 11394 3596
rect 11532 3593 11560 3624
rect 12618 3612 12624 3664
rect 12676 3652 12682 3664
rect 13078 3652 13084 3664
rect 12676 3624 13084 3652
rect 12676 3612 12682 3624
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 11517 3587 11575 3593
rect 11517 3553 11529 3587
rect 11563 3553 11575 3587
rect 11517 3547 11575 3553
rect 11606 3544 11612 3596
rect 11664 3584 11670 3596
rect 11773 3587 11831 3593
rect 11773 3584 11785 3587
rect 11664 3556 11785 3584
rect 11664 3544 11670 3556
rect 11773 3553 11785 3556
rect 11819 3553 11831 3587
rect 11773 3547 11831 3553
rect 7064 3488 7696 3516
rect 7745 3519 7803 3525
rect 7064 3476 7070 3488
rect 7745 3485 7757 3519
rect 7791 3516 7803 3519
rect 7834 3516 7840 3528
rect 7791 3488 7840 3516
rect 7791 3485 7803 3488
rect 7745 3479 7803 3485
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 9640 3488 10425 3516
rect 9640 3476 9646 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 11149 3519 11207 3525
rect 11149 3516 11161 3519
rect 11020 3488 11161 3516
rect 11020 3476 11026 3488
rect 11149 3485 11161 3488
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 11241 3519 11299 3525
rect 11241 3485 11253 3519
rect 11287 3516 11299 3519
rect 11422 3516 11428 3528
rect 11287 3488 11428 3516
rect 11287 3485 11299 3488
rect 11241 3479 11299 3485
rect 11422 3476 11428 3488
rect 11480 3476 11486 3528
rect 7101 3451 7159 3457
rect 3559 3420 5672 3448
rect 3559 3417 3571 3420
rect 3513 3411 3571 3417
rect 1394 3340 1400 3392
rect 1452 3380 1458 3392
rect 2225 3383 2283 3389
rect 2225 3380 2237 3383
rect 1452 3352 2237 3380
rect 1452 3340 1458 3352
rect 2225 3349 2237 3352
rect 2271 3349 2283 3383
rect 2225 3343 2283 3349
rect 2314 3340 2320 3392
rect 2372 3380 2378 3392
rect 2777 3383 2835 3389
rect 2777 3380 2789 3383
rect 2372 3352 2789 3380
rect 2372 3340 2378 3352
rect 2777 3349 2789 3352
rect 2823 3380 2835 3383
rect 3528 3380 3556 3411
rect 4430 3380 4436 3392
rect 2823 3352 3556 3380
rect 4391 3352 4436 3380
rect 2823 3349 2835 3352
rect 2777 3343 2835 3349
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 4706 3340 4712 3392
rect 4764 3380 4770 3392
rect 5258 3380 5264 3392
rect 4764 3352 5264 3380
rect 4764 3340 4770 3352
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5445 3383 5503 3389
rect 5445 3349 5457 3383
rect 5491 3380 5503 3383
rect 5534 3380 5540 3392
rect 5491 3352 5540 3380
rect 5491 3349 5503 3352
rect 5445 3343 5503 3349
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 5644 3380 5672 3420
rect 7101 3417 7113 3451
rect 7147 3448 7159 3451
rect 7282 3448 7288 3460
rect 7147 3420 7288 3448
rect 7147 3417 7159 3420
rect 7101 3411 7159 3417
rect 7282 3408 7288 3420
rect 7340 3408 7346 3460
rect 7466 3408 7472 3460
rect 7524 3448 7530 3460
rect 7650 3448 7656 3460
rect 7524 3420 7656 3448
rect 7524 3408 7530 3420
rect 7650 3408 7656 3420
rect 7708 3448 7714 3460
rect 7929 3451 7987 3457
rect 7929 3448 7941 3451
rect 7708 3420 7941 3448
rect 7708 3408 7714 3420
rect 7929 3417 7941 3420
rect 7975 3417 7987 3451
rect 7929 3411 7987 3417
rect 6546 3380 6552 3392
rect 5644 3352 6552 3380
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 7009 3383 7067 3389
rect 7009 3349 7021 3383
rect 7055 3380 7067 3383
rect 7374 3380 7380 3392
rect 7055 3352 7380 3380
rect 7055 3349 7067 3352
rect 7009 3343 7067 3349
rect 7374 3340 7380 3352
rect 7432 3380 7438 3392
rect 7834 3380 7840 3392
rect 7432 3352 7840 3380
rect 7432 3340 7438 3352
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 7944 3380 7972 3411
rect 9214 3380 9220 3392
rect 7944 3352 9220 3380
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 9490 3380 9496 3392
rect 9451 3352 9496 3380
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 9858 3340 9864 3392
rect 9916 3380 9922 3392
rect 10321 3383 10379 3389
rect 10321 3380 10333 3383
rect 9916 3352 10333 3380
rect 9916 3340 9922 3352
rect 10321 3349 10333 3352
rect 10367 3380 10379 3383
rect 11698 3380 11704 3392
rect 10367 3352 11704 3380
rect 10367 3349 10379 3352
rect 10321 3343 10379 3349
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 1104 3290 16008 3312
rect 1104 3238 3480 3290
rect 3532 3238 3544 3290
rect 3596 3238 3608 3290
rect 3660 3238 3672 3290
rect 3724 3238 8478 3290
rect 8530 3238 8542 3290
rect 8594 3238 8606 3290
rect 8658 3238 8670 3290
rect 8722 3238 13475 3290
rect 13527 3238 13539 3290
rect 13591 3238 13603 3290
rect 13655 3238 13667 3290
rect 13719 3238 16008 3290
rect 1104 3216 16008 3238
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 4433 3179 4491 3185
rect 3292 3148 4016 3176
rect 3292 3136 3298 3148
rect 3988 3108 4016 3148
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 4706 3176 4712 3188
rect 4479 3148 4712 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 4706 3136 4712 3148
rect 4764 3176 4770 3188
rect 4982 3176 4988 3188
rect 4764 3148 4988 3176
rect 4764 3136 4770 3148
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 5350 3176 5356 3188
rect 5311 3148 5356 3176
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 6454 3176 6460 3188
rect 5868 3148 6460 3176
rect 5868 3136 5874 3148
rect 6454 3136 6460 3148
rect 6512 3136 6518 3188
rect 6641 3179 6699 3185
rect 6641 3145 6653 3179
rect 6687 3176 6699 3179
rect 6822 3176 6828 3188
rect 6687 3148 6828 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 6822 3136 6828 3148
rect 6880 3176 6886 3188
rect 8018 3176 8024 3188
rect 6880 3148 8024 3176
rect 6880 3136 6886 3148
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8297 3179 8355 3185
rect 8297 3176 8309 3179
rect 8168 3148 8309 3176
rect 8168 3136 8174 3148
rect 8297 3145 8309 3148
rect 8343 3145 8355 3179
rect 8297 3139 8355 3145
rect 9122 3136 9128 3188
rect 9180 3176 9186 3188
rect 9217 3179 9275 3185
rect 9217 3176 9229 3179
rect 9180 3148 9229 3176
rect 9180 3136 9186 3148
rect 9217 3145 9229 3148
rect 9263 3145 9275 3179
rect 10962 3176 10968 3188
rect 10923 3148 10968 3176
rect 9217 3139 9275 3145
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 11514 3136 11520 3188
rect 11572 3176 11578 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 11572 3148 12449 3176
rect 11572 3136 11578 3148
rect 12437 3145 12449 3148
rect 12483 3145 12495 3179
rect 12437 3139 12495 3145
rect 4798 3108 4804 3120
rect 3988 3080 4804 3108
rect 4798 3068 4804 3080
rect 4856 3068 4862 3120
rect 4890 3068 4896 3120
rect 4948 3108 4954 3120
rect 6365 3111 6423 3117
rect 6365 3108 6377 3111
rect 4948 3080 6377 3108
rect 4948 3068 4954 3080
rect 6365 3077 6377 3080
rect 6411 3077 6423 3111
rect 8202 3108 8208 3120
rect 8163 3080 8208 3108
rect 6365 3071 6423 3077
rect 8202 3068 8208 3080
rect 8260 3068 8266 3120
rect 8570 3068 8576 3120
rect 8628 3108 8634 3120
rect 9030 3108 9036 3120
rect 8628 3080 9036 3108
rect 8628 3068 8634 3080
rect 9030 3068 9036 3080
rect 9088 3068 9094 3120
rect 10781 3111 10839 3117
rect 10781 3077 10793 3111
rect 10827 3108 10839 3111
rect 10827 3080 11560 3108
rect 10827 3077 10839 3080
rect 10781 3071 10839 3077
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 5074 3040 5080 3052
rect 1544 3012 1624 3040
rect 1544 3000 1550 3012
rect 1596 2981 1624 3012
rect 4816 3012 5080 3040
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2972 1639 2975
rect 3053 2975 3111 2981
rect 3053 2972 3065 2975
rect 1627 2944 3065 2972
rect 1627 2941 1639 2944
rect 1581 2935 1639 2941
rect 3053 2941 3065 2944
rect 3099 2941 3111 2975
rect 4816 2972 4844 3012
rect 5074 3000 5080 3012
rect 5132 3040 5138 3052
rect 5905 3043 5963 3049
rect 5905 3040 5917 3043
rect 5132 3012 5917 3040
rect 5132 3000 5138 3012
rect 5905 3009 5917 3012
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 6454 3000 6460 3052
rect 6512 3000 6518 3052
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3040 6883 3043
rect 6871 3012 6960 3040
rect 6871 3009 6883 3012
rect 6825 3003 6883 3009
rect 3053 2935 3111 2941
rect 3344 2944 4844 2972
rect 4985 2975 5043 2981
rect 1486 2904 1492 2916
rect 1399 2876 1492 2904
rect 1486 2864 1492 2876
rect 1544 2904 1550 2916
rect 3344 2913 3372 2944
rect 4985 2941 4997 2975
rect 5031 2972 5043 2975
rect 5810 2972 5816 2984
rect 5031 2944 5816 2972
rect 5031 2941 5043 2944
rect 4985 2935 5043 2941
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 6178 2972 6184 2984
rect 6139 2944 6184 2972
rect 6178 2932 6184 2944
rect 6236 2932 6242 2984
rect 6472 2972 6500 3000
rect 6730 2972 6736 2984
rect 6472 2944 6736 2972
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 1826 2907 1884 2913
rect 1826 2904 1838 2907
rect 1544 2876 1838 2904
rect 1544 2864 1550 2876
rect 1826 2873 1838 2876
rect 1872 2873 1884 2907
rect 3298 2907 3372 2913
rect 3298 2904 3310 2907
rect 1826 2867 1884 2873
rect 2976 2876 3310 2904
rect 2976 2845 3004 2876
rect 3298 2873 3310 2876
rect 3344 2876 3372 2907
rect 6454 2904 6460 2916
rect 3436 2876 6460 2904
rect 3344 2873 3356 2876
rect 3298 2867 3356 2873
rect 2961 2839 3019 2845
rect 2961 2805 2973 2839
rect 3007 2805 3019 2839
rect 2961 2799 3019 2805
rect 3142 2796 3148 2848
rect 3200 2836 3206 2848
rect 3436 2836 3464 2876
rect 6454 2864 6460 2876
rect 6512 2864 6518 2916
rect 6932 2904 6960 3012
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 7892 3012 8861 3040
rect 7892 3000 7898 3012
rect 8849 3009 8861 3012
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 8956 3012 9352 3040
rect 7092 2975 7150 2981
rect 7092 2941 7104 2975
rect 7138 2972 7150 2975
rect 7374 2972 7380 2984
rect 7138 2944 7380 2972
rect 7138 2941 7150 2944
rect 7092 2935 7150 2941
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 8956 2972 8984 3012
rect 7484 2944 8984 2972
rect 9324 2972 9352 3012
rect 9398 3000 9404 3052
rect 9456 3040 9462 3052
rect 11532 3049 11560 3080
rect 11517 3043 11575 3049
rect 9456 3012 9501 3040
rect 9456 3000 9462 3012
rect 11517 3009 11529 3043
rect 11563 3040 11575 3043
rect 11606 3040 11612 3052
rect 11563 3012 11612 3040
rect 11563 3009 11575 3012
rect 11517 3003 11575 3009
rect 11606 3000 11612 3012
rect 11664 3040 11670 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 11664 3012 13001 3040
rect 11664 3000 11670 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3040 14611 3043
rect 16942 3040 16948 3052
rect 14599 3012 16948 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 16942 3000 16948 3012
rect 17000 3000 17006 3052
rect 9950 2972 9956 2984
rect 9324 2944 9956 2972
rect 7006 2904 7012 2916
rect 6932 2876 7012 2904
rect 7006 2864 7012 2876
rect 7064 2864 7070 2916
rect 7190 2864 7196 2916
rect 7248 2904 7254 2916
rect 7484 2904 7512 2944
rect 9950 2932 9956 2944
rect 10008 2932 10014 2984
rect 14274 2972 14280 2984
rect 14235 2944 14280 2972
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 14642 2932 14648 2984
rect 14700 2972 14706 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14700 2944 14841 2972
rect 14700 2932 14706 2944
rect 14829 2941 14841 2944
rect 14875 2972 14887 2975
rect 15381 2975 15439 2981
rect 15381 2972 15393 2975
rect 14875 2944 15393 2972
rect 14875 2941 14887 2944
rect 14829 2935 14887 2941
rect 15381 2941 15393 2944
rect 15427 2941 15439 2975
rect 15381 2935 15439 2941
rect 8662 2904 8668 2916
rect 7248 2876 7512 2904
rect 8623 2876 8668 2904
rect 7248 2864 7254 2876
rect 8662 2864 8668 2876
rect 8720 2864 8726 2916
rect 8846 2864 8852 2916
rect 8904 2904 8910 2916
rect 9490 2904 9496 2916
rect 8904 2876 9496 2904
rect 8904 2864 8910 2876
rect 9490 2864 9496 2876
rect 9548 2904 9554 2916
rect 9646 2907 9704 2913
rect 9646 2904 9658 2907
rect 9548 2876 9658 2904
rect 9548 2864 9554 2876
rect 9646 2873 9658 2876
rect 9692 2873 9704 2907
rect 9646 2867 9704 2873
rect 9766 2864 9772 2916
rect 9824 2904 9830 2916
rect 11425 2907 11483 2913
rect 11425 2904 11437 2907
rect 9824 2876 11437 2904
rect 9824 2864 9830 2876
rect 11425 2873 11437 2876
rect 11471 2904 11483 2907
rect 11793 2907 11851 2913
rect 11793 2904 11805 2907
rect 11471 2876 11805 2904
rect 11471 2873 11483 2876
rect 11425 2867 11483 2873
rect 11793 2873 11805 2876
rect 11839 2873 11851 2907
rect 12158 2904 12164 2916
rect 12119 2876 12164 2904
rect 11793 2867 11851 2873
rect 12158 2864 12164 2876
rect 12216 2904 12222 2916
rect 12897 2907 12955 2913
rect 12897 2904 12909 2907
rect 12216 2876 12909 2904
rect 12216 2864 12222 2876
rect 12897 2873 12909 2876
rect 12943 2873 12955 2907
rect 12897 2867 12955 2873
rect 3200 2808 3464 2836
rect 3200 2796 3206 2808
rect 4522 2796 4528 2848
rect 4580 2836 4586 2848
rect 4580 2808 4625 2836
rect 4580 2796 4586 2808
rect 4798 2796 4804 2848
rect 4856 2836 4862 2848
rect 4893 2839 4951 2845
rect 4893 2836 4905 2839
rect 4856 2808 4905 2836
rect 4856 2796 4862 2808
rect 4893 2805 4905 2808
rect 4939 2805 4951 2839
rect 4893 2799 4951 2805
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 5721 2839 5779 2845
rect 5721 2836 5733 2839
rect 5500 2808 5733 2836
rect 5500 2796 5506 2808
rect 5721 2805 5733 2808
rect 5767 2805 5779 2839
rect 5721 2799 5779 2805
rect 5813 2839 5871 2845
rect 5813 2805 5825 2839
rect 5859 2836 5871 2839
rect 6822 2836 6828 2848
rect 5859 2808 6828 2836
rect 5859 2805 5871 2808
rect 5813 2799 5871 2805
rect 6822 2796 6828 2808
rect 6880 2796 6886 2848
rect 8754 2836 8760 2848
rect 8667 2808 8760 2836
rect 8754 2796 8760 2808
rect 8812 2836 8818 2848
rect 10226 2836 10232 2848
rect 8812 2808 10232 2836
rect 8812 2796 8818 2808
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 11333 2839 11391 2845
rect 11333 2805 11345 2839
rect 11379 2836 11391 2839
rect 11977 2839 12035 2845
rect 11977 2836 11989 2839
rect 11379 2808 11989 2836
rect 11379 2805 11391 2808
rect 11333 2799 11391 2805
rect 11977 2805 11989 2808
rect 12023 2836 12035 2839
rect 12250 2836 12256 2848
rect 12023 2808 12256 2836
rect 12023 2805 12035 2808
rect 11977 2799 12035 2805
rect 12250 2796 12256 2808
rect 12308 2796 12314 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12805 2839 12863 2845
rect 12805 2836 12817 2839
rect 12492 2808 12817 2836
rect 12492 2796 12498 2808
rect 12805 2805 12817 2808
rect 12851 2836 12863 2839
rect 12986 2836 12992 2848
rect 12851 2808 12992 2836
rect 12851 2805 12863 2808
rect 12805 2799 12863 2805
rect 12986 2796 12992 2808
rect 13044 2836 13050 2848
rect 13265 2839 13323 2845
rect 13265 2836 13277 2839
rect 13044 2808 13277 2836
rect 13044 2796 13050 2808
rect 13265 2805 13277 2808
rect 13311 2805 13323 2839
rect 14292 2836 14320 2932
rect 15105 2907 15163 2913
rect 15105 2873 15117 2907
rect 15151 2904 15163 2907
rect 15930 2904 15936 2916
rect 15151 2876 15936 2904
rect 15151 2873 15163 2876
rect 15105 2867 15163 2873
rect 15930 2864 15936 2876
rect 15988 2864 15994 2916
rect 15194 2836 15200 2848
rect 14292 2808 15200 2836
rect 13265 2799 13323 2805
rect 15194 2796 15200 2808
rect 15252 2836 15258 2848
rect 15565 2839 15623 2845
rect 15565 2836 15577 2839
rect 15252 2808 15577 2836
rect 15252 2796 15258 2808
rect 15565 2805 15577 2808
rect 15611 2805 15623 2839
rect 15565 2799 15623 2805
rect 1104 2746 16008 2768
rect 1104 2694 5979 2746
rect 6031 2694 6043 2746
rect 6095 2694 6107 2746
rect 6159 2694 6171 2746
rect 6223 2694 10976 2746
rect 11028 2694 11040 2746
rect 11092 2694 11104 2746
rect 11156 2694 11168 2746
rect 11220 2694 16008 2746
rect 1104 2672 16008 2694
rect 382 2592 388 2644
rect 440 2632 446 2644
rect 2133 2635 2191 2641
rect 2133 2632 2145 2635
rect 440 2604 2145 2632
rect 440 2592 446 2604
rect 2133 2601 2145 2604
rect 2179 2601 2191 2635
rect 2133 2595 2191 2601
rect 2501 2635 2559 2641
rect 2501 2601 2513 2635
rect 2547 2601 2559 2635
rect 2501 2595 2559 2601
rect 750 2524 756 2576
rect 808 2564 814 2576
rect 2516 2564 2544 2595
rect 3878 2592 3884 2644
rect 3936 2632 3942 2644
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 3936 2604 4077 2632
rect 3936 2592 3942 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 4522 2632 4528 2644
rect 4483 2604 4528 2632
rect 4065 2595 4123 2601
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 4614 2592 4620 2644
rect 4672 2632 4678 2644
rect 5813 2635 5871 2641
rect 5813 2632 5825 2635
rect 4672 2604 5825 2632
rect 4672 2592 4678 2604
rect 5813 2601 5825 2604
rect 5859 2601 5871 2635
rect 5813 2595 5871 2601
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6454 2632 6460 2644
rect 6411 2604 6460 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 6914 2632 6920 2644
rect 6875 2604 6920 2632
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2632 7435 2635
rect 7742 2632 7748 2644
rect 7423 2604 7748 2632
rect 7423 2601 7435 2604
rect 7377 2595 7435 2601
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 8202 2632 8208 2644
rect 8163 2604 8208 2632
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8570 2632 8576 2644
rect 8531 2604 8576 2632
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2632 9091 2635
rect 9582 2632 9588 2644
rect 9079 2604 9588 2632
rect 9079 2601 9091 2604
rect 9033 2595 9091 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 9950 2592 9956 2644
rect 10008 2632 10014 2644
rect 10045 2635 10103 2641
rect 10045 2632 10057 2635
rect 10008 2604 10057 2632
rect 10008 2592 10014 2604
rect 10045 2601 10057 2604
rect 10091 2601 10103 2635
rect 10045 2595 10103 2601
rect 10965 2635 11023 2641
rect 10965 2601 10977 2635
rect 11011 2632 11023 2635
rect 11330 2632 11336 2644
rect 11011 2604 11336 2632
rect 11011 2601 11023 2604
rect 10965 2595 11023 2601
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 11422 2592 11428 2644
rect 11480 2632 11486 2644
rect 12066 2632 12072 2644
rect 11480 2604 12072 2632
rect 11480 2592 11486 2604
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 12802 2632 12808 2644
rect 12763 2604 12808 2632
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 12894 2592 12900 2644
rect 12952 2632 12958 2644
rect 12989 2635 13047 2641
rect 12989 2632 13001 2635
rect 12952 2604 13001 2632
rect 12952 2592 12958 2604
rect 12989 2601 13001 2604
rect 13035 2601 13047 2635
rect 12989 2595 13047 2601
rect 14090 2592 14096 2644
rect 14148 2632 14154 2644
rect 14826 2632 14832 2644
rect 14148 2604 14832 2632
rect 14148 2592 14154 2604
rect 14826 2592 14832 2604
rect 14884 2632 14890 2644
rect 15473 2635 15531 2641
rect 15473 2632 15485 2635
rect 14884 2604 15485 2632
rect 14884 2592 14890 2604
rect 15473 2601 15485 2604
rect 15519 2601 15531 2635
rect 15473 2595 15531 2601
rect 808 2536 2544 2564
rect 808 2524 814 2536
rect 2590 2524 2596 2576
rect 2648 2564 2654 2576
rect 4430 2564 4436 2576
rect 2648 2536 3372 2564
rect 4391 2536 4436 2564
rect 2648 2524 2654 2536
rect 1489 2499 1547 2505
rect 1489 2465 1501 2499
rect 1535 2496 1547 2499
rect 1578 2496 1584 2508
rect 1535 2468 1584 2496
rect 1535 2465 1547 2468
rect 1489 2459 1547 2465
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 1946 2496 1952 2508
rect 1907 2468 1952 2496
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2314 2496 2320 2508
rect 2275 2468 2320 2496
rect 2314 2456 2320 2468
rect 2372 2456 2378 2508
rect 2682 2496 2688 2508
rect 2643 2468 2688 2496
rect 2682 2456 2688 2468
rect 2740 2456 2746 2508
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 3234 2496 3240 2508
rect 3191 2468 3240 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 3234 2456 3240 2468
rect 3292 2456 3298 2508
rect 3344 2496 3372 2536
rect 4430 2524 4436 2536
rect 4488 2524 4494 2576
rect 8113 2567 8171 2573
rect 4816 2536 5304 2564
rect 3513 2499 3571 2505
rect 3513 2496 3525 2499
rect 3344 2468 3525 2496
rect 3513 2465 3525 2468
rect 3559 2465 3571 2499
rect 3513 2459 3571 2465
rect 4338 2456 4344 2508
rect 4396 2496 4402 2508
rect 4816 2496 4844 2536
rect 4396 2468 4844 2496
rect 4893 2499 4951 2505
rect 4396 2456 4402 2468
rect 4893 2465 4905 2499
rect 4939 2496 4951 2499
rect 5166 2496 5172 2508
rect 4939 2468 5172 2496
rect 4939 2465 4951 2468
rect 4893 2459 4951 2465
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 5276 2505 5304 2536
rect 6012 2536 6960 2564
rect 5261 2499 5319 2505
rect 5261 2465 5273 2499
rect 5307 2465 5319 2499
rect 5626 2496 5632 2508
rect 5587 2468 5632 2496
rect 5261 2459 5319 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 6012 2505 6040 2536
rect 6932 2508 6960 2536
rect 8113 2533 8125 2567
rect 8159 2564 8171 2567
rect 9401 2567 9459 2573
rect 9401 2564 9413 2567
rect 8159 2536 9413 2564
rect 8159 2533 8171 2536
rect 8113 2527 8171 2533
rect 9401 2533 9413 2536
rect 9447 2533 9459 2567
rect 11974 2564 11980 2576
rect 9401 2527 9459 2533
rect 10244 2536 11980 2564
rect 5997 2499 6055 2505
rect 5997 2496 6009 2499
rect 5868 2468 6009 2496
rect 5868 2456 5874 2468
rect 5997 2465 6009 2468
rect 6043 2465 6055 2499
rect 6178 2496 6184 2508
rect 6139 2468 6184 2496
rect 5997 2459 6055 2465
rect 6178 2456 6184 2468
rect 6236 2456 6242 2508
rect 6914 2456 6920 2508
rect 6972 2456 6978 2508
rect 7285 2499 7343 2505
rect 7285 2465 7297 2499
rect 7331 2496 7343 2499
rect 8386 2496 8392 2508
rect 7331 2468 8392 2496
rect 7331 2465 7343 2468
rect 7285 2459 7343 2465
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 8941 2499 8999 2505
rect 8941 2465 8953 2499
rect 8987 2496 8999 2499
rect 9214 2496 9220 2508
rect 8987 2468 9220 2496
rect 8987 2465 8999 2468
rect 8941 2459 8999 2465
rect 9214 2456 9220 2468
rect 9272 2496 9278 2508
rect 9490 2496 9496 2508
rect 9272 2468 9496 2496
rect 9272 2456 9278 2468
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 9858 2496 9864 2508
rect 9819 2468 9864 2496
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 10244 2505 10272 2536
rect 11974 2524 11980 2536
rect 12032 2524 12038 2576
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2465 10287 2499
rect 10229 2459 10287 2465
rect 10597 2499 10655 2505
rect 10597 2465 10609 2499
rect 10643 2465 10655 2499
rect 10597 2459 10655 2465
rect 11333 2499 11391 2505
rect 11333 2465 11345 2499
rect 11379 2496 11391 2499
rect 11790 2496 11796 2508
rect 11379 2468 11796 2496
rect 11379 2465 11391 2468
rect 11333 2459 11391 2465
rect 2130 2388 2136 2440
rect 2188 2428 2194 2440
rect 4706 2428 4712 2440
rect 2188 2400 3740 2428
rect 4667 2400 4712 2428
rect 2188 2388 2194 2400
rect 106 2320 112 2372
rect 164 2360 170 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 164 2332 1777 2360
rect 164 2320 170 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 1854 2320 1860 2372
rect 1912 2360 1918 2372
rect 3712 2369 3740 2400
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 4798 2388 4804 2440
rect 4856 2428 4862 2440
rect 5718 2428 5724 2440
rect 4856 2400 5724 2428
rect 4856 2388 4862 2400
rect 5718 2388 5724 2400
rect 5776 2428 5782 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 5776 2400 6561 2428
rect 5776 2388 5782 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 2869 2363 2927 2369
rect 2869 2360 2881 2363
rect 1912 2332 2881 2360
rect 1912 2320 1918 2332
rect 2869 2329 2881 2332
rect 2915 2329 2927 2363
rect 2869 2323 2927 2329
rect 3697 2363 3755 2369
rect 3697 2329 3709 2363
rect 3743 2329 3755 2363
rect 3697 2323 3755 2329
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 5445 2363 5503 2369
rect 5445 2360 5457 2363
rect 4212 2332 5457 2360
rect 4212 2320 4218 2332
rect 5445 2329 5457 2332
rect 5491 2329 5503 2363
rect 7576 2360 7604 2391
rect 7834 2388 7840 2440
rect 7892 2428 7898 2440
rect 8297 2431 8355 2437
rect 8297 2428 8309 2431
rect 7892 2400 8309 2428
rect 7892 2388 7898 2400
rect 8297 2397 8309 2400
rect 8343 2428 8355 2431
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8343 2400 9137 2428
rect 8343 2397 8355 2400
rect 8297 2391 8355 2397
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 8846 2360 8852 2372
rect 7576 2332 8852 2360
rect 5445 2323 5503 2329
rect 8846 2320 8852 2332
rect 8904 2320 8910 2372
rect 10612 2360 10640 2459
rect 11790 2456 11796 2468
rect 11848 2496 11854 2508
rect 12161 2499 12219 2505
rect 12161 2496 12173 2499
rect 11848 2468 12173 2496
rect 11848 2456 11854 2468
rect 12161 2465 12173 2468
rect 12207 2465 12219 2499
rect 12161 2459 12219 2465
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 12912 2496 12940 2592
rect 14369 2567 14427 2573
rect 14369 2533 14381 2567
rect 14415 2564 14427 2567
rect 16574 2564 16580 2576
rect 14415 2536 16580 2564
rect 14415 2533 14427 2536
rect 14369 2527 14427 2533
rect 16574 2524 16580 2536
rect 16632 2524 16638 2576
rect 14090 2496 14096 2508
rect 12667 2468 12940 2496
rect 14051 2468 14096 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 14090 2456 14096 2468
rect 14148 2456 14154 2508
rect 14642 2496 14648 2508
rect 14603 2468 14648 2496
rect 14642 2456 14648 2468
rect 14700 2496 14706 2508
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 14700 2468 15209 2496
rect 14700 2456 14706 2468
rect 15197 2465 15209 2468
rect 15243 2465 15255 2499
rect 15197 2459 15255 2465
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 11425 2431 11483 2437
rect 11425 2428 11437 2431
rect 11296 2400 11437 2428
rect 11296 2388 11302 2400
rect 11425 2397 11437 2400
rect 11471 2397 11483 2431
rect 11606 2428 11612 2440
rect 11567 2400 11612 2428
rect 11425 2391 11483 2397
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 15562 2428 15568 2440
rect 14967 2400 15568 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 12434 2360 12440 2372
rect 10612 2332 12440 2360
rect 12434 2320 12440 2332
rect 12492 2320 12498 2372
rect 1118 2252 1124 2304
rect 1176 2292 1182 2304
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 1176 2264 3341 2292
rect 1176 2252 1182 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 3786 2252 3792 2304
rect 3844 2292 3850 2304
rect 5077 2295 5135 2301
rect 5077 2292 5089 2295
rect 3844 2264 5089 2292
rect 3844 2252 3850 2264
rect 5077 2261 5089 2264
rect 5123 2261 5135 2295
rect 5077 2255 5135 2261
rect 7745 2295 7803 2301
rect 7745 2261 7757 2295
rect 7791 2292 7803 2295
rect 8938 2292 8944 2304
rect 7791 2264 8944 2292
rect 7791 2261 7803 2264
rect 7745 2255 7803 2261
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 9122 2252 9128 2304
rect 9180 2292 9186 2304
rect 10413 2295 10471 2301
rect 10413 2292 10425 2295
rect 9180 2264 10425 2292
rect 9180 2252 9186 2264
rect 10413 2261 10425 2264
rect 10459 2261 10471 2295
rect 10778 2292 10784 2304
rect 10739 2264 10784 2292
rect 10413 2255 10471 2261
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 11238 2252 11244 2304
rect 11296 2292 11302 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11296 2264 11805 2292
rect 11296 2252 11302 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 11974 2252 11980 2304
rect 12032 2292 12038 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12032 2264 13185 2292
rect 12032 2252 12038 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 1104 2202 16008 2224
rect 1104 2150 3480 2202
rect 3532 2150 3544 2202
rect 3596 2150 3608 2202
rect 3660 2150 3672 2202
rect 3724 2150 8478 2202
rect 8530 2150 8542 2202
rect 8594 2150 8606 2202
rect 8658 2150 8670 2202
rect 8722 2150 13475 2202
rect 13527 2150 13539 2202
rect 13591 2150 13603 2202
rect 13655 2150 13667 2202
rect 13719 2150 16008 2202
rect 1104 2128 16008 2150
rect 3878 2048 3884 2100
rect 3936 2088 3942 2100
rect 9122 2088 9128 2100
rect 3936 2060 9128 2088
rect 3936 2048 3942 2060
rect 9122 2048 9128 2060
rect 9180 2048 9186 2100
rect 10686 2088 10692 2100
rect 9324 2060 10692 2088
rect 8018 1980 8024 2032
rect 8076 2020 8082 2032
rect 9324 2020 9352 2060
rect 10686 2048 10692 2060
rect 10744 2088 10750 2100
rect 11238 2088 11244 2100
rect 10744 2060 11244 2088
rect 10744 2048 10750 2060
rect 11238 2048 11244 2060
rect 11296 2048 11302 2100
rect 8076 1992 9352 2020
rect 8076 1980 8082 1992
rect 9490 1980 9496 2032
rect 9548 2020 9554 2032
rect 11698 2020 11704 2032
rect 9548 1992 11704 2020
rect 9548 1980 9554 1992
rect 11698 1980 11704 1992
rect 11756 1980 11762 2032
rect 2498 1912 2504 1964
rect 2556 1952 2562 1964
rect 10778 1952 10784 1964
rect 2556 1924 10784 1952
rect 2556 1912 2562 1924
rect 10778 1912 10784 1924
rect 10836 1912 10842 1964
rect 6178 1844 6184 1896
rect 6236 1884 6242 1896
rect 7558 1884 7564 1896
rect 6236 1856 7564 1884
rect 6236 1844 6242 1856
rect 7558 1844 7564 1856
rect 7616 1884 7622 1896
rect 11974 1884 11980 1896
rect 7616 1856 11980 1884
rect 7616 1844 7622 1856
rect 11974 1844 11980 1856
rect 12032 1844 12038 1896
rect 7098 1776 7104 1828
rect 7156 1816 7162 1828
rect 8662 1816 8668 1828
rect 7156 1788 8668 1816
rect 7156 1776 7162 1788
rect 8662 1776 8668 1788
rect 8720 1776 8726 1828
rect 10318 1776 10324 1828
rect 10376 1816 10382 1828
rect 12434 1816 12440 1828
rect 10376 1788 12440 1816
rect 10376 1776 10382 1788
rect 12434 1776 12440 1788
rect 12492 1776 12498 1828
rect 9306 1708 9312 1760
rect 9364 1748 9370 1760
rect 12158 1748 12164 1760
rect 9364 1720 12164 1748
rect 9364 1708 9370 1720
rect 12158 1708 12164 1720
rect 12216 1708 12222 1760
rect 5258 1504 5264 1556
rect 5316 1544 5322 1556
rect 7190 1544 7196 1556
rect 5316 1516 7196 1544
rect 5316 1504 5322 1516
rect 7190 1504 7196 1516
rect 7248 1504 7254 1556
<< via1 >>
rect 7564 17688 7616 17740
rect 15016 17688 15068 17740
rect 5264 17620 5316 17672
rect 6368 17620 6420 17672
rect 11980 17620 12032 17672
rect 1308 17552 1360 17604
rect 14648 17552 14700 17604
rect 6828 17484 6880 17536
rect 7748 17484 7800 17536
rect 10048 17484 10100 17536
rect 3480 17382 3532 17434
rect 3544 17382 3596 17434
rect 3608 17382 3660 17434
rect 3672 17382 3724 17434
rect 8478 17382 8530 17434
rect 8542 17382 8594 17434
rect 8606 17382 8658 17434
rect 8670 17382 8722 17434
rect 13475 17382 13527 17434
rect 13539 17382 13591 17434
rect 13603 17382 13655 17434
rect 13667 17382 13719 17434
rect 4620 17280 4672 17332
rect 5724 17280 5776 17332
rect 6368 17323 6420 17332
rect 6368 17289 6377 17323
rect 6377 17289 6411 17323
rect 6411 17289 6420 17323
rect 6368 17280 6420 17289
rect 6920 17280 6972 17332
rect 7288 17280 7340 17332
rect 7748 17323 7800 17332
rect 7748 17289 7757 17323
rect 7757 17289 7791 17323
rect 7791 17289 7800 17323
rect 7748 17280 7800 17289
rect 8300 17280 8352 17332
rect 8852 17280 8904 17332
rect 9128 17280 9180 17332
rect 940 17212 992 17264
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 2504 17212 2556 17264
rect 7564 17212 7616 17264
rect 8024 17212 8076 17264
rect 4436 17144 4488 17196
rect 7932 17144 7984 17196
rect 1584 17076 1636 17128
rect 1952 17076 2004 17128
rect 5264 17119 5316 17128
rect 2504 17008 2556 17060
rect 5264 17085 5273 17119
rect 5273 17085 5307 17119
rect 5307 17085 5316 17119
rect 5264 17076 5316 17085
rect 7472 17076 7524 17128
rect 8392 17076 8444 17128
rect 8484 17119 8536 17128
rect 8484 17085 8493 17119
rect 8493 17085 8527 17119
rect 8527 17085 8536 17119
rect 8484 17076 8536 17085
rect 8668 17076 8720 17128
rect 8944 17051 8996 17060
rect 8944 17017 8953 17051
rect 8953 17017 8987 17051
rect 8987 17017 8996 17051
rect 8944 17008 8996 17017
rect 3976 16940 4028 16992
rect 4988 16940 5040 16992
rect 5816 16940 5868 16992
rect 6276 16940 6328 16992
rect 6644 16983 6696 16992
rect 6644 16949 6653 16983
rect 6653 16949 6687 16983
rect 6687 16949 6696 16983
rect 6644 16940 6696 16949
rect 7748 16940 7800 16992
rect 9404 16940 9456 16992
rect 10324 16940 10376 16992
rect 14280 17076 14332 17128
rect 14832 17051 14884 17060
rect 14832 17017 14841 17051
rect 14841 17017 14875 17051
rect 14875 17017 14884 17051
rect 14832 17008 14884 17017
rect 11704 16940 11756 16992
rect 5979 16838 6031 16890
rect 6043 16838 6095 16890
rect 6107 16838 6159 16890
rect 6171 16838 6223 16890
rect 10976 16838 11028 16890
rect 11040 16838 11092 16890
rect 11104 16838 11156 16890
rect 11168 16838 11220 16890
rect 2504 16779 2556 16788
rect 2504 16745 2513 16779
rect 2513 16745 2547 16779
rect 2547 16745 2556 16779
rect 2504 16736 2556 16745
rect 2780 16736 2832 16788
rect 3792 16736 3844 16788
rect 4344 16736 4396 16788
rect 6552 16736 6604 16788
rect 7656 16736 7708 16788
rect 10140 16736 10192 16788
rect 2044 16668 2096 16720
rect 5540 16668 5592 16720
rect 3424 16643 3476 16652
rect 3424 16609 3433 16643
rect 3433 16609 3467 16643
rect 3467 16609 3476 16643
rect 3424 16600 3476 16609
rect 4436 16643 4488 16652
rect 3792 16575 3844 16584
rect 3792 16541 3801 16575
rect 3801 16541 3835 16575
rect 3835 16541 3844 16575
rect 3792 16532 3844 16541
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 4804 16643 4856 16652
rect 4804 16609 4813 16643
rect 4813 16609 4847 16643
rect 4847 16609 4856 16643
rect 4804 16600 4856 16609
rect 6000 16600 6052 16652
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 7564 16600 7616 16652
rect 5356 16575 5408 16584
rect 3148 16464 3200 16516
rect 3884 16464 3936 16516
rect 5356 16541 5365 16575
rect 5365 16541 5399 16575
rect 5399 16541 5408 16575
rect 5356 16532 5408 16541
rect 7748 16532 7800 16584
rect 6368 16464 6420 16516
rect 9680 16668 9732 16720
rect 8116 16600 8168 16652
rect 9496 16600 9548 16652
rect 9956 16643 10008 16652
rect 8944 16575 8996 16584
rect 8944 16541 8953 16575
rect 8953 16541 8987 16575
rect 8987 16541 8996 16575
rect 8944 16532 8996 16541
rect 9956 16609 9990 16643
rect 9990 16609 10008 16643
rect 9956 16600 10008 16609
rect 10232 16668 10284 16720
rect 11152 16668 11204 16720
rect 11612 16668 11664 16720
rect 12072 16600 12124 16652
rect 13268 16643 13320 16652
rect 13268 16609 13277 16643
rect 13277 16609 13311 16643
rect 13311 16609 13320 16643
rect 13268 16600 13320 16609
rect 14096 16600 14148 16652
rect 14648 16643 14700 16652
rect 14648 16609 14657 16643
rect 14657 16609 14691 16643
rect 14691 16609 14700 16643
rect 14648 16600 14700 16609
rect 9680 16575 9732 16584
rect 9680 16541 9689 16575
rect 9689 16541 9723 16575
rect 9723 16541 9732 16575
rect 11152 16575 11204 16584
rect 9680 16532 9732 16541
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 11428 16464 11480 16516
rect 12992 16464 13044 16516
rect 4988 16396 5040 16448
rect 6736 16439 6788 16448
rect 6736 16405 6745 16439
rect 6745 16405 6779 16439
rect 6779 16405 6788 16439
rect 6736 16396 6788 16405
rect 8300 16396 8352 16448
rect 3480 16294 3532 16346
rect 3544 16294 3596 16346
rect 3608 16294 3660 16346
rect 3672 16294 3724 16346
rect 8478 16294 8530 16346
rect 8542 16294 8594 16346
rect 8606 16294 8658 16346
rect 8670 16294 8722 16346
rect 13475 16294 13527 16346
rect 13539 16294 13591 16346
rect 13603 16294 13655 16346
rect 13667 16294 13719 16346
rect 1492 16192 1544 16244
rect 5632 16192 5684 16244
rect 6000 16235 6052 16244
rect 6000 16201 6009 16235
rect 6009 16201 6043 16235
rect 6043 16201 6052 16235
rect 6000 16192 6052 16201
rect 7748 16192 7800 16244
rect 8852 16192 8904 16244
rect 9956 16192 10008 16244
rect 10876 16192 10928 16244
rect 15108 16192 15160 16244
rect 204 16056 256 16108
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 10232 16124 10284 16176
rect 12256 16124 12308 16176
rect 2688 15988 2740 16040
rect 4620 16031 4672 16040
rect 4620 15997 4629 16031
rect 4629 15997 4663 16031
rect 4663 15997 4672 16031
rect 4620 15988 4672 15997
rect 5356 15988 5408 16040
rect 7748 16031 7800 16040
rect 7748 15997 7757 16031
rect 7757 15997 7791 16031
rect 7791 15997 7800 16031
rect 7748 15988 7800 15997
rect 10784 16056 10836 16108
rect 11612 16099 11664 16108
rect 11612 16065 11621 16099
rect 11621 16065 11655 16099
rect 11655 16065 11664 16099
rect 11612 16056 11664 16065
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 8300 15988 8352 16040
rect 9772 15988 9824 16040
rect 3332 15920 3384 15972
rect 9036 15920 9088 15972
rect 2320 15852 2372 15904
rect 4712 15852 4764 15904
rect 6460 15895 6512 15904
rect 6460 15861 6469 15895
rect 6469 15861 6503 15895
rect 6503 15861 6512 15895
rect 6460 15852 6512 15861
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 7288 15895 7340 15904
rect 7288 15861 7297 15895
rect 7297 15861 7331 15895
rect 7331 15861 7340 15895
rect 9956 15920 10008 15972
rect 7288 15852 7340 15861
rect 9588 15852 9640 15904
rect 10140 15852 10192 15904
rect 10508 15852 10560 15904
rect 11152 15988 11204 16040
rect 11888 15988 11940 16040
rect 13360 15988 13412 16040
rect 12624 15852 12676 15904
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 5979 15750 6031 15802
rect 6043 15750 6095 15802
rect 6107 15750 6159 15802
rect 6171 15750 6223 15802
rect 10976 15750 11028 15802
rect 11040 15750 11092 15802
rect 11104 15750 11156 15802
rect 11168 15750 11220 15802
rect 2412 15648 2464 15700
rect 1492 15555 1544 15564
rect 1492 15521 1501 15555
rect 1501 15521 1535 15555
rect 1535 15521 1544 15555
rect 1492 15512 1544 15521
rect 2964 15555 3016 15564
rect 2964 15521 2973 15555
rect 2973 15521 3007 15555
rect 3007 15521 3016 15555
rect 2964 15512 3016 15521
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 2872 15376 2924 15428
rect 4804 15580 4856 15632
rect 5264 15580 5316 15632
rect 6460 15648 6512 15700
rect 6552 15648 6604 15700
rect 6736 15623 6788 15632
rect 6736 15589 6748 15623
rect 6748 15589 6788 15623
rect 6736 15580 6788 15589
rect 7196 15580 7248 15632
rect 8208 15580 8260 15632
rect 8944 15648 8996 15700
rect 4988 15512 5040 15564
rect 5908 15512 5960 15564
rect 4344 15444 4396 15496
rect 4528 15487 4580 15496
rect 4528 15453 4537 15487
rect 4537 15453 4571 15487
rect 4571 15453 4580 15487
rect 4528 15444 4580 15453
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 7288 15512 7340 15564
rect 9220 15512 9272 15564
rect 9588 15580 9640 15632
rect 10416 15648 10468 15700
rect 10692 15648 10744 15700
rect 12808 15648 12860 15700
rect 10232 15580 10284 15632
rect 10600 15580 10652 15632
rect 11796 15580 11848 15632
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 11336 15555 11388 15564
rect 10048 15512 10100 15521
rect 4712 15444 4764 15453
rect 5356 15376 5408 15428
rect 5540 15376 5592 15428
rect 7748 15444 7800 15496
rect 9128 15487 9180 15496
rect 7932 15419 7984 15428
rect 4804 15308 4856 15360
rect 4988 15351 5040 15360
rect 4988 15317 4997 15351
rect 4997 15317 5031 15351
rect 5031 15317 5040 15351
rect 4988 15308 5040 15317
rect 5448 15351 5500 15360
rect 5448 15317 5457 15351
rect 5457 15317 5491 15351
rect 5491 15317 5500 15351
rect 5448 15308 5500 15317
rect 5908 15308 5960 15360
rect 6276 15351 6328 15360
rect 6276 15317 6285 15351
rect 6285 15317 6319 15351
rect 6319 15317 6328 15351
rect 6276 15308 6328 15317
rect 6368 15308 6420 15360
rect 7932 15385 7941 15419
rect 7941 15385 7975 15419
rect 7975 15385 7984 15419
rect 7932 15376 7984 15385
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9956 15444 10008 15496
rect 10140 15444 10192 15496
rect 11336 15521 11345 15555
rect 11345 15521 11379 15555
rect 11379 15521 11388 15555
rect 14372 15623 14424 15632
rect 14372 15589 14381 15623
rect 14381 15589 14415 15623
rect 14415 15589 14424 15623
rect 14372 15580 14424 15589
rect 11336 15512 11388 15521
rect 10968 15444 11020 15496
rect 9680 15376 9732 15428
rect 10048 15376 10100 15428
rect 10876 15376 10928 15428
rect 7840 15351 7892 15360
rect 7840 15317 7849 15351
rect 7849 15317 7883 15351
rect 7883 15317 7892 15351
rect 7840 15308 7892 15317
rect 8944 15308 8996 15360
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 11796 15444 11848 15496
rect 13176 15512 13228 15564
rect 12256 15487 12308 15496
rect 12256 15453 12265 15487
rect 12265 15453 12299 15487
rect 12299 15453 12308 15487
rect 12256 15444 12308 15453
rect 11428 15308 11480 15360
rect 14924 15308 14976 15360
rect 3480 15206 3532 15258
rect 3544 15206 3596 15258
rect 3608 15206 3660 15258
rect 3672 15206 3724 15258
rect 8478 15206 8530 15258
rect 8542 15206 8594 15258
rect 8606 15206 8658 15258
rect 8670 15206 8722 15258
rect 13475 15206 13527 15258
rect 13539 15206 13591 15258
rect 13603 15206 13655 15258
rect 13667 15206 13719 15258
rect 3332 15104 3384 15156
rect 4528 15104 4580 15156
rect 4804 15104 4856 15156
rect 9128 15104 9180 15156
rect 9496 15104 9548 15156
rect 4436 15036 4488 15088
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 9772 15036 9824 15088
rect 5540 15011 5592 15020
rect 5540 14977 5549 15011
rect 5549 14977 5583 15011
rect 5583 14977 5592 15011
rect 5540 14968 5592 14977
rect 6736 14968 6788 15020
rect 7380 15011 7432 15020
rect 5448 14900 5500 14952
rect 6828 14900 6880 14952
rect 7380 14977 7389 15011
rect 7389 14977 7423 15011
rect 7423 14977 7432 15011
rect 7380 14968 7432 14977
rect 7840 14968 7892 15020
rect 9036 15011 9088 15020
rect 9036 14977 9045 15011
rect 9045 14977 9079 15011
rect 9079 14977 9088 15011
rect 10232 15036 10284 15088
rect 9036 14968 9088 14977
rect 9956 14968 10008 15020
rect 10140 14900 10192 14952
rect 13176 15104 13228 15156
rect 16580 15104 16632 15156
rect 11336 15036 11388 15088
rect 12900 15036 12952 15088
rect 13084 15036 13136 15088
rect 11428 15011 11480 15020
rect 11428 14977 11437 15011
rect 11437 14977 11471 15011
rect 11471 14977 11480 15011
rect 11428 14968 11480 14977
rect 11612 15011 11664 15020
rect 11612 14977 11621 15011
rect 11621 14977 11655 15011
rect 11655 14977 11664 15011
rect 11612 14968 11664 14977
rect 12256 14968 12308 15020
rect 3240 14832 3292 14884
rect 4436 14832 4488 14884
rect 2688 14764 2740 14816
rect 3792 14764 3844 14816
rect 4252 14807 4304 14816
rect 4252 14773 4261 14807
rect 4261 14773 4295 14807
rect 4295 14773 4304 14807
rect 4252 14764 4304 14773
rect 5356 14764 5408 14816
rect 7012 14764 7064 14816
rect 7472 14764 7524 14816
rect 7932 14764 7984 14816
rect 8760 14764 8812 14816
rect 10692 14832 10744 14884
rect 12348 14832 12400 14884
rect 9680 14807 9732 14816
rect 9680 14773 9689 14807
rect 9689 14773 9723 14807
rect 9723 14773 9732 14807
rect 9680 14764 9732 14773
rect 10416 14764 10468 14816
rect 11796 14807 11848 14816
rect 11796 14773 11805 14807
rect 11805 14773 11839 14807
rect 11839 14773 11848 14807
rect 11796 14764 11848 14773
rect 12440 14807 12492 14816
rect 12440 14773 12449 14807
rect 12449 14773 12483 14807
rect 12483 14773 12492 14807
rect 12440 14764 12492 14773
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 12808 14764 12860 14773
rect 13544 14764 13596 14816
rect 5979 14662 6031 14714
rect 6043 14662 6095 14714
rect 6107 14662 6159 14714
rect 6171 14662 6223 14714
rect 10976 14662 11028 14714
rect 11040 14662 11092 14714
rect 11104 14662 11156 14714
rect 11168 14662 11220 14714
rect 2872 14424 2924 14476
rect 3056 14467 3108 14476
rect 3056 14433 3065 14467
rect 3065 14433 3099 14467
rect 3099 14433 3108 14467
rect 3056 14424 3108 14433
rect 5080 14467 5132 14476
rect 5080 14433 5089 14467
rect 5089 14433 5123 14467
rect 5123 14433 5132 14467
rect 5080 14424 5132 14433
rect 5724 14467 5776 14476
rect 5724 14433 5733 14467
rect 5733 14433 5767 14467
rect 5767 14433 5776 14467
rect 5724 14424 5776 14433
rect 5816 14424 5868 14476
rect 7012 14603 7064 14612
rect 7012 14569 7021 14603
rect 7021 14569 7055 14603
rect 7055 14569 7064 14603
rect 7012 14560 7064 14569
rect 7104 14560 7156 14612
rect 7840 14535 7892 14544
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 4068 14288 4120 14340
rect 4896 14356 4948 14408
rect 6644 14424 6696 14476
rect 7840 14501 7874 14535
rect 7874 14501 7892 14535
rect 7840 14492 7892 14501
rect 9036 14560 9088 14612
rect 8760 14492 8812 14544
rect 6920 14424 6972 14476
rect 7656 14424 7708 14476
rect 7104 14356 7156 14408
rect 9680 14560 9732 14612
rect 9772 14560 9824 14612
rect 11428 14560 11480 14612
rect 12348 14603 12400 14612
rect 12348 14569 12357 14603
rect 12357 14569 12391 14603
rect 12391 14569 12400 14603
rect 12348 14560 12400 14569
rect 12808 14560 12860 14612
rect 13544 14603 13596 14612
rect 13544 14569 13553 14603
rect 13553 14569 13587 14603
rect 13587 14569 13596 14603
rect 13544 14560 13596 14569
rect 10324 14424 10376 14476
rect 11612 14492 11664 14544
rect 11152 14424 11204 14476
rect 11888 14424 11940 14476
rect 12716 14467 12768 14476
rect 12716 14433 12725 14467
rect 12725 14433 12759 14467
rect 12759 14433 12768 14467
rect 12716 14424 12768 14433
rect 12900 14492 12952 14544
rect 16948 14492 17000 14544
rect 12992 14424 13044 14476
rect 10416 14288 10468 14340
rect 1584 14220 1636 14272
rect 4620 14220 4672 14272
rect 4988 14220 5040 14272
rect 5172 14263 5224 14272
rect 5172 14229 5181 14263
rect 5181 14229 5215 14263
rect 5215 14229 5224 14263
rect 5172 14220 5224 14229
rect 5264 14220 5316 14272
rect 7380 14220 7432 14272
rect 12072 14288 12124 14340
rect 12716 14288 12768 14340
rect 15476 14288 15528 14340
rect 12256 14220 12308 14272
rect 12808 14220 12860 14272
rect 13268 14220 13320 14272
rect 3480 14118 3532 14170
rect 3544 14118 3596 14170
rect 3608 14118 3660 14170
rect 3672 14118 3724 14170
rect 8478 14118 8530 14170
rect 8542 14118 8594 14170
rect 8606 14118 8658 14170
rect 8670 14118 8722 14170
rect 13475 14118 13527 14170
rect 13539 14118 13591 14170
rect 13603 14118 13655 14170
rect 13667 14118 13719 14170
rect 2964 14016 3016 14068
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 4712 14016 4764 14068
rect 2688 13923 2740 13932
rect 2688 13889 2697 13923
rect 2697 13889 2731 13923
rect 2731 13889 2740 13923
rect 2688 13880 2740 13889
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 4896 13880 4948 13932
rect 3976 13744 4028 13796
rect 5172 13812 5224 13864
rect 5264 13812 5316 13864
rect 4160 13719 4212 13728
rect 4160 13685 4169 13719
rect 4169 13685 4203 13719
rect 4203 13685 4212 13719
rect 4160 13676 4212 13685
rect 4620 13676 4672 13728
rect 5264 13719 5316 13728
rect 5264 13685 5273 13719
rect 5273 13685 5307 13719
rect 5307 13685 5316 13719
rect 5264 13676 5316 13685
rect 6368 13948 6420 14000
rect 5540 13880 5592 13932
rect 6644 13948 6696 14000
rect 8852 14016 8904 14068
rect 9772 14016 9824 14068
rect 10140 14059 10192 14068
rect 10140 14025 10149 14059
rect 10149 14025 10183 14059
rect 10183 14025 10192 14059
rect 10140 14016 10192 14025
rect 11152 14016 11204 14068
rect 6920 13923 6972 13932
rect 6920 13889 6929 13923
rect 6929 13889 6963 13923
rect 6963 13889 6972 13923
rect 6920 13880 6972 13889
rect 5724 13812 5776 13864
rect 6552 13812 6604 13864
rect 7472 13812 7524 13864
rect 8944 13880 8996 13932
rect 10784 13880 10836 13932
rect 11060 13948 11112 14000
rect 11612 13948 11664 14000
rect 8024 13812 8076 13864
rect 9864 13812 9916 13864
rect 10416 13812 10468 13864
rect 7380 13744 7432 13796
rect 8852 13787 8904 13796
rect 6736 13676 6788 13728
rect 7104 13676 7156 13728
rect 8852 13753 8861 13787
rect 8861 13753 8895 13787
rect 8895 13753 8904 13787
rect 8852 13744 8904 13753
rect 11060 13744 11112 13796
rect 11336 13812 11388 13864
rect 12256 14016 12308 14068
rect 12256 13880 12308 13932
rect 12072 13812 12124 13864
rect 16212 13744 16264 13796
rect 12624 13676 12676 13728
rect 13268 13676 13320 13728
rect 5979 13574 6031 13626
rect 6043 13574 6095 13626
rect 6107 13574 6159 13626
rect 6171 13574 6223 13626
rect 10976 13574 11028 13626
rect 11040 13574 11092 13626
rect 11104 13574 11156 13626
rect 11168 13574 11220 13626
rect 3240 13472 3292 13524
rect 4528 13472 4580 13524
rect 5264 13472 5316 13524
rect 6644 13472 6696 13524
rect 4068 13404 4120 13456
rect 5540 13404 5592 13456
rect 2596 13336 2648 13388
rect 5264 13336 5316 13388
rect 6920 13404 6972 13456
rect 9220 13472 9272 13524
rect 11428 13472 11480 13524
rect 11612 13515 11664 13524
rect 11612 13481 11621 13515
rect 11621 13481 11655 13515
rect 11655 13481 11664 13515
rect 11612 13472 11664 13481
rect 8208 13336 8260 13388
rect 4344 13268 4396 13320
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 4896 13268 4948 13277
rect 4988 13268 5040 13320
rect 4896 13132 4948 13184
rect 7380 13132 7432 13184
rect 8300 13132 8352 13184
rect 9496 13379 9548 13388
rect 9496 13345 9505 13379
rect 9505 13345 9539 13379
rect 9539 13345 9548 13379
rect 9496 13336 9548 13345
rect 11336 13336 11388 13388
rect 12440 13404 12492 13456
rect 15844 13336 15896 13388
rect 8852 13200 8904 13252
rect 9312 13268 9364 13320
rect 9404 13268 9456 13320
rect 10232 13268 10284 13320
rect 10784 13311 10836 13320
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 10876 13311 10928 13320
rect 10876 13277 10885 13311
rect 10885 13277 10919 13311
rect 10919 13277 10928 13311
rect 10876 13268 10928 13277
rect 13268 13268 13320 13320
rect 9404 13132 9456 13184
rect 10324 13175 10376 13184
rect 10324 13141 10333 13175
rect 10333 13141 10367 13175
rect 10367 13141 10376 13175
rect 10324 13132 10376 13141
rect 3480 13030 3532 13082
rect 3544 13030 3596 13082
rect 3608 13030 3660 13082
rect 3672 13030 3724 13082
rect 8478 13030 8530 13082
rect 8542 13030 8594 13082
rect 8606 13030 8658 13082
rect 8670 13030 8722 13082
rect 13475 13030 13527 13082
rect 13539 13030 13591 13082
rect 13603 13030 13655 13082
rect 13667 13030 13719 13082
rect 3056 12928 3108 12980
rect 5080 12928 5132 12980
rect 5264 12971 5316 12980
rect 5264 12937 5273 12971
rect 5273 12937 5307 12971
rect 5307 12937 5316 12971
rect 5264 12928 5316 12937
rect 4068 12792 4120 12844
rect 6644 12860 6696 12912
rect 4896 12792 4948 12844
rect 5540 12792 5592 12844
rect 6460 12792 6512 12844
rect 6920 12792 6972 12844
rect 4160 12724 4212 12776
rect 4344 12767 4396 12776
rect 4344 12733 4353 12767
rect 4353 12733 4387 12767
rect 4387 12733 4396 12767
rect 4344 12724 4396 12733
rect 10324 12928 10376 12980
rect 10784 12928 10836 12980
rect 9036 12860 9088 12912
rect 9312 12860 9364 12912
rect 7380 12835 7432 12844
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 4068 12656 4120 12708
rect 4620 12656 4672 12708
rect 5540 12588 5592 12640
rect 8300 12724 8352 12776
rect 7380 12656 7432 12708
rect 8760 12656 8812 12708
rect 6460 12588 6512 12640
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 11428 12835 11480 12844
rect 11428 12801 11437 12835
rect 11437 12801 11471 12835
rect 11471 12801 11480 12835
rect 11428 12792 11480 12801
rect 9128 12656 9180 12708
rect 9404 12724 9456 12776
rect 9680 12656 9732 12708
rect 9864 12656 9916 12708
rect 12440 12928 12492 12980
rect 13820 12928 13872 12980
rect 10876 12588 10928 12640
rect 11796 12631 11848 12640
rect 11796 12597 11805 12631
rect 11805 12597 11839 12631
rect 11839 12597 11848 12631
rect 11796 12588 11848 12597
rect 5979 12486 6031 12538
rect 6043 12486 6095 12538
rect 6107 12486 6159 12538
rect 6171 12486 6223 12538
rect 10976 12486 11028 12538
rect 11040 12486 11092 12538
rect 11104 12486 11156 12538
rect 11168 12486 11220 12538
rect 1768 12359 1820 12368
rect 1768 12325 1777 12359
rect 1777 12325 1811 12359
rect 1811 12325 1820 12359
rect 1768 12316 1820 12325
rect 5356 12384 5408 12436
rect 7380 12427 7432 12436
rect 6828 12316 6880 12368
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 8668 12384 8720 12436
rect 8760 12427 8812 12436
rect 8760 12393 8769 12427
rect 8769 12393 8803 12427
rect 8803 12393 8812 12427
rect 8760 12384 8812 12393
rect 9036 12384 9088 12436
rect 9404 12384 9456 12436
rect 11336 12427 11388 12436
rect 11336 12393 11345 12427
rect 11345 12393 11379 12427
rect 11379 12393 11388 12427
rect 11336 12384 11388 12393
rect 12716 12384 12768 12436
rect 8392 12359 8444 12368
rect 8392 12325 8401 12359
rect 8401 12325 8435 12359
rect 8435 12325 8444 12359
rect 8392 12316 8444 12325
rect 8944 12316 8996 12368
rect 9588 12316 9640 12368
rect 9864 12316 9916 12368
rect 6184 12291 6236 12300
rect 5172 12180 5224 12232
rect 1492 12044 1544 12096
rect 6184 12257 6218 12291
rect 6218 12257 6236 12291
rect 6184 12248 6236 12257
rect 6460 12248 6512 12300
rect 6736 12248 6788 12300
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 7564 12248 7616 12257
rect 5908 12223 5960 12232
rect 5908 12189 5917 12223
rect 5917 12189 5951 12223
rect 5951 12189 5960 12223
rect 5908 12180 5960 12189
rect 7012 12180 7064 12232
rect 8208 12248 8260 12300
rect 9956 12248 10008 12300
rect 10140 12291 10192 12300
rect 10140 12257 10174 12291
rect 10174 12257 10192 12291
rect 10140 12248 10192 12257
rect 5816 12112 5868 12164
rect 11612 12180 11664 12232
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 9036 12044 9088 12096
rect 9772 12044 9824 12096
rect 11428 12112 11480 12164
rect 10140 12044 10192 12096
rect 11704 12044 11756 12096
rect 12716 12044 12768 12096
rect 3480 11942 3532 11994
rect 3544 11942 3596 11994
rect 3608 11942 3660 11994
rect 3672 11942 3724 11994
rect 8478 11942 8530 11994
rect 8542 11942 8594 11994
rect 8606 11942 8658 11994
rect 8670 11942 8722 11994
rect 13475 11942 13527 11994
rect 13539 11942 13591 11994
rect 13603 11942 13655 11994
rect 13667 11942 13719 11994
rect 6736 11840 6788 11892
rect 7104 11840 7156 11892
rect 8208 11772 8260 11824
rect 8852 11840 8904 11892
rect 9772 11840 9824 11892
rect 10508 11840 10560 11892
rect 10600 11772 10652 11824
rect 10140 11704 10192 11756
rect 1492 11679 1544 11688
rect 1492 11645 1501 11679
rect 1501 11645 1535 11679
rect 1535 11645 1544 11679
rect 1492 11636 1544 11645
rect 2044 11679 2096 11688
rect 2044 11645 2053 11679
rect 2053 11645 2087 11679
rect 2087 11645 2096 11679
rect 2044 11636 2096 11645
rect 2412 11636 2464 11688
rect 4804 11636 4856 11688
rect 5908 11636 5960 11688
rect 7104 11636 7156 11688
rect 7288 11636 7340 11688
rect 8944 11636 8996 11688
rect 9496 11636 9548 11688
rect 1768 11611 1820 11620
rect 1768 11577 1777 11611
rect 1777 11577 1811 11611
rect 1811 11577 1820 11611
rect 1768 11568 1820 11577
rect 2780 11568 2832 11620
rect 3792 11568 3844 11620
rect 4988 11611 5040 11620
rect 3148 11543 3200 11552
rect 3148 11509 3157 11543
rect 3157 11509 3191 11543
rect 3191 11509 3200 11543
rect 3148 11500 3200 11509
rect 4988 11577 5022 11611
rect 5022 11577 5040 11611
rect 4988 11568 5040 11577
rect 4896 11500 4948 11552
rect 7012 11568 7064 11620
rect 8300 11568 8352 11620
rect 6276 11500 6328 11552
rect 6736 11500 6788 11552
rect 7656 11500 7708 11552
rect 9128 11568 9180 11620
rect 9772 11568 9824 11620
rect 10324 11704 10376 11756
rect 5979 11398 6031 11450
rect 6043 11398 6095 11450
rect 6107 11398 6159 11450
rect 6171 11398 6223 11450
rect 10976 11398 11028 11450
rect 11040 11398 11092 11450
rect 11104 11398 11156 11450
rect 11168 11398 11220 11450
rect 2044 11296 2096 11348
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 4620 11296 4672 11348
rect 5632 11296 5684 11348
rect 5724 11296 5776 11348
rect 7656 11339 7708 11348
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 1584 11092 1636 11144
rect 2964 11160 3016 11212
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 4436 11024 4488 11076
rect 6460 11228 6512 11280
rect 7656 11305 7665 11339
rect 7665 11305 7699 11339
rect 7699 11305 7708 11339
rect 7656 11296 7708 11305
rect 9864 11296 9916 11348
rect 7840 11228 7892 11280
rect 8116 11228 8168 11280
rect 8300 11271 8352 11280
rect 8300 11237 8309 11271
rect 8309 11237 8343 11271
rect 8343 11237 8352 11271
rect 8300 11228 8352 11237
rect 5080 11203 5132 11212
rect 5080 11169 5089 11203
rect 5089 11169 5123 11203
rect 5123 11169 5132 11203
rect 5080 11160 5132 11169
rect 5540 11160 5592 11212
rect 5908 11203 5960 11212
rect 5908 11169 5917 11203
rect 5917 11169 5951 11203
rect 5951 11169 5960 11203
rect 5908 11160 5960 11169
rect 4988 11092 5040 11144
rect 6736 11092 6788 11144
rect 9220 11228 9272 11280
rect 4804 11024 4856 11076
rect 5540 11024 5592 11076
rect 7196 11024 7248 11076
rect 8944 11092 8996 11144
rect 9128 11092 9180 11144
rect 10048 11160 10100 11212
rect 12992 11160 13044 11212
rect 9956 11092 10008 11144
rect 10140 11092 10192 11144
rect 10784 11092 10836 11144
rect 11060 11024 11112 11076
rect 7288 10999 7340 11008
rect 7288 10965 7297 10999
rect 7297 10965 7331 10999
rect 7331 10965 7340 10999
rect 7288 10956 7340 10965
rect 8300 10956 8352 11008
rect 9036 10956 9088 11008
rect 9220 10999 9272 11008
rect 9220 10965 9229 10999
rect 9229 10965 9263 10999
rect 9263 10965 9272 10999
rect 9220 10956 9272 10965
rect 12716 10999 12768 11008
rect 12716 10965 12725 10999
rect 12725 10965 12759 10999
rect 12759 10965 12768 10999
rect 12716 10956 12768 10965
rect 3480 10854 3532 10906
rect 3544 10854 3596 10906
rect 3608 10854 3660 10906
rect 3672 10854 3724 10906
rect 8478 10854 8530 10906
rect 8542 10854 8594 10906
rect 8606 10854 8658 10906
rect 8670 10854 8722 10906
rect 13475 10854 13527 10906
rect 13539 10854 13591 10906
rect 13603 10854 13655 10906
rect 13667 10854 13719 10906
rect 1860 10752 1912 10804
rect 4620 10752 4672 10804
rect 5172 10795 5224 10804
rect 5172 10761 5181 10795
rect 5181 10761 5215 10795
rect 5215 10761 5224 10795
rect 5172 10752 5224 10761
rect 5816 10752 5868 10804
rect 7104 10752 7156 10804
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 3148 10684 3200 10736
rect 5724 10684 5776 10736
rect 3700 10659 3752 10668
rect 2596 10548 2648 10600
rect 3700 10625 3709 10659
rect 3709 10625 3743 10659
rect 3743 10625 3752 10659
rect 3700 10616 3752 10625
rect 4436 10659 4488 10668
rect 4436 10625 4445 10659
rect 4445 10625 4479 10659
rect 4479 10625 4488 10659
rect 4436 10616 4488 10625
rect 4988 10616 5040 10668
rect 5172 10616 5224 10668
rect 6276 10616 6328 10668
rect 8208 10659 8260 10668
rect 8208 10625 8217 10659
rect 8217 10625 8251 10659
rect 8251 10625 8260 10659
rect 8208 10616 8260 10625
rect 5356 10548 5408 10600
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 5908 10548 5960 10600
rect 6736 10548 6788 10600
rect 7288 10548 7340 10600
rect 8300 10548 8352 10600
rect 9864 10752 9916 10804
rect 11336 10727 11388 10736
rect 11336 10693 11345 10727
rect 11345 10693 11379 10727
rect 11379 10693 11388 10727
rect 11336 10684 11388 10693
rect 9864 10616 9916 10668
rect 11060 10616 11112 10668
rect 12716 10616 12768 10668
rect 9036 10548 9088 10600
rect 10784 10548 10836 10600
rect 2228 10412 2280 10464
rect 3332 10480 3384 10532
rect 4252 10480 4304 10532
rect 4620 10480 4672 10532
rect 3056 10412 3108 10464
rect 6920 10480 6972 10532
rect 6460 10412 6512 10464
rect 6736 10412 6788 10464
rect 7196 10412 7248 10464
rect 7380 10412 7432 10464
rect 8300 10412 8352 10464
rect 9128 10480 9180 10532
rect 8852 10412 8904 10464
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 11428 10455 11480 10464
rect 11428 10421 11437 10455
rect 11437 10421 11471 10455
rect 11471 10421 11480 10455
rect 11428 10412 11480 10421
rect 12624 10480 12676 10532
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 13360 10412 13412 10464
rect 5979 10310 6031 10362
rect 6043 10310 6095 10362
rect 6107 10310 6159 10362
rect 6171 10310 6223 10362
rect 10976 10310 11028 10362
rect 11040 10310 11092 10362
rect 11104 10310 11156 10362
rect 11168 10310 11220 10362
rect 2964 10251 3016 10260
rect 2964 10217 2973 10251
rect 2973 10217 3007 10251
rect 3007 10217 3016 10251
rect 2964 10208 3016 10217
rect 4528 10208 4580 10260
rect 6920 10208 6972 10260
rect 7656 10208 7708 10260
rect 8760 10208 8812 10260
rect 12624 10208 12676 10260
rect 12808 10208 12860 10260
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 16212 10208 16264 10260
rect 2412 10140 2464 10192
rect 3884 10140 3936 10192
rect 2136 10072 2188 10124
rect 4344 10072 4396 10124
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 3792 10004 3844 10013
rect 2964 9868 3016 9920
rect 4804 10072 4856 10124
rect 5540 10140 5592 10192
rect 6736 10140 6788 10192
rect 9404 10140 9456 10192
rect 11336 10140 11388 10192
rect 11980 10140 12032 10192
rect 12440 10140 12492 10192
rect 7196 10072 7248 10124
rect 9496 10072 9548 10124
rect 9956 10072 10008 10124
rect 7472 10004 7524 10056
rect 6920 9936 6972 9988
rect 8116 9936 8168 9988
rect 8760 9936 8812 9988
rect 9956 9936 10008 9988
rect 12992 10004 13044 10056
rect 12808 9936 12860 9988
rect 5080 9911 5132 9920
rect 5080 9877 5089 9911
rect 5089 9877 5123 9911
rect 5123 9877 5132 9911
rect 5080 9868 5132 9877
rect 5356 9868 5408 9920
rect 7012 9868 7064 9920
rect 7564 9868 7616 9920
rect 9128 9868 9180 9920
rect 3480 9766 3532 9818
rect 3544 9766 3596 9818
rect 3608 9766 3660 9818
rect 3672 9766 3724 9818
rect 8478 9766 8530 9818
rect 8542 9766 8594 9818
rect 8606 9766 8658 9818
rect 8670 9766 8722 9818
rect 13475 9766 13527 9818
rect 13539 9766 13591 9818
rect 13603 9766 13655 9818
rect 13667 9766 13719 9818
rect 3792 9596 3844 9648
rect 6552 9596 6604 9648
rect 8116 9664 8168 9716
rect 9772 9664 9824 9716
rect 11612 9664 11664 9716
rect 3700 9571 3752 9580
rect 3700 9537 3709 9571
rect 3709 9537 3743 9571
rect 3743 9537 3752 9571
rect 3700 9528 3752 9537
rect 8300 9596 8352 9648
rect 8760 9596 8812 9648
rect 9220 9596 9272 9648
rect 10048 9639 10100 9648
rect 10048 9605 10057 9639
rect 10057 9605 10091 9639
rect 10091 9605 10100 9639
rect 10048 9596 10100 9605
rect 1492 9503 1544 9512
rect 1492 9469 1501 9503
rect 1501 9469 1535 9503
rect 1535 9469 1544 9503
rect 1492 9460 1544 9469
rect 2044 9503 2096 9512
rect 2044 9469 2053 9503
rect 2053 9469 2087 9503
rect 2087 9469 2096 9503
rect 2044 9460 2096 9469
rect 3148 9460 3200 9512
rect 4252 9460 4304 9512
rect 4804 9460 4856 9512
rect 1768 9435 1820 9444
rect 1768 9401 1777 9435
rect 1777 9401 1811 9435
rect 1811 9401 1820 9435
rect 1768 9392 1820 9401
rect 2596 9392 2648 9444
rect 4988 9460 5040 9512
rect 5356 9503 5408 9512
rect 5356 9469 5390 9503
rect 5390 9469 5408 9503
rect 5356 9460 5408 9469
rect 5632 9460 5684 9512
rect 7104 9435 7156 9444
rect 7104 9401 7138 9435
rect 7138 9401 7156 9435
rect 7104 9392 7156 9401
rect 2136 9324 2188 9376
rect 4252 9367 4304 9376
rect 4252 9333 4261 9367
rect 4261 9333 4295 9367
rect 4295 9333 4304 9367
rect 4252 9324 4304 9333
rect 4620 9367 4672 9376
rect 4620 9333 4629 9367
rect 4629 9333 4663 9367
rect 4663 9333 4672 9367
rect 4620 9324 4672 9333
rect 6368 9324 6420 9376
rect 7656 9324 7708 9376
rect 8116 9324 8168 9376
rect 8852 9528 8904 9580
rect 9128 9571 9180 9580
rect 9128 9537 9137 9571
rect 9137 9537 9171 9571
rect 9171 9537 9180 9571
rect 9128 9528 9180 9537
rect 10324 9528 10376 9580
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 12716 9528 12768 9580
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 9220 9460 9272 9512
rect 9496 9460 9548 9512
rect 8392 9435 8444 9444
rect 8392 9401 8401 9435
rect 8401 9401 8435 9435
rect 8435 9401 8444 9435
rect 8392 9392 8444 9401
rect 9680 9392 9732 9444
rect 9404 9324 9456 9376
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 11612 9460 11664 9512
rect 12072 9460 12124 9512
rect 13084 9460 13136 9512
rect 15016 9503 15068 9512
rect 11336 9435 11388 9444
rect 11336 9401 11345 9435
rect 11345 9401 11379 9435
rect 11379 9401 11388 9435
rect 11336 9392 11388 9401
rect 11428 9392 11480 9444
rect 10048 9324 10100 9376
rect 10232 9324 10284 9376
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 13820 9324 13872 9376
rect 15016 9469 15025 9503
rect 15025 9469 15059 9503
rect 15059 9469 15068 9503
rect 15016 9460 15068 9469
rect 5979 9222 6031 9274
rect 6043 9222 6095 9274
rect 6107 9222 6159 9274
rect 6171 9222 6223 9274
rect 10976 9222 11028 9274
rect 11040 9222 11092 9274
rect 11104 9222 11156 9274
rect 11168 9222 11220 9274
rect 1584 9120 1636 9172
rect 2228 9120 2280 9172
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 4252 9120 4304 9172
rect 4344 9120 4396 9172
rect 8392 9120 8444 9172
rect 10140 9120 10192 9172
rect 10324 9120 10376 9172
rect 2872 9052 2924 9104
rect 3332 9052 3384 9104
rect 6736 9052 6788 9104
rect 7380 9052 7432 9104
rect 2688 9027 2740 9036
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 2688 8984 2740 8993
rect 2780 9027 2832 9036
rect 2780 8993 2789 9027
rect 2789 8993 2823 9027
rect 2823 8993 2832 9027
rect 2780 8984 2832 8993
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 2596 8916 2648 8968
rect 5448 8984 5500 9036
rect 5540 8984 5592 9036
rect 6368 8984 6420 9036
rect 9496 9052 9548 9104
rect 9772 9052 9824 9104
rect 12256 9120 12308 9172
rect 12532 9120 12584 9172
rect 12900 9120 12952 9172
rect 12992 9120 13044 9172
rect 10692 9052 10744 9104
rect 3056 8848 3108 8900
rect 5724 8916 5776 8968
rect 5816 8916 5868 8968
rect 6184 8959 6236 8968
rect 6184 8925 6193 8959
rect 6193 8925 6227 8959
rect 6227 8925 6236 8959
rect 6184 8916 6236 8925
rect 7104 8959 7156 8968
rect 7104 8925 7113 8959
rect 7113 8925 7147 8959
rect 7147 8925 7156 8959
rect 7748 8959 7800 8968
rect 7104 8916 7156 8925
rect 2688 8780 2740 8832
rect 4252 8780 4304 8832
rect 4528 8823 4580 8832
rect 4528 8789 4537 8823
rect 4537 8789 4571 8823
rect 4571 8789 4580 8823
rect 4528 8780 4580 8789
rect 4620 8780 4672 8832
rect 6552 8780 6604 8832
rect 7748 8925 7757 8959
rect 7757 8925 7791 8959
rect 7791 8925 7800 8959
rect 7748 8916 7800 8925
rect 8208 8984 8260 9036
rect 9864 8984 9916 9036
rect 10140 8984 10192 9036
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 10416 8916 10468 8968
rect 10692 8959 10744 8968
rect 10692 8925 10701 8959
rect 10701 8925 10735 8959
rect 10735 8925 10744 8959
rect 10692 8916 10744 8925
rect 11244 8984 11296 9036
rect 12716 8984 12768 9036
rect 11336 8848 11388 8900
rect 10140 8780 10192 8832
rect 12992 8780 13044 8832
rect 3480 8678 3532 8730
rect 3544 8678 3596 8730
rect 3608 8678 3660 8730
rect 3672 8678 3724 8730
rect 8478 8678 8530 8730
rect 8542 8678 8594 8730
rect 8606 8678 8658 8730
rect 8670 8678 8722 8730
rect 13475 8678 13527 8730
rect 13539 8678 13591 8730
rect 13603 8678 13655 8730
rect 13667 8678 13719 8730
rect 7196 8576 7248 8628
rect 7748 8576 7800 8628
rect 9496 8619 9548 8628
rect 9496 8585 9505 8619
rect 9505 8585 9539 8619
rect 9539 8585 9548 8619
rect 9496 8576 9548 8585
rect 9956 8576 10008 8628
rect 4896 8508 4948 8560
rect 6184 8508 6236 8560
rect 6920 8508 6972 8560
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 2044 8372 2096 8424
rect 3332 8347 3384 8356
rect 3332 8313 3366 8347
rect 3366 8313 3384 8347
rect 3332 8304 3384 8313
rect 3056 8236 3108 8288
rect 4988 8440 5040 8492
rect 6276 8440 6328 8492
rect 6644 8440 6696 8492
rect 8484 8508 8536 8560
rect 9772 8508 9824 8560
rect 10508 8576 10560 8628
rect 12164 8576 12216 8628
rect 11244 8508 11296 8560
rect 12348 8508 12400 8560
rect 4528 8372 4580 8424
rect 6368 8372 6420 8424
rect 8300 8440 8352 8492
rect 8116 8372 8168 8424
rect 9128 8440 9180 8492
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 11428 8483 11480 8492
rect 11428 8449 11437 8483
rect 11437 8449 11471 8483
rect 11471 8449 11480 8483
rect 11428 8440 11480 8449
rect 12716 8440 12768 8492
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 8668 8372 8720 8424
rect 10324 8372 10376 8424
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 9312 8304 9364 8356
rect 10600 8304 10652 8356
rect 11796 8372 11848 8424
rect 12072 8415 12124 8424
rect 12072 8381 12081 8415
rect 12081 8381 12115 8415
rect 12115 8381 12124 8415
rect 12808 8415 12860 8424
rect 12072 8372 12124 8381
rect 12808 8381 12817 8415
rect 12817 8381 12851 8415
rect 12851 8381 12860 8415
rect 12808 8372 12860 8381
rect 13912 8372 13964 8424
rect 6644 8279 6696 8288
rect 6644 8245 6653 8279
rect 6653 8245 6687 8279
rect 6687 8245 6696 8279
rect 6644 8236 6696 8245
rect 7472 8236 7524 8288
rect 7564 8236 7616 8288
rect 7748 8236 7800 8288
rect 8392 8236 8444 8288
rect 9956 8236 10008 8288
rect 10324 8236 10376 8288
rect 10416 8236 10468 8288
rect 12440 8236 12492 8288
rect 12808 8236 12860 8288
rect 13176 8304 13228 8356
rect 13360 8347 13412 8356
rect 13360 8313 13369 8347
rect 13369 8313 13403 8347
rect 13403 8313 13412 8347
rect 13360 8304 13412 8313
rect 5979 8134 6031 8186
rect 6043 8134 6095 8186
rect 6107 8134 6159 8186
rect 6171 8134 6223 8186
rect 10976 8134 11028 8186
rect 11040 8134 11092 8186
rect 11104 8134 11156 8186
rect 11168 8134 11220 8186
rect 1584 8032 1636 8084
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 5724 8032 5776 8084
rect 7932 8032 7984 8084
rect 8484 8075 8536 8084
rect 2044 7896 2096 7948
rect 3240 7896 3292 7948
rect 4712 7896 4764 7948
rect 4804 7896 4856 7948
rect 5908 7939 5960 7948
rect 5908 7905 5917 7939
rect 5917 7905 5951 7939
rect 5951 7905 5960 7939
rect 5908 7896 5960 7905
rect 3884 7828 3936 7880
rect 3332 7803 3384 7812
rect 3332 7769 3341 7803
rect 3341 7769 3375 7803
rect 3375 7769 3384 7803
rect 5080 7828 5132 7880
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 6092 7828 6144 7880
rect 6368 7828 6420 7880
rect 3332 7760 3384 7769
rect 2872 7692 2924 7744
rect 4620 7692 4672 7744
rect 6368 7735 6420 7744
rect 6368 7701 6377 7735
rect 6377 7701 6411 7735
rect 6411 7701 6420 7735
rect 6368 7692 6420 7701
rect 6736 7964 6788 8016
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 9312 8032 9364 8084
rect 9588 8032 9640 8084
rect 9956 8075 10008 8084
rect 9956 8041 9965 8075
rect 9965 8041 9999 8075
rect 9999 8041 10008 8075
rect 9956 8032 10008 8041
rect 10784 8032 10836 8084
rect 11336 8032 11388 8084
rect 11428 8032 11480 8084
rect 12164 8032 12216 8084
rect 12716 8032 12768 8084
rect 8300 7964 8352 8016
rect 8760 7964 8812 8016
rect 9128 7964 9180 8016
rect 9772 7964 9824 8016
rect 6552 7939 6604 7948
rect 6552 7905 6561 7939
rect 6561 7905 6595 7939
rect 6595 7905 6604 7939
rect 6920 7939 6972 7948
rect 6552 7896 6604 7905
rect 6920 7905 6954 7939
rect 6954 7905 6972 7939
rect 6920 7896 6972 7905
rect 8944 7896 8996 7948
rect 10692 7939 10744 7948
rect 10692 7905 10701 7939
rect 10701 7905 10735 7939
rect 10735 7905 10744 7939
rect 10692 7896 10744 7905
rect 11336 7896 11388 7948
rect 6552 7760 6604 7812
rect 9404 7828 9456 7880
rect 10600 7828 10652 7880
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 10140 7760 10192 7812
rect 7656 7692 7708 7744
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 3480 7590 3532 7642
rect 3544 7590 3596 7642
rect 3608 7590 3660 7642
rect 3672 7590 3724 7642
rect 8478 7590 8530 7642
rect 8542 7590 8594 7642
rect 8606 7590 8658 7642
rect 8670 7590 8722 7642
rect 13475 7590 13527 7642
rect 13539 7590 13591 7642
rect 13603 7590 13655 7642
rect 13667 7590 13719 7642
rect 3884 7531 3936 7540
rect 3884 7497 3893 7531
rect 3893 7497 3927 7531
rect 3927 7497 3936 7531
rect 3884 7488 3936 7497
rect 4712 7531 4764 7540
rect 4712 7497 4721 7531
rect 4721 7497 4755 7531
rect 4755 7497 4764 7531
rect 4712 7488 4764 7497
rect 5816 7531 5868 7540
rect 5816 7497 5825 7531
rect 5825 7497 5859 7531
rect 5859 7497 5868 7531
rect 5816 7488 5868 7497
rect 6552 7488 6604 7540
rect 10324 7488 10376 7540
rect 10692 7488 10744 7540
rect 10140 7420 10192 7472
rect 14832 7420 14884 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 3148 7284 3200 7336
rect 3240 7284 3292 7336
rect 3792 7284 3844 7336
rect 5080 7327 5132 7336
rect 4068 7216 4120 7268
rect 4620 7216 4672 7268
rect 5080 7293 5089 7327
rect 5089 7293 5123 7327
rect 5123 7293 5132 7327
rect 5080 7284 5132 7293
rect 5172 7327 5224 7336
rect 5172 7293 5181 7327
rect 5181 7293 5215 7327
rect 5215 7293 5224 7327
rect 5816 7352 5868 7404
rect 6460 7395 6512 7404
rect 6460 7361 6469 7395
rect 6469 7361 6503 7395
rect 6503 7361 6512 7395
rect 6460 7352 6512 7361
rect 6920 7352 6972 7404
rect 7012 7352 7064 7404
rect 5172 7284 5224 7293
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 5908 7284 5960 7336
rect 7104 7284 7156 7336
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 6552 7216 6604 7268
rect 6644 7216 6696 7268
rect 7380 7216 7432 7268
rect 2688 7191 2740 7200
rect 2688 7157 2697 7191
rect 2697 7157 2731 7191
rect 2731 7157 2740 7191
rect 2688 7148 2740 7157
rect 3148 7191 3200 7200
rect 3148 7157 3157 7191
rect 3157 7157 3191 7191
rect 3191 7157 3200 7191
rect 4252 7191 4304 7200
rect 3148 7148 3200 7157
rect 4252 7157 4261 7191
rect 4261 7157 4295 7191
rect 4295 7157 4304 7191
rect 4252 7148 4304 7157
rect 5632 7148 5684 7200
rect 7748 7284 7800 7336
rect 7932 7327 7984 7336
rect 7932 7293 7966 7327
rect 7966 7293 7984 7327
rect 7932 7284 7984 7293
rect 9772 7284 9824 7336
rect 7748 7148 7800 7200
rect 9312 7216 9364 7268
rect 9864 7148 9916 7200
rect 11336 7352 11388 7404
rect 10600 7284 10652 7336
rect 11428 7284 11480 7336
rect 11888 7284 11940 7336
rect 12072 7284 12124 7336
rect 10692 7216 10744 7268
rect 10876 7216 10928 7268
rect 12440 7216 12492 7268
rect 10600 7191 10652 7200
rect 10600 7157 10609 7191
rect 10609 7157 10643 7191
rect 10643 7157 10652 7191
rect 11888 7191 11940 7200
rect 10600 7148 10652 7157
rect 11888 7157 11897 7191
rect 11897 7157 11931 7191
rect 11931 7157 11940 7191
rect 11888 7148 11940 7157
rect 5979 7046 6031 7098
rect 6043 7046 6095 7098
rect 6107 7046 6159 7098
rect 6171 7046 6223 7098
rect 10976 7046 11028 7098
rect 11040 7046 11092 7098
rect 11104 7046 11156 7098
rect 11168 7046 11220 7098
rect 2688 6944 2740 6996
rect 3148 6944 3200 6996
rect 3792 6987 3844 6996
rect 3792 6953 3801 6987
rect 3801 6953 3835 6987
rect 3835 6953 3844 6987
rect 3792 6944 3844 6953
rect 4068 6987 4120 6996
rect 4068 6953 4077 6987
rect 4077 6953 4111 6987
rect 4111 6953 4120 6987
rect 4068 6944 4120 6953
rect 5448 6987 5500 6996
rect 5448 6953 5457 6987
rect 5457 6953 5491 6987
rect 5491 6953 5500 6987
rect 5448 6944 5500 6953
rect 6552 6987 6604 6996
rect 6552 6953 6561 6987
rect 6561 6953 6595 6987
rect 6595 6953 6604 6987
rect 6552 6944 6604 6953
rect 6920 6944 6972 6996
rect 8116 6987 8168 6996
rect 8116 6953 8125 6987
rect 8125 6953 8159 6987
rect 8159 6953 8168 6987
rect 8116 6944 8168 6953
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 11428 6987 11480 6996
rect 11428 6953 11437 6987
rect 11437 6953 11471 6987
rect 11471 6953 11480 6987
rect 11428 6944 11480 6953
rect 11888 6944 11940 6996
rect 12440 6987 12492 6996
rect 12440 6953 12449 6987
rect 12449 6953 12483 6987
rect 12483 6953 12492 6987
rect 12440 6944 12492 6953
rect 2872 6876 2924 6928
rect 3240 6876 3292 6928
rect 3332 6808 3384 6860
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 4988 6876 5040 6928
rect 4068 6740 4120 6792
rect 6368 6876 6420 6928
rect 5908 6851 5960 6860
rect 5908 6817 5917 6851
rect 5917 6817 5951 6851
rect 5951 6817 5960 6851
rect 5908 6808 5960 6817
rect 6828 6808 6880 6860
rect 7012 6851 7064 6860
rect 7012 6817 7046 6851
rect 7046 6817 7064 6851
rect 7012 6808 7064 6817
rect 7380 6876 7432 6928
rect 10140 6876 10192 6928
rect 10692 6876 10744 6928
rect 11796 6876 11848 6928
rect 13176 6876 13228 6928
rect 9128 6851 9180 6860
rect 9128 6817 9137 6851
rect 9137 6817 9171 6851
rect 9171 6817 9180 6851
rect 9128 6808 9180 6817
rect 9772 6851 9824 6860
rect 9772 6817 9781 6851
rect 9781 6817 9815 6851
rect 9815 6817 9824 6851
rect 9772 6808 9824 6817
rect 9864 6808 9916 6860
rect 12072 6851 12124 6860
rect 4344 6672 4396 6724
rect 5724 6672 5776 6724
rect 1492 6604 1544 6656
rect 4528 6604 4580 6656
rect 5264 6647 5316 6656
rect 5264 6613 5273 6647
rect 5273 6613 5307 6647
rect 5307 6613 5316 6647
rect 5264 6604 5316 6613
rect 5632 6604 5684 6656
rect 5816 6604 5868 6656
rect 6368 6647 6420 6656
rect 6368 6613 6377 6647
rect 6377 6613 6411 6647
rect 6411 6613 6420 6647
rect 6368 6604 6420 6613
rect 9312 6783 9364 6792
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 12072 6817 12081 6851
rect 12081 6817 12115 6851
rect 12115 6817 12124 6851
rect 12072 6808 12124 6817
rect 12808 6851 12860 6860
rect 12808 6817 12817 6851
rect 12817 6817 12851 6851
rect 12851 6817 12860 6851
rect 12808 6808 12860 6817
rect 12532 6740 12584 6792
rect 13360 6808 13412 6860
rect 7656 6604 7708 6656
rect 9680 6604 9732 6656
rect 9956 6604 10008 6656
rect 10508 6604 10560 6656
rect 11152 6647 11204 6656
rect 11152 6613 11161 6647
rect 11161 6613 11195 6647
rect 11195 6613 11204 6647
rect 11152 6604 11204 6613
rect 12072 6604 12124 6656
rect 13176 6604 13228 6656
rect 3480 6502 3532 6554
rect 3544 6502 3596 6554
rect 3608 6502 3660 6554
rect 3672 6502 3724 6554
rect 8478 6502 8530 6554
rect 8542 6502 8594 6554
rect 8606 6502 8658 6554
rect 8670 6502 8722 6554
rect 13475 6502 13527 6554
rect 13539 6502 13591 6554
rect 13603 6502 13655 6554
rect 13667 6502 13719 6554
rect 4068 6400 4120 6452
rect 5908 6400 5960 6452
rect 7104 6400 7156 6452
rect 8024 6400 8076 6452
rect 8208 6400 8260 6452
rect 6460 6332 6512 6384
rect 8300 6332 8352 6384
rect 8760 6332 8812 6384
rect 3056 6264 3108 6316
rect 6276 6264 6328 6316
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 10784 6400 10836 6452
rect 9312 6264 9364 6316
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 9864 6307 9916 6316
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 9864 6264 9916 6273
rect 11152 6264 11204 6316
rect 12808 6264 12860 6316
rect 1492 6239 1544 6248
rect 1492 6205 1501 6239
rect 1501 6205 1535 6239
rect 1535 6205 1544 6239
rect 1492 6196 1544 6205
rect 4896 6239 4948 6248
rect 4896 6205 4930 6239
rect 4930 6205 4948 6239
rect 2964 6128 3016 6180
rect 3424 6171 3476 6180
rect 3424 6137 3458 6171
rect 3458 6137 3476 6171
rect 3424 6128 3476 6137
rect 4896 6196 4948 6205
rect 5448 6128 5500 6180
rect 6644 6128 6696 6180
rect 5172 6060 5224 6112
rect 7104 6196 7156 6248
rect 8944 6196 8996 6248
rect 9220 6196 9272 6248
rect 10600 6239 10652 6248
rect 10600 6205 10609 6239
rect 10609 6205 10643 6239
rect 10643 6205 10652 6239
rect 10600 6196 10652 6205
rect 7196 6103 7248 6112
rect 7196 6069 7205 6103
rect 7205 6069 7239 6103
rect 7239 6069 7248 6103
rect 7196 6060 7248 6069
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7748 6103 7800 6112
rect 7288 6060 7340 6069
rect 7748 6069 7757 6103
rect 7757 6069 7791 6103
rect 7791 6069 7800 6103
rect 7748 6060 7800 6069
rect 8300 6060 8352 6112
rect 9496 6060 9548 6112
rect 5979 5958 6031 6010
rect 6043 5958 6095 6010
rect 6107 5958 6159 6010
rect 6171 5958 6223 6010
rect 10976 5958 11028 6010
rect 11040 5958 11092 6010
rect 11104 5958 11156 6010
rect 11168 5958 11220 6010
rect 3332 5856 3384 5908
rect 4712 5856 4764 5908
rect 6828 5856 6880 5908
rect 8760 5856 8812 5908
rect 10048 5856 10100 5908
rect 3056 5788 3108 5840
rect 5724 5831 5776 5840
rect 2136 5720 2188 5772
rect 2780 5720 2832 5772
rect 3240 5720 3292 5772
rect 5172 5763 5224 5772
rect 5172 5729 5181 5763
rect 5181 5729 5215 5763
rect 5215 5729 5224 5763
rect 5172 5720 5224 5729
rect 5724 5797 5758 5831
rect 5758 5797 5776 5831
rect 5724 5788 5776 5797
rect 7932 5788 7984 5840
rect 10324 5788 10376 5840
rect 10692 5788 10744 5840
rect 7380 5763 7432 5772
rect 7380 5729 7389 5763
rect 7389 5729 7423 5763
rect 7423 5729 7432 5763
rect 7380 5720 7432 5729
rect 8852 5720 8904 5772
rect 9128 5720 9180 5772
rect 9404 5720 9456 5772
rect 9864 5720 9916 5772
rect 10048 5720 10100 5772
rect 5448 5695 5500 5704
rect 3424 5627 3476 5636
rect 3424 5593 3433 5627
rect 3433 5593 3467 5627
rect 3467 5593 3476 5627
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 6920 5652 6972 5704
rect 7472 5652 7524 5704
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 3424 5584 3476 5593
rect 7012 5584 7064 5636
rect 8208 5584 8260 5636
rect 4712 5516 4764 5568
rect 7748 5516 7800 5568
rect 9128 5516 9180 5568
rect 9496 5516 9548 5568
rect 3480 5414 3532 5466
rect 3544 5414 3596 5466
rect 3608 5414 3660 5466
rect 3672 5414 3724 5466
rect 8478 5414 8530 5466
rect 8542 5414 8594 5466
rect 8606 5414 8658 5466
rect 8670 5414 8722 5466
rect 13475 5414 13527 5466
rect 13539 5414 13591 5466
rect 13603 5414 13655 5466
rect 13667 5414 13719 5466
rect 5632 5312 5684 5364
rect 5724 5312 5776 5364
rect 6368 5355 6420 5364
rect 6368 5321 6377 5355
rect 6377 5321 6411 5355
rect 6411 5321 6420 5355
rect 6368 5312 6420 5321
rect 7472 5312 7524 5364
rect 6828 5244 6880 5296
rect 2228 5219 2280 5228
rect 2228 5185 2237 5219
rect 2237 5185 2271 5219
rect 2271 5185 2280 5219
rect 2228 5176 2280 5185
rect 6736 5176 6788 5228
rect 2136 5108 2188 5160
rect 4528 5151 4580 5160
rect 1768 5083 1820 5092
rect 1768 5049 1777 5083
rect 1777 5049 1811 5083
rect 1811 5049 1820 5083
rect 1768 5040 1820 5049
rect 4160 5040 4212 5092
rect 3332 4972 3384 5024
rect 3976 4972 4028 5024
rect 4528 5117 4537 5151
rect 4537 5117 4571 5151
rect 4571 5117 4580 5151
rect 4528 5108 4580 5117
rect 5448 5108 5500 5160
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 8944 5312 8996 5364
rect 9496 5312 9548 5364
rect 9680 5312 9732 5364
rect 12072 5312 12124 5364
rect 14832 5355 14884 5364
rect 14832 5321 14841 5355
rect 14841 5321 14875 5355
rect 14875 5321 14884 5355
rect 14832 5312 14884 5321
rect 12348 5176 12400 5228
rect 13360 5176 13412 5228
rect 6920 5040 6972 5092
rect 8208 5040 8260 5092
rect 9312 5108 9364 5160
rect 10048 5151 10100 5160
rect 10048 5117 10057 5151
rect 10057 5117 10091 5151
rect 10091 5117 10100 5151
rect 10048 5108 10100 5117
rect 11336 5108 11388 5160
rect 12440 5108 12492 5160
rect 12900 5151 12952 5160
rect 12900 5117 12909 5151
rect 12909 5117 12943 5151
rect 12943 5117 12952 5151
rect 12900 5108 12952 5117
rect 14832 5108 14884 5160
rect 9404 5040 9456 5092
rect 10324 5083 10376 5092
rect 10324 5049 10358 5083
rect 10358 5049 10376 5083
rect 10324 5040 10376 5049
rect 16212 5040 16264 5092
rect 5264 4972 5316 5024
rect 7012 4972 7064 5024
rect 8576 4972 8628 5024
rect 10692 4972 10744 5024
rect 12624 4972 12676 5024
rect 5979 4870 6031 4922
rect 6043 4870 6095 4922
rect 6107 4870 6159 4922
rect 6171 4870 6223 4922
rect 10976 4870 11028 4922
rect 11040 4870 11092 4922
rect 11104 4870 11156 4922
rect 11168 4870 11220 4922
rect 2780 4811 2832 4820
rect 2780 4777 2789 4811
rect 2789 4777 2823 4811
rect 2823 4777 2832 4811
rect 2780 4768 2832 4777
rect 4804 4811 4856 4820
rect 4804 4777 4813 4811
rect 4813 4777 4847 4811
rect 4847 4777 4856 4811
rect 4804 4768 4856 4777
rect 2136 4700 2188 4752
rect 5264 4768 5316 4820
rect 6276 4768 6328 4820
rect 6552 4811 6604 4820
rect 6552 4777 6561 4811
rect 6561 4777 6595 4811
rect 6595 4777 6604 4811
rect 6552 4768 6604 4777
rect 7288 4768 7340 4820
rect 7380 4768 7432 4820
rect 8300 4768 8352 4820
rect 8852 4768 8904 4820
rect 9220 4811 9272 4820
rect 9220 4777 9229 4811
rect 9229 4777 9263 4811
rect 9263 4777 9272 4811
rect 9220 4768 9272 4777
rect 9588 4768 9640 4820
rect 1492 4632 1544 4684
rect 4252 4675 4304 4684
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 6644 4632 6696 4684
rect 7840 4675 7892 4684
rect 7840 4641 7849 4675
rect 7849 4641 7883 4675
rect 7883 4641 7892 4675
rect 7840 4632 7892 4641
rect 3976 4564 4028 4616
rect 4160 4564 4212 4616
rect 7472 4607 7524 4616
rect 2688 4428 2740 4480
rect 3148 4471 3200 4480
rect 3148 4437 3157 4471
rect 3157 4437 3191 4471
rect 3191 4437 3200 4471
rect 3148 4428 3200 4437
rect 4988 4496 5040 4548
rect 4620 4428 4672 4480
rect 6276 4471 6328 4480
rect 6276 4437 6285 4471
rect 6285 4437 6319 4471
rect 6319 4437 6328 4471
rect 6276 4428 6328 4437
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 8576 4607 8628 4616
rect 8576 4573 8585 4607
rect 8585 4573 8619 4607
rect 8619 4573 8628 4607
rect 8576 4564 8628 4573
rect 7656 4496 7708 4548
rect 10140 4700 10192 4752
rect 11428 4768 11480 4820
rect 12716 4768 12768 4820
rect 13452 4768 13504 4820
rect 10324 4700 10376 4752
rect 9956 4632 10008 4684
rect 10784 4675 10836 4684
rect 10784 4641 10793 4675
rect 10793 4641 10827 4675
rect 10827 4641 10836 4675
rect 10784 4632 10836 4641
rect 9312 4607 9364 4616
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 9588 4564 9640 4616
rect 10416 4564 10468 4616
rect 10876 4607 10928 4616
rect 10876 4573 10885 4607
rect 10885 4573 10919 4607
rect 10919 4573 10928 4607
rect 10876 4564 10928 4573
rect 12808 4700 12860 4752
rect 14740 4768 14792 4820
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 12348 4632 12400 4684
rect 12716 4632 12768 4684
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 10324 4496 10376 4548
rect 13452 4496 13504 4548
rect 7932 4428 7984 4480
rect 9404 4428 9456 4480
rect 10416 4471 10468 4480
rect 10416 4437 10425 4471
rect 10425 4437 10459 4471
rect 10459 4437 10468 4471
rect 10416 4428 10468 4437
rect 12716 4471 12768 4480
rect 12716 4437 12725 4471
rect 12725 4437 12759 4471
rect 12759 4437 12768 4471
rect 12716 4428 12768 4437
rect 12808 4471 12860 4480
rect 12808 4437 12817 4471
rect 12817 4437 12851 4471
rect 12851 4437 12860 4471
rect 12808 4428 12860 4437
rect 13360 4428 13412 4480
rect 3480 4326 3532 4378
rect 3544 4326 3596 4378
rect 3608 4326 3660 4378
rect 3672 4326 3724 4378
rect 8478 4326 8530 4378
rect 8542 4326 8594 4378
rect 8606 4326 8658 4378
rect 8670 4326 8722 4378
rect 13475 4326 13527 4378
rect 13539 4326 13591 4378
rect 13603 4326 13655 4378
rect 13667 4326 13719 4378
rect 2504 4224 2556 4276
rect 3332 4224 3384 4276
rect 10784 4267 10836 4276
rect 10784 4233 10793 4267
rect 10793 4233 10827 4267
rect 10827 4233 10836 4267
rect 10784 4224 10836 4233
rect 2780 4156 2832 4208
rect 5540 4156 5592 4208
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 3148 4020 3200 4072
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 5540 4063 5592 4072
rect 2412 3884 2464 3936
rect 2780 3884 2832 3936
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 5356 3884 5408 3936
rect 5540 3884 5592 3936
rect 6368 4156 6420 4208
rect 6460 4131 6512 4140
rect 6460 4097 6469 4131
rect 6469 4097 6503 4131
rect 6503 4097 6512 4131
rect 6460 4088 6512 4097
rect 6736 4088 6788 4140
rect 7656 4156 7708 4208
rect 8760 4156 8812 4208
rect 10232 4156 10284 4208
rect 8208 4088 8260 4140
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 10692 4156 10744 4208
rect 12716 4156 12768 4208
rect 11428 4131 11480 4140
rect 11428 4097 11437 4131
rect 11437 4097 11471 4131
rect 11471 4097 11480 4131
rect 11428 4088 11480 4097
rect 12348 4088 12400 4140
rect 12808 4088 12860 4140
rect 6368 4020 6420 4072
rect 7380 4020 7432 4072
rect 6000 3952 6052 4004
rect 9036 4020 9088 4072
rect 9956 4020 10008 4072
rect 12072 4020 12124 4072
rect 5816 3884 5868 3936
rect 6552 3884 6604 3936
rect 7196 3884 7248 3936
rect 7288 3884 7340 3936
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 8300 3884 8352 3936
rect 8944 3927 8996 3936
rect 8944 3893 8953 3927
rect 8953 3893 8987 3927
rect 8987 3893 8996 3927
rect 8944 3884 8996 3893
rect 9036 3927 9088 3936
rect 9036 3893 9045 3927
rect 9045 3893 9079 3927
rect 9079 3893 9088 3927
rect 9036 3884 9088 3893
rect 9220 3884 9272 3936
rect 10508 3884 10560 3936
rect 10692 3884 10744 3936
rect 11520 3884 11572 3936
rect 12072 3884 12124 3936
rect 12624 3952 12676 4004
rect 5979 3782 6031 3834
rect 6043 3782 6095 3834
rect 6107 3782 6159 3834
rect 6171 3782 6223 3834
rect 10976 3782 11028 3834
rect 11040 3782 11092 3834
rect 11104 3782 11156 3834
rect 11168 3782 11220 3834
rect 3240 3680 3292 3732
rect 5264 3680 5316 3732
rect 4436 3612 4488 3664
rect 1860 3544 1912 3596
rect 2412 3544 2464 3596
rect 3056 3587 3108 3596
rect 3056 3553 3065 3587
rect 3065 3553 3099 3587
rect 3099 3553 3108 3587
rect 3056 3544 3108 3553
rect 4528 3544 4580 3596
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 2780 3476 2832 3528
rect 3148 3476 3200 3528
rect 4712 3476 4764 3528
rect 1952 3408 2004 3460
rect 5816 3680 5868 3732
rect 7932 3680 7984 3732
rect 8760 3680 8812 3732
rect 8852 3680 8904 3732
rect 10140 3723 10192 3732
rect 10140 3689 10149 3723
rect 10149 3689 10183 3723
rect 10183 3689 10192 3723
rect 10140 3680 10192 3689
rect 10876 3680 10928 3732
rect 11336 3680 11388 3732
rect 11612 3680 11664 3732
rect 11796 3680 11848 3732
rect 12348 3680 12400 3732
rect 6460 3612 6512 3664
rect 7472 3655 7524 3664
rect 7472 3621 7481 3655
rect 7481 3621 7515 3655
rect 7515 3621 7524 3655
rect 7472 3612 7524 3621
rect 7196 3544 7248 3596
rect 7656 3612 7708 3664
rect 8208 3612 8260 3664
rect 9496 3612 9548 3664
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 5172 3476 5224 3528
rect 5448 3476 5500 3528
rect 7012 3476 7064 3528
rect 9404 3544 9456 3596
rect 9772 3544 9824 3596
rect 10876 3544 10928 3596
rect 11336 3544 11388 3596
rect 12624 3612 12676 3664
rect 13084 3612 13136 3664
rect 11612 3544 11664 3596
rect 7840 3476 7892 3528
rect 9588 3476 9640 3528
rect 10968 3476 11020 3528
rect 11428 3476 11480 3528
rect 1400 3340 1452 3392
rect 2320 3340 2372 3392
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 4712 3340 4764 3392
rect 5264 3340 5316 3392
rect 5540 3340 5592 3392
rect 7288 3408 7340 3460
rect 7472 3408 7524 3460
rect 7656 3408 7708 3460
rect 6552 3340 6604 3392
rect 7380 3340 7432 3392
rect 7840 3340 7892 3392
rect 9220 3340 9272 3392
rect 9496 3383 9548 3392
rect 9496 3349 9505 3383
rect 9505 3349 9539 3383
rect 9539 3349 9548 3383
rect 9496 3340 9548 3349
rect 9864 3340 9916 3392
rect 11704 3340 11756 3392
rect 3480 3238 3532 3290
rect 3544 3238 3596 3290
rect 3608 3238 3660 3290
rect 3672 3238 3724 3290
rect 8478 3238 8530 3290
rect 8542 3238 8594 3290
rect 8606 3238 8658 3290
rect 8670 3238 8722 3290
rect 13475 3238 13527 3290
rect 13539 3238 13591 3290
rect 13603 3238 13655 3290
rect 13667 3238 13719 3290
rect 3240 3136 3292 3188
rect 4712 3136 4764 3188
rect 4988 3136 5040 3188
rect 5356 3179 5408 3188
rect 5356 3145 5365 3179
rect 5365 3145 5399 3179
rect 5399 3145 5408 3179
rect 5356 3136 5408 3145
rect 5816 3136 5868 3188
rect 6460 3136 6512 3188
rect 6828 3136 6880 3188
rect 8024 3136 8076 3188
rect 8116 3136 8168 3188
rect 9128 3136 9180 3188
rect 10968 3179 11020 3188
rect 10968 3145 10977 3179
rect 10977 3145 11011 3179
rect 11011 3145 11020 3179
rect 10968 3136 11020 3145
rect 11520 3136 11572 3188
rect 4804 3068 4856 3120
rect 4896 3068 4948 3120
rect 8208 3111 8260 3120
rect 8208 3077 8217 3111
rect 8217 3077 8251 3111
rect 8251 3077 8260 3111
rect 8208 3068 8260 3077
rect 8576 3068 8628 3120
rect 9036 3068 9088 3120
rect 1492 3000 1544 3052
rect 5080 3043 5132 3052
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 6460 3000 6512 3052
rect 1492 2907 1544 2916
rect 1492 2873 1501 2907
rect 1501 2873 1535 2907
rect 1535 2873 1544 2907
rect 5816 2932 5868 2984
rect 6184 2975 6236 2984
rect 6184 2941 6193 2975
rect 6193 2941 6227 2975
rect 6227 2941 6236 2975
rect 6184 2932 6236 2941
rect 6736 2932 6788 2984
rect 1492 2864 1544 2873
rect 3148 2796 3200 2848
rect 6460 2864 6512 2916
rect 7840 3000 7892 3052
rect 7380 2932 7432 2984
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 11612 3000 11664 3052
rect 16948 3000 17000 3052
rect 7012 2864 7064 2916
rect 7196 2864 7248 2916
rect 9956 2932 10008 2984
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 14648 2932 14700 2984
rect 8668 2907 8720 2916
rect 8668 2873 8677 2907
rect 8677 2873 8711 2907
rect 8711 2873 8720 2907
rect 8668 2864 8720 2873
rect 8852 2864 8904 2916
rect 9496 2864 9548 2916
rect 9772 2864 9824 2916
rect 12164 2907 12216 2916
rect 12164 2873 12173 2907
rect 12173 2873 12207 2907
rect 12207 2873 12216 2907
rect 12164 2864 12216 2873
rect 4528 2839 4580 2848
rect 4528 2805 4537 2839
rect 4537 2805 4571 2839
rect 4571 2805 4580 2839
rect 4528 2796 4580 2805
rect 4804 2796 4856 2848
rect 5448 2796 5500 2848
rect 6828 2796 6880 2848
rect 8760 2839 8812 2848
rect 8760 2805 8769 2839
rect 8769 2805 8803 2839
rect 8803 2805 8812 2839
rect 8760 2796 8812 2805
rect 10232 2796 10284 2848
rect 12256 2796 12308 2848
rect 12440 2796 12492 2848
rect 12992 2796 13044 2848
rect 15936 2864 15988 2916
rect 15200 2796 15252 2848
rect 5979 2694 6031 2746
rect 6043 2694 6095 2746
rect 6107 2694 6159 2746
rect 6171 2694 6223 2746
rect 10976 2694 11028 2746
rect 11040 2694 11092 2746
rect 11104 2694 11156 2746
rect 11168 2694 11220 2746
rect 388 2592 440 2644
rect 756 2524 808 2576
rect 3884 2592 3936 2644
rect 4528 2635 4580 2644
rect 4528 2601 4537 2635
rect 4537 2601 4571 2635
rect 4571 2601 4580 2635
rect 4528 2592 4580 2601
rect 4620 2592 4672 2644
rect 6460 2592 6512 2644
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 7748 2592 7800 2644
rect 8208 2635 8260 2644
rect 8208 2601 8217 2635
rect 8217 2601 8251 2635
rect 8251 2601 8260 2635
rect 8208 2592 8260 2601
rect 8576 2635 8628 2644
rect 8576 2601 8585 2635
rect 8585 2601 8619 2635
rect 8619 2601 8628 2635
rect 8576 2592 8628 2601
rect 9588 2592 9640 2644
rect 9956 2592 10008 2644
rect 11336 2592 11388 2644
rect 11428 2592 11480 2644
rect 12072 2592 12124 2644
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 12808 2635 12860 2644
rect 12808 2601 12817 2635
rect 12817 2601 12851 2635
rect 12851 2601 12860 2635
rect 12808 2592 12860 2601
rect 12900 2592 12952 2644
rect 14096 2592 14148 2644
rect 14832 2592 14884 2644
rect 2596 2524 2648 2576
rect 4436 2567 4488 2576
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 1952 2499 2004 2508
rect 1952 2465 1961 2499
rect 1961 2465 1995 2499
rect 1995 2465 2004 2499
rect 1952 2456 2004 2465
rect 2320 2499 2372 2508
rect 2320 2465 2329 2499
rect 2329 2465 2363 2499
rect 2363 2465 2372 2499
rect 2320 2456 2372 2465
rect 2688 2499 2740 2508
rect 2688 2465 2697 2499
rect 2697 2465 2731 2499
rect 2731 2465 2740 2499
rect 2688 2456 2740 2465
rect 3240 2456 3292 2508
rect 4436 2533 4445 2567
rect 4445 2533 4479 2567
rect 4479 2533 4488 2567
rect 4436 2524 4488 2533
rect 4344 2456 4396 2508
rect 5172 2456 5224 2508
rect 5632 2499 5684 2508
rect 5632 2465 5641 2499
rect 5641 2465 5675 2499
rect 5675 2465 5684 2499
rect 5632 2456 5684 2465
rect 5816 2456 5868 2508
rect 11980 2567 12032 2576
rect 6184 2499 6236 2508
rect 6184 2465 6193 2499
rect 6193 2465 6227 2499
rect 6227 2465 6236 2499
rect 6184 2456 6236 2465
rect 6920 2456 6972 2508
rect 8392 2456 8444 2508
rect 9220 2456 9272 2508
rect 9496 2456 9548 2508
rect 9864 2499 9916 2508
rect 9864 2465 9873 2499
rect 9873 2465 9907 2499
rect 9907 2465 9916 2499
rect 9864 2456 9916 2465
rect 11980 2533 11989 2567
rect 11989 2533 12023 2567
rect 12023 2533 12032 2567
rect 11980 2524 12032 2533
rect 2136 2388 2188 2440
rect 4712 2431 4764 2440
rect 112 2320 164 2372
rect 1860 2320 1912 2372
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 4804 2388 4856 2440
rect 5724 2388 5776 2440
rect 4160 2320 4212 2372
rect 7840 2388 7892 2440
rect 8852 2320 8904 2372
rect 11796 2456 11848 2508
rect 16580 2524 16632 2576
rect 14096 2499 14148 2508
rect 14096 2465 14105 2499
rect 14105 2465 14139 2499
rect 14139 2465 14148 2499
rect 14096 2456 14148 2465
rect 14648 2499 14700 2508
rect 14648 2465 14657 2499
rect 14657 2465 14691 2499
rect 14691 2465 14700 2499
rect 14648 2456 14700 2465
rect 11244 2388 11296 2440
rect 11612 2431 11664 2440
rect 11612 2397 11621 2431
rect 11621 2397 11655 2431
rect 11655 2397 11664 2431
rect 11612 2388 11664 2397
rect 15568 2388 15620 2440
rect 12440 2320 12492 2372
rect 1124 2252 1176 2304
rect 3792 2252 3844 2304
rect 8944 2252 8996 2304
rect 9128 2252 9180 2304
rect 10784 2295 10836 2304
rect 10784 2261 10793 2295
rect 10793 2261 10827 2295
rect 10827 2261 10836 2295
rect 10784 2252 10836 2261
rect 11244 2252 11296 2304
rect 11980 2252 12032 2304
rect 3480 2150 3532 2202
rect 3544 2150 3596 2202
rect 3608 2150 3660 2202
rect 3672 2150 3724 2202
rect 8478 2150 8530 2202
rect 8542 2150 8594 2202
rect 8606 2150 8658 2202
rect 8670 2150 8722 2202
rect 13475 2150 13527 2202
rect 13539 2150 13591 2202
rect 13603 2150 13655 2202
rect 13667 2150 13719 2202
rect 3884 2048 3936 2100
rect 9128 2048 9180 2100
rect 8024 1980 8076 2032
rect 10692 2048 10744 2100
rect 11244 2048 11296 2100
rect 9496 1980 9548 2032
rect 11704 1980 11756 2032
rect 2504 1912 2556 1964
rect 10784 1912 10836 1964
rect 6184 1844 6236 1896
rect 7564 1844 7616 1896
rect 11980 1844 12032 1896
rect 7104 1776 7156 1828
rect 8668 1776 8720 1828
rect 10324 1776 10376 1828
rect 12440 1776 12492 1828
rect 9312 1708 9364 1760
rect 12164 1708 12216 1760
rect 5264 1504 5316 1556
rect 7196 1504 7248 1556
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 938 19200 994 20000
rect 1306 19200 1362 20000
rect 1674 19200 1730 20000
rect 1950 19408 2006 19417
rect 1950 19343 2006 19352
rect 216 16114 244 19200
rect 204 16108 256 16114
rect 204 16050 256 16056
rect 584 16017 612 19200
rect 952 17270 980 19200
rect 1320 17610 1348 19200
rect 1688 18578 1716 19200
rect 1688 18550 1808 18578
rect 1674 18456 1730 18465
rect 1674 18391 1730 18400
rect 1308 17604 1360 17610
rect 1308 17546 1360 17552
rect 940 17264 992 17270
rect 940 17206 992 17212
rect 1688 17202 1716 18391
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1596 16538 1624 17070
rect 1780 16561 1808 18550
rect 1964 17134 1992 19343
rect 2042 19200 2098 20000
rect 2410 19200 2466 20000
rect 2778 19200 2834 20000
rect 3146 19200 3202 20000
rect 3514 19200 3570 20000
rect 3882 19200 3938 20000
rect 4250 19200 4306 20000
rect 4618 19200 4674 20000
rect 4986 19200 5042 20000
rect 5354 19200 5410 20000
rect 5722 19200 5778 20000
rect 6182 19200 6238 20000
rect 6550 19200 6606 20000
rect 6918 19200 6974 20000
rect 7286 19200 7342 20000
rect 7654 19200 7710 20000
rect 8022 19200 8078 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 9126 19200 9182 20000
rect 9494 19200 9550 20000
rect 9862 19200 9918 20000
rect 10230 19200 10286 20000
rect 10598 19200 10654 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11794 19200 11850 20000
rect 12162 19200 12218 20000
rect 12530 19200 12586 20000
rect 12898 19200 12954 20000
rect 13266 19200 13322 20000
rect 13634 19200 13690 20000
rect 14002 19200 14058 20000
rect 14370 19200 14426 20000
rect 14738 19200 14794 20000
rect 15106 19200 15162 20000
rect 15474 19200 15530 20000
rect 15842 19200 15898 20000
rect 16210 19200 16266 20000
rect 16578 19200 16634 20000
rect 16946 19200 17002 20000
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 2056 16726 2084 19200
rect 2044 16720 2096 16726
rect 2044 16662 2096 16668
rect 1412 16510 1624 16538
rect 1766 16552 1822 16561
rect 570 16008 626 16017
rect 570 15943 626 15952
rect 1412 8412 1440 16510
rect 1766 16487 1822 16496
rect 1766 16416 1822 16425
rect 1766 16351 1822 16360
rect 1492 16244 1544 16250
rect 1492 16186 1544 16192
rect 1504 15570 1532 16186
rect 1492 15564 1544 15570
rect 1492 15506 1544 15512
rect 1676 15496 1728 15502
rect 1674 15464 1676 15473
rect 1728 15464 1730 15473
rect 1674 15399 1730 15408
rect 1780 14958 1808 16351
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1676 14408 1728 14414
rect 1674 14376 1676 14385
rect 1728 14376 1730 14385
rect 1674 14311 1730 14320
rect 1584 14272 1636 14278
rect 1584 14214 1636 14220
rect 1596 13870 1624 14214
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1872 13433 1900 13806
rect 1858 13424 1914 13433
rect 1858 13359 1914 13368
rect 1766 12472 1822 12481
rect 1766 12407 1822 12416
rect 1780 12374 1808 12407
rect 1768 12368 1820 12374
rect 1768 12310 1820 12316
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11694 1532 12038
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 1768 11620 1820 11626
rect 1768 11562 1820 11568
rect 1780 11393 1808 11562
rect 1766 11384 1822 11393
rect 2056 11354 2084 11630
rect 1766 11319 1822 11328
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1490 9616 1546 9625
rect 1490 9551 1546 9560
rect 1504 9518 1532 9551
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1596 9178 1624 11086
rect 1872 10810 1900 11154
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2148 10130 2176 10610
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 1768 9444 1820 9450
rect 1768 9386 1820 9392
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1584 8424 1636 8430
rect 1412 8384 1584 8412
rect 1780 8401 1808 9386
rect 2056 8430 2084 9454
rect 2148 9382 2176 10066
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2148 8974 2176 9318
rect 2240 9178 2268 10406
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2044 8424 2096 8430
rect 1584 8366 1636 8372
rect 1766 8392 1822 8401
rect 1596 8090 1624 8366
rect 2044 8366 2096 8372
rect 1766 8327 1822 8336
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 2056 7954 2084 8366
rect 2044 7948 2096 7954
rect 2044 7890 2096 7896
rect 1674 7440 1730 7449
rect 1674 7375 1676 7384
rect 1728 7375 1730 7384
rect 1676 7346 1728 7352
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1504 6254 1532 6598
rect 1688 6497 1716 6734
rect 1674 6488 1730 6497
rect 1674 6423 1730 6432
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2148 5166 2176 5714
rect 2226 5400 2282 5409
rect 2226 5335 2282 5344
rect 2240 5234 2268 5335
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 1768 5092 1820 5098
rect 1768 5034 1820 5040
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 388 2644 440 2650
rect 388 2586 440 2592
rect 112 2372 164 2378
rect 112 2314 164 2320
rect 124 800 152 2314
rect 400 800 428 2586
rect 756 2576 808 2582
rect 756 2518 808 2524
rect 768 800 796 2518
rect 1124 2304 1176 2310
rect 1124 2246 1176 2252
rect 1136 800 1164 2246
rect 1412 800 1440 3334
rect 1504 3058 1532 4626
rect 1780 4457 1808 5034
rect 2148 4758 2176 5102
rect 2136 4752 2188 4758
rect 2332 4729 2360 15846
rect 2424 15706 2452 19200
rect 2504 17264 2556 17270
rect 2504 17206 2556 17212
rect 2516 17066 2544 17206
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 2516 16794 2544 17002
rect 2792 16794 2820 19200
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 3160 16522 3188 19200
rect 3528 17626 3556 19200
rect 3528 17598 3832 17626
rect 3454 17436 3750 17456
rect 3510 17434 3534 17436
rect 3590 17434 3614 17436
rect 3670 17434 3694 17436
rect 3532 17382 3534 17434
rect 3596 17382 3608 17434
rect 3670 17382 3672 17434
rect 3510 17380 3534 17382
rect 3590 17380 3614 17382
rect 3670 17380 3694 17382
rect 3454 17360 3750 17380
rect 3804 16794 3832 17598
rect 3792 16788 3844 16794
rect 3792 16730 3844 16736
rect 3422 16688 3478 16697
rect 3422 16623 3424 16632
rect 3476 16623 3478 16632
rect 3424 16594 3476 16600
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3148 16516 3200 16522
rect 3148 16458 3200 16464
rect 3454 16348 3750 16368
rect 3510 16346 3534 16348
rect 3590 16346 3614 16348
rect 3670 16346 3694 16348
rect 3532 16294 3534 16346
rect 3596 16294 3608 16346
rect 3670 16294 3672 16346
rect 3510 16292 3534 16294
rect 3590 16292 3614 16294
rect 3670 16292 3694 16294
rect 3454 16272 3750 16292
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2700 14822 2728 15982
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2872 15428 2924 15434
rect 2872 15370 2924 15376
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2700 13938 2728 14758
rect 2884 14482 2912 15370
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2976 14074 3004 15506
rect 3344 15162 3372 15914
rect 3454 15260 3750 15280
rect 3510 15258 3534 15260
rect 3590 15258 3614 15260
rect 3670 15258 3694 15260
rect 3532 15206 3534 15258
rect 3596 15206 3608 15258
rect 3670 15206 3672 15258
rect 3510 15204 3534 15206
rect 3590 15204 3614 15206
rect 3670 15204 3694 15206
rect 3454 15184 3750 15204
rect 3332 15156 3384 15162
rect 3332 15098 3384 15104
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2700 13410 2728 13874
rect 2608 13394 2728 13410
rect 2596 13388 2728 13394
rect 2648 13382 2728 13388
rect 2596 13330 2648 13336
rect 3068 12986 3096 14418
rect 3252 14414 3280 14826
rect 3804 14822 3832 16526
rect 3896 16522 3924 19200
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3988 16697 4016 16934
rect 4264 16776 4292 19200
rect 4632 17338 4660 19200
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 4344 16788 4396 16794
rect 4264 16748 4344 16776
rect 4344 16730 4396 16736
rect 3974 16688 4030 16697
rect 4448 16658 4476 17138
rect 5000 16998 5028 19200
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 5368 17626 5396 19200
rect 5276 17134 5304 17614
rect 5368 17598 5580 17626
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5552 16726 5580 17598
rect 5736 17338 5764 19200
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 6196 17082 6224 19200
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6380 17338 6408 17614
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6196 17054 6408 17082
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 3974 16623 4030 16632
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 3884 16516 3936 16522
rect 3884 16458 3936 16464
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4356 15178 4384 15438
rect 4356 15150 4476 15178
rect 4540 15162 4568 15438
rect 4448 15094 4476 15150
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4436 15088 4488 15094
rect 4436 15030 4488 15036
rect 4436 14884 4488 14890
rect 4436 14826 4488 14832
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3252 13530 3280 14350
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 3454 14172 3750 14192
rect 3510 14170 3534 14172
rect 3590 14170 3614 14172
rect 3670 14170 3694 14172
rect 3532 14118 3534 14170
rect 3596 14118 3608 14170
rect 3670 14118 3672 14170
rect 3510 14116 3534 14118
rect 3590 14116 3614 14118
rect 3670 14116 3694 14118
rect 3454 14096 3750 14116
rect 4080 14074 4108 14282
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3454 13084 3750 13104
rect 3510 13082 3534 13084
rect 3590 13082 3614 13084
rect 3670 13082 3694 13084
rect 3532 13030 3534 13082
rect 3596 13030 3608 13082
rect 3670 13030 3672 13082
rect 3510 13028 3534 13030
rect 3590 13028 3614 13030
rect 3670 13028 3694 13030
rect 3454 13008 3750 13028
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 3454 11996 3750 12016
rect 3510 11994 3534 11996
rect 3590 11994 3614 11996
rect 3670 11994 3694 11996
rect 3532 11942 3534 11994
rect 3596 11942 3608 11994
rect 3670 11942 3672 11994
rect 3510 11940 3534 11942
rect 3590 11940 3614 11942
rect 3670 11940 3694 11942
rect 3454 11920 3750 11940
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2424 11150 2452 11630
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 3792 11620 3844 11626
rect 3792 11562 3844 11568
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2424 10198 2452 11086
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2412 10192 2464 10198
rect 2412 10134 2464 10140
rect 2608 9450 2636 10542
rect 2792 10441 2820 11562
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 2778 10432 2834 10441
rect 2778 10367 2834 10376
rect 2976 10266 3004 11154
rect 3160 10742 3188 11494
rect 3804 11354 3832 11562
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3454 10908 3750 10928
rect 3510 10906 3534 10908
rect 3590 10906 3614 10908
rect 3670 10906 3694 10908
rect 3532 10854 3534 10906
rect 3596 10854 3608 10906
rect 3670 10854 3672 10906
rect 3510 10852 3534 10854
rect 3590 10852 3614 10854
rect 3670 10852 3694 10854
rect 3454 10832 3750 10852
rect 3148 10736 3200 10742
rect 3148 10678 3200 10684
rect 3700 10668 3752 10674
rect 3752 10628 3832 10656
rect 3700 10610 3752 10616
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2976 9568 3004 9862
rect 2884 9540 3004 9568
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 2502 9072 2558 9081
rect 2502 9007 2558 9016
rect 2136 4694 2188 4700
rect 2318 4720 2374 4729
rect 2318 4655 2374 4664
rect 1766 4448 1822 4457
rect 1766 4383 1822 4392
rect 2516 4282 2544 9007
rect 2608 8974 2636 9386
rect 2884 9110 2912 9540
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2700 8838 2728 8978
rect 2792 8945 2820 8978
rect 2778 8936 2834 8945
rect 3068 8906 3096 10406
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3160 9178 3188 9454
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3344 9110 3372 10474
rect 3804 10062 3832 10628
rect 3884 10192 3936 10198
rect 3884 10134 3936 10140
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3454 9820 3750 9840
rect 3510 9818 3534 9820
rect 3590 9818 3614 9820
rect 3670 9818 3694 9820
rect 3532 9766 3534 9818
rect 3596 9766 3608 9818
rect 3670 9766 3672 9818
rect 3510 9764 3534 9766
rect 3590 9764 3614 9766
rect 3670 9764 3694 9766
rect 3454 9744 3750 9764
rect 3804 9654 3832 9998
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3712 9489 3740 9522
rect 3698 9480 3754 9489
rect 3698 9415 3754 9424
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 2778 8871 2834 8880
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 3454 8732 3750 8752
rect 3510 8730 3534 8732
rect 3590 8730 3614 8732
rect 3670 8730 3694 8732
rect 3532 8678 3534 8730
rect 3596 8678 3608 8730
rect 3670 8678 3672 8730
rect 3510 8676 3534 8678
rect 3590 8676 3614 8678
rect 3670 8676 3694 8678
rect 3454 8656 3750 8676
rect 3896 8514 3924 10134
rect 3988 8537 4016 13738
rect 4080 13462 4108 14010
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 4080 12850 4108 13398
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4172 12782 4200 13670
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 3804 8486 3924 8514
rect 3974 8528 4030 8537
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2700 7002 2728 7142
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2884 6934 2912 7686
rect 2872 6928 2924 6934
rect 2872 6870 2924 6876
rect 2780 6792 2832 6798
rect 2778 6760 2780 6769
rect 2832 6760 2834 6769
rect 2778 6695 2834 6704
rect 3068 6322 3096 8230
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3146 7440 3202 7449
rect 3146 7375 3202 7384
rect 3160 7342 3188 7375
rect 3252 7342 3280 7890
rect 3344 7818 3372 8298
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3344 7410 3372 7754
rect 3454 7644 3750 7664
rect 3510 7642 3534 7644
rect 3590 7642 3614 7644
rect 3670 7642 3694 7644
rect 3532 7590 3534 7642
rect 3596 7590 3608 7642
rect 3670 7590 3672 7642
rect 3510 7588 3534 7590
rect 3590 7588 3614 7590
rect 3670 7588 3694 7590
rect 3454 7568 3750 7588
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3804 7342 3832 8486
rect 3974 8463 4030 8472
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3896 7546 3924 7822
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 4080 7392 4108 12650
rect 4264 10656 4292 14758
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4356 12782 4384 13262
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4448 11506 4476 14826
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4540 13530 4568 14350
rect 4632 14278 4660 15982
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4724 15502 4752 15846
rect 4816 15638 4844 16594
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 5000 15570 5028 16390
rect 5368 16046 5396 16526
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 5356 16040 5408 16046
rect 5408 16000 5488 16028
rect 5356 15982 5408 15988
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 4988 15564 5040 15570
rect 4988 15506 5040 15512
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 5000 15366 5028 15506
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 4816 15162 4844 15302
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 5000 15065 5028 15302
rect 4986 15056 5042 15065
rect 4986 14991 5042 15000
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4632 12714 4660 13670
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 4724 12594 4752 14010
rect 4908 13938 4936 14350
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 4908 13326 4936 13874
rect 5000 13326 5028 14214
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 4908 13190 4936 13262
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4908 12850 4936 13126
rect 5092 12986 5120 14418
rect 5276 14362 5304 15574
rect 5460 15450 5488 16000
rect 5460 15434 5580 15450
rect 5356 15428 5408 15434
rect 5460 15428 5592 15434
rect 5460 15422 5540 15428
rect 5356 15370 5408 15376
rect 5540 15370 5592 15376
rect 5368 14822 5396 15370
rect 5448 15360 5500 15366
rect 5644 15314 5672 16186
rect 5448 15302 5500 15308
rect 5460 14958 5488 15302
rect 5552 15286 5672 15314
rect 5552 15026 5580 15286
rect 5540 15020 5592 15026
rect 5540 14962 5592 14968
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5828 14482 5856 16934
rect 5953 16892 6249 16912
rect 6009 16890 6033 16892
rect 6089 16890 6113 16892
rect 6169 16890 6193 16892
rect 6031 16838 6033 16890
rect 6095 16838 6107 16890
rect 6169 16838 6171 16890
rect 6009 16836 6033 16838
rect 6089 16836 6113 16838
rect 6169 16836 6193 16838
rect 5953 16816 6249 16836
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 6012 16250 6040 16594
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5953 15804 6249 15824
rect 6009 15802 6033 15804
rect 6089 15802 6113 15804
rect 6169 15802 6193 15804
rect 6031 15750 6033 15802
rect 6095 15750 6107 15802
rect 6169 15750 6171 15802
rect 6009 15748 6033 15750
rect 6089 15748 6113 15750
rect 6169 15748 6193 15750
rect 5953 15728 6249 15748
rect 5908 15564 5960 15570
rect 5908 15506 5960 15512
rect 5920 15366 5948 15506
rect 6288 15484 6316 16934
rect 6380 16522 6408 17054
rect 6564 16794 6592 19200
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6368 16516 6420 16522
rect 6368 16458 6420 16464
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6472 15706 6500 15846
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6472 15609 6500 15642
rect 6458 15600 6514 15609
rect 6458 15535 6514 15544
rect 6564 15484 6592 15642
rect 6288 15456 6592 15484
rect 6288 15366 6316 15456
rect 5908 15360 5960 15366
rect 5908 15302 5960 15308
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 5953 14716 6249 14736
rect 6009 14714 6033 14716
rect 6089 14714 6113 14716
rect 6169 14714 6193 14716
rect 6031 14662 6033 14714
rect 6095 14662 6107 14714
rect 6169 14662 6171 14714
rect 6009 14660 6033 14662
rect 6089 14660 6113 14662
rect 6169 14660 6193 14662
rect 5953 14640 6249 14660
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5276 14334 5396 14362
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5184 13870 5212 14214
rect 5276 13870 5304 14214
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5264 13728 5316 13734
rect 5264 13670 5316 13676
rect 5276 13530 5304 13670
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5276 12986 5304 13330
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4632 12566 4752 12594
rect 4448 11478 4568 11506
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4448 10674 4476 11018
rect 4436 10668 4488 10674
rect 4264 10628 4384 10656
rect 4252 10532 4304 10538
rect 4252 10474 4304 10480
rect 4264 9518 4292 10474
rect 4356 10130 4384 10628
rect 4436 10610 4488 10616
rect 4540 10266 4568 11478
rect 4632 11354 4660 12566
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4816 11082 4844 11630
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4632 10538 4660 10746
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4816 10130 4844 11018
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4264 9178 4292 9318
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4080 7364 4200 7392
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3160 7002 3188 7142
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3252 6934 3280 7278
rect 3804 7002 3832 7278
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4080 7002 4108 7210
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 2964 6180 3016 6186
rect 2964 6122 3016 6128
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2792 4826 2820 5714
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2504 4276 2556 4282
rect 2556 4236 2636 4264
rect 2504 4218 2556 4224
rect 2608 4185 2636 4236
rect 2594 4176 2650 4185
rect 2594 4111 2650 4120
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2424 3602 2452 3878
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 1676 3528 1728 3534
rect 1674 3496 1676 3505
rect 1728 3496 1730 3505
rect 1674 3431 1730 3440
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1872 2961 1900 3538
rect 2424 3505 2452 3538
rect 2410 3496 2466 3505
rect 1952 3460 2004 3466
rect 2410 3431 2466 3440
rect 1952 3402 2004 3408
rect 1858 2952 1914 2961
rect 1492 2916 1544 2922
rect 1858 2887 1914 2896
rect 1492 2858 1544 2864
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1504 513 1532 2858
rect 1582 2816 1638 2825
rect 1582 2751 1638 2760
rect 1596 2514 1624 2751
rect 1964 2514 1992 3402
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 2514 2360 3334
rect 2608 2582 2636 4111
rect 2596 2576 2648 2582
rect 2596 2518 2648 2524
rect 2700 2514 2728 4422
rect 2792 4214 2820 4762
rect 2780 4208 2832 4214
rect 2780 4150 2832 4156
rect 2780 3936 2832 3942
rect 2832 3896 2912 3924
rect 2780 3878 2832 3884
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 1872 1170 1900 2314
rect 1780 1142 1900 1170
rect 1780 800 1808 1142
rect 2148 800 2176 2382
rect 2504 1964 2556 1970
rect 2504 1906 2556 1912
rect 2516 800 2544 1906
rect 2792 800 2820 3470
rect 2884 1465 2912 3896
rect 2976 2417 3004 6122
rect 3344 5914 3372 6802
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3454 6556 3750 6576
rect 3510 6554 3534 6556
rect 3590 6554 3614 6556
rect 3670 6554 3694 6556
rect 3532 6502 3534 6554
rect 3596 6502 3608 6554
rect 3670 6502 3672 6554
rect 3510 6500 3534 6502
rect 3590 6500 3614 6502
rect 3670 6500 3694 6502
rect 3454 6480 3750 6500
rect 4080 6458 4108 6734
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3056 5840 3108 5846
rect 3056 5782 3108 5788
rect 3068 3602 3096 5782
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3160 4078 3188 4422
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3252 3738 3280 5714
rect 3436 5642 3464 6122
rect 4172 5930 4200 7364
rect 4264 7206 4292 8774
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4356 6730 4384 9114
rect 4526 8936 4582 8945
rect 4526 8871 4582 8880
rect 4540 8838 4568 8871
rect 4632 8838 4660 9318
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4434 8528 4490 8537
rect 4540 8514 4568 8774
rect 4540 8486 4660 8514
rect 4434 8463 4490 8472
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4172 5902 4292 5930
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 3454 5468 3750 5488
rect 3510 5466 3534 5468
rect 3590 5466 3614 5468
rect 3670 5466 3694 5468
rect 3532 5414 3534 5466
rect 3596 5414 3608 5466
rect 3670 5414 3672 5466
rect 3510 5412 3534 5414
rect 3590 5412 3614 5414
rect 3670 5412 3694 5414
rect 3454 5392 3750 5412
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3344 4282 3372 4966
rect 3988 4622 4016 4966
rect 4172 4622 4200 5034
rect 4264 4690 4292 5902
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 3454 4380 3750 4400
rect 3510 4378 3534 4380
rect 3590 4378 3614 4380
rect 3670 4378 3694 4380
rect 3532 4326 3534 4378
rect 3596 4326 3608 4378
rect 3670 4326 3672 4378
rect 3510 4324 3534 4326
rect 3590 4324 3614 4326
rect 3670 4324 3694 4326
rect 3454 4304 3750 4324
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3988 4146 4016 4558
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3332 4072 3384 4078
rect 3330 4040 3332 4049
rect 3384 4040 3386 4049
rect 3330 3975 3386 3984
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3148 3528 3200 3534
rect 3200 3476 3280 3482
rect 3148 3470 3280 3476
rect 3160 3454 3280 3470
rect 3252 3194 3280 3454
rect 3454 3292 3750 3312
rect 3510 3290 3534 3292
rect 3590 3290 3614 3292
rect 3670 3290 3694 3292
rect 3532 3238 3534 3290
rect 3596 3238 3608 3290
rect 3670 3238 3672 3290
rect 3510 3236 3534 3238
rect 3590 3236 3614 3238
rect 3670 3236 3694 3238
rect 3454 3216 3750 3236
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 2962 2408 3018 2417
rect 2962 2343 3018 2352
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 3160 800 3188 2790
rect 3252 2514 3280 3130
rect 3896 2650 3924 3878
rect 4448 3670 4476 8463
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4540 6662 4568 8366
rect 4632 7750 4660 8486
rect 4816 7954 4844 9454
rect 4908 8945 4936 11494
rect 5000 11150 5028 11562
rect 5092 11218 5120 12922
rect 5368 12442 5396 14334
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5552 13462 5580 13874
rect 5736 13870 5764 14418
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5552 12850 5580 13398
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5000 10674 5028 11086
rect 5184 10810 5212 12174
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5080 9920 5132 9926
rect 5078 9888 5080 9897
rect 5132 9888 5134 9897
rect 5078 9823 5134 9832
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4894 8936 4950 8945
rect 4894 8871 4950 8880
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4632 7274 4660 7686
rect 4724 7546 4752 7890
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4540 5166 4568 6598
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4632 4486 4660 7210
rect 4908 6769 4936 8502
rect 5000 8498 5028 9454
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5000 7721 5028 8434
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 4986 7712 5042 7721
rect 4986 7647 5042 7656
rect 5092 7342 5120 7822
rect 5184 7342 5212 10610
rect 5368 10606 5396 12378
rect 5552 11218 5580 12582
rect 5828 12322 5856 14418
rect 6288 13852 6316 15302
rect 6380 14006 6408 15302
rect 6656 14906 6684 16934
rect 6840 16658 6868 17478
rect 6932 17338 6960 19200
rect 7300 17338 7328 19200
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7576 17270 7604 17682
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7102 16688 7158 16697
rect 6828 16652 6880 16658
rect 7102 16623 7158 16632
rect 6828 16594 6880 16600
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6748 15638 6776 16390
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6564 14878 6684 14906
rect 6368 14000 6420 14006
rect 6368 13942 6420 13948
rect 6564 13870 6592 14878
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6656 14006 6684 14418
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6552 13864 6604 13870
rect 6288 13824 6408 13852
rect 5953 13628 6249 13648
rect 6009 13626 6033 13628
rect 6089 13626 6113 13628
rect 6169 13626 6193 13628
rect 6031 13574 6033 13626
rect 6095 13574 6107 13626
rect 6169 13574 6171 13626
rect 6009 13572 6033 13574
rect 6089 13572 6113 13574
rect 6169 13572 6193 13574
rect 5953 13552 6249 13572
rect 5953 12540 6249 12560
rect 6009 12538 6033 12540
rect 6089 12538 6113 12540
rect 6169 12538 6193 12540
rect 6031 12486 6033 12538
rect 6095 12486 6107 12538
rect 6169 12486 6171 12538
rect 6009 12484 6033 12486
rect 6089 12484 6113 12486
rect 6169 12484 6193 12486
rect 5953 12464 6249 12484
rect 5736 12294 5856 12322
rect 6184 12300 6236 12306
rect 5736 11354 5764 12294
rect 6184 12242 6236 12248
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 6196 12186 6224 12242
rect 5816 12164 5868 12170
rect 5816 12106 5868 12112
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5644 11257 5672 11290
rect 5630 11248 5686 11257
rect 5540 11212 5592 11218
rect 5630 11183 5686 11192
rect 5540 11154 5592 11160
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 10606 5580 11018
rect 5736 10742 5764 11290
rect 5828 10810 5856 12106
rect 5920 11694 5948 12174
rect 6196 12158 6316 12186
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 6288 11558 6316 12158
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 5953 11452 6249 11472
rect 6009 11450 6033 11452
rect 6089 11450 6113 11452
rect 6169 11450 6193 11452
rect 6031 11398 6033 11450
rect 6095 11398 6107 11450
rect 6169 11398 6171 11450
rect 6009 11396 6033 11398
rect 6089 11396 6113 11398
rect 6169 11396 6193 11398
rect 5953 11376 6249 11396
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5814 10704 5870 10713
rect 5814 10639 5870 10648
rect 5356 10600 5408 10606
rect 5276 10560 5356 10588
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 4894 6760 4950 6769
rect 4894 6695 4950 6704
rect 4908 6254 4936 6695
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4724 5574 4752 5850
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4802 5264 4858 5273
rect 4802 5199 4858 5208
rect 4816 4826 4844 5199
rect 4804 4820 4856 4826
rect 4724 4780 4804 4808
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4436 3664 4488 3670
rect 4356 3624 4436 3652
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 4356 2514 4384 3624
rect 4436 3606 4488 3612
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4448 2582 4476 3334
rect 4540 3233 4568 3538
rect 4724 3534 4752 4780
rect 4804 4762 4856 4768
rect 5000 4706 5028 6870
rect 5276 6662 5304 10560
rect 5356 10542 5408 10548
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 9518 5396 9862
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5552 9466 5580 10134
rect 5632 9512 5684 9518
rect 5552 9460 5632 9466
rect 5552 9454 5684 9460
rect 5552 9438 5672 9454
rect 5552 9160 5580 9438
rect 5460 9132 5580 9160
rect 5460 9042 5488 9132
rect 5828 9081 5856 10639
rect 5920 10606 5948 11154
rect 6288 10674 6316 11494
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5953 10364 6249 10384
rect 6009 10362 6033 10364
rect 6089 10362 6113 10364
rect 6169 10362 6193 10364
rect 6031 10310 6033 10362
rect 6095 10310 6107 10362
rect 6169 10310 6171 10362
rect 6009 10308 6033 10310
rect 6089 10308 6113 10310
rect 6169 10308 6193 10310
rect 5953 10288 6249 10308
rect 6380 9466 6408 13824
rect 6552 13806 6604 13812
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6472 12646 6500 12786
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6472 11286 6500 12242
rect 6460 11280 6512 11286
rect 6460 11222 6512 11228
rect 6472 10470 6500 11222
rect 6460 10464 6512 10470
rect 6458 10432 6460 10441
rect 6512 10432 6514 10441
rect 6458 10367 6514 10376
rect 6564 9654 6592 13806
rect 6748 13734 6776 14962
rect 6840 14958 6868 15846
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7024 14618 7052 14758
rect 7116 14618 7144 16623
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7196 15904 7248 15910
rect 7288 15904 7340 15910
rect 7196 15846 7248 15852
rect 7286 15872 7288 15881
rect 7340 15872 7342 15881
rect 7208 15638 7236 15846
rect 7286 15807 7342 15816
rect 7196 15632 7248 15638
rect 7196 15574 7248 15580
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7116 14498 7144 14554
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 7024 14470 7144 14498
rect 6932 13938 6960 14418
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6656 12918 6684 13466
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6380 9438 6500 9466
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 5953 9276 6249 9296
rect 6009 9274 6033 9276
rect 6089 9274 6113 9276
rect 6169 9274 6193 9276
rect 6031 9222 6033 9274
rect 6095 9222 6107 9274
rect 6169 9222 6171 9274
rect 6009 9220 6033 9222
rect 6089 9220 6113 9222
rect 6169 9220 6193 9222
rect 5953 9200 6249 9220
rect 5814 9072 5870 9081
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5540 9036 5592 9042
rect 6380 9042 6408 9318
rect 5814 9007 5870 9016
rect 6368 9036 6420 9042
rect 5540 8978 5592 8984
rect 6368 8978 6420 8984
rect 5552 8090 5580 8978
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 5736 8090 5764 8910
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5460 7002 5488 7822
rect 5828 7546 5856 8910
rect 6196 8566 6224 8910
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 5953 8188 6249 8208
rect 6009 8186 6033 8188
rect 6089 8186 6113 8188
rect 6169 8186 6193 8188
rect 6031 8134 6033 8186
rect 6095 8134 6107 8186
rect 6169 8134 6171 8186
rect 6009 8132 6033 8134
rect 6089 8132 6113 8134
rect 6169 8132 6193 8134
rect 5953 8112 6249 8132
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5632 7336 5684 7342
rect 5630 7304 5632 7313
rect 5684 7304 5686 7313
rect 5630 7239 5686 7248
rect 5644 7206 5672 7239
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5184 5778 5212 6054
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5276 5030 5304 6598
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5460 5710 5488 6122
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5460 5166 5488 5646
rect 5644 5370 5672 6598
rect 5736 5846 5764 6666
rect 5828 6662 5856 7346
rect 5920 7342 5948 7890
rect 6092 7880 6144 7886
rect 6090 7848 6092 7857
rect 6144 7848 6146 7857
rect 6090 7783 6146 7792
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5953 7100 6249 7120
rect 6009 7098 6033 7100
rect 6089 7098 6113 7100
rect 6169 7098 6193 7100
rect 6031 7046 6033 7098
rect 6095 7046 6107 7098
rect 6169 7046 6171 7098
rect 6009 7044 6033 7046
rect 6089 7044 6113 7046
rect 6169 7044 6193 7046
rect 5953 7024 6249 7044
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5920 6458 5948 6802
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 6288 6322 6316 8434
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6380 7886 6408 8366
rect 6472 8276 6500 9438
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6564 8401 6592 8774
rect 6656 8498 6684 12854
rect 6748 12306 6776 13670
rect 6932 13462 6960 13874
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6920 12844 6972 12850
rect 7024 12832 7052 14470
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7116 13734 7144 14350
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 6972 12804 7052 12832
rect 6920 12786 6972 12792
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6840 12374 6868 12582
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6748 11558 6776 11834
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6748 11150 6776 11494
rect 6826 11248 6882 11257
rect 6826 11183 6882 11192
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 10713 6776 11086
rect 6734 10704 6790 10713
rect 6734 10639 6790 10648
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6748 10470 6776 10542
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6748 10198 6776 10406
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6550 8392 6606 8401
rect 6550 8327 6606 8336
rect 6644 8288 6696 8294
rect 6472 8248 6644 8276
rect 6644 8230 6696 8236
rect 6550 7984 6606 7993
rect 6550 7919 6552 7928
rect 6604 7919 6606 7928
rect 6552 7890 6604 7896
rect 6368 7880 6420 7886
rect 6420 7840 6500 7868
rect 6368 7822 6420 7828
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6380 6934 6408 7686
rect 6472 7410 6500 7840
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6564 7721 6592 7754
rect 6550 7712 6606 7721
rect 6550 7647 6606 7656
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6564 7449 6592 7482
rect 6550 7440 6606 7449
rect 6460 7404 6512 7410
rect 6550 7375 6606 7384
rect 6460 7346 6512 7352
rect 6656 7274 6684 8230
rect 6748 8022 6776 9046
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6564 7002 6592 7210
rect 6642 7168 6698 7177
rect 6642 7103 6698 7112
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6550 6896 6606 6905
rect 6550 6831 6606 6840
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 5953 6012 6249 6032
rect 6009 6010 6033 6012
rect 6089 6010 6113 6012
rect 6169 6010 6193 6012
rect 6031 5958 6033 6010
rect 6095 5958 6107 6010
rect 6169 5958 6171 6010
rect 6009 5956 6033 5958
rect 6089 5956 6113 5958
rect 6169 5956 6193 5958
rect 5953 5936 6249 5956
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5736 5370 5764 5782
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 4908 4678 5028 4706
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4712 3528 4764 3534
rect 4816 3505 4844 3878
rect 4712 3470 4764 3476
rect 4802 3496 4858 3505
rect 4724 3398 4752 3470
rect 4802 3431 4858 3440
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4526 3224 4582 3233
rect 4908 3210 4936 4678
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 5000 4146 5028 4490
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4526 3159 4582 3168
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4816 3182 4936 3210
rect 5000 3194 5028 4082
rect 5276 3738 5304 4762
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 4988 3188 5040 3194
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4540 2650 4568 2790
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4436 2576 4488 2582
rect 4436 2518 4488 2524
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3454 2204 3750 2224
rect 3510 2202 3534 2204
rect 3590 2202 3614 2204
rect 3670 2202 3694 2204
rect 3532 2150 3534 2202
rect 3596 2150 3608 2202
rect 3670 2150 3672 2202
rect 3510 2148 3534 2150
rect 3590 2148 3614 2150
rect 3670 2148 3694 2150
rect 3454 2128 3750 2148
rect 3804 1170 3832 2246
rect 3884 2100 3936 2106
rect 3884 2042 3936 2048
rect 3528 1142 3832 1170
rect 3528 800 3556 1142
rect 3896 800 3924 2042
rect 4172 800 4200 2314
rect 4632 1170 4660 2586
rect 4724 2446 4752 3130
rect 4816 3126 4844 3182
rect 4988 3130 5040 3136
rect 4804 3120 4856 3126
rect 4804 3062 4856 3068
rect 4896 3120 4948 3126
rect 4896 3062 4948 3068
rect 4804 2848 4856 2854
rect 4802 2816 4804 2825
rect 4856 2816 4858 2825
rect 4802 2751 4858 2760
rect 4816 2446 4844 2751
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 4540 1142 4660 1170
rect 4540 800 4568 1142
rect 4908 800 4936 3062
rect 5092 3058 5120 3470
rect 5184 3233 5212 3470
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5170 3224 5226 3233
rect 5170 3159 5226 3168
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5172 2508 5224 2514
rect 5276 2496 5304 3334
rect 5368 3194 5396 3878
rect 5460 3534 5488 5102
rect 5953 4924 6249 4944
rect 6009 4922 6033 4924
rect 6089 4922 6113 4924
rect 6169 4922 6193 4924
rect 6031 4870 6033 4922
rect 6095 4870 6107 4922
rect 6169 4870 6171 4922
rect 6009 4868 6033 4870
rect 6089 4868 6113 4870
rect 6169 4868 6193 4870
rect 5953 4848 6249 4868
rect 6288 4826 6316 6258
rect 6380 5370 6408 6598
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5552 4214 5580 4626
rect 6380 4593 6408 5306
rect 6366 4584 6422 4593
rect 6366 4519 6422 4528
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5540 4072 5592 4078
rect 5538 4040 5540 4049
rect 5592 4040 5594 4049
rect 5538 3975 5594 3984
rect 5736 4010 6040 4026
rect 5736 4004 6052 4010
rect 5736 3998 6000 4004
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3652 5580 3878
rect 5552 3624 5672 3652
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5540 3392 5592 3398
rect 5446 3360 5502 3369
rect 5540 3334 5592 3340
rect 5446 3295 5502 3304
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5460 2854 5488 3295
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5224 2468 5304 2496
rect 5172 2450 5224 2456
rect 5264 1556 5316 1562
rect 5264 1498 5316 1504
rect 5276 800 5304 1498
rect 5552 800 5580 3334
rect 5644 2514 5672 3624
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5736 2446 5764 3998
rect 6000 3946 6052 3952
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5828 3738 5856 3878
rect 5953 3836 6249 3856
rect 6009 3834 6033 3836
rect 6089 3834 6113 3836
rect 6169 3834 6193 3836
rect 6031 3782 6033 3834
rect 6095 3782 6107 3834
rect 6169 3782 6171 3834
rect 6009 3780 6033 3782
rect 6089 3780 6113 3782
rect 6169 3780 6193 3782
rect 5953 3760 6249 3780
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5828 2990 5856 3130
rect 6182 3088 6238 3097
rect 6182 3023 6238 3032
rect 6196 2990 6224 3023
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 5828 2514 5856 2926
rect 5953 2748 6249 2768
rect 6009 2746 6033 2748
rect 6089 2746 6113 2748
rect 6169 2746 6193 2748
rect 6031 2694 6033 2746
rect 6095 2694 6107 2746
rect 6169 2694 6171 2746
rect 6009 2692 6033 2694
rect 6089 2692 6113 2694
rect 6169 2692 6193 2694
rect 5953 2672 6249 2692
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6196 1902 6224 2450
rect 6184 1896 6236 1902
rect 6184 1838 6236 1844
rect 6288 1578 6316 4422
rect 6380 4214 6408 4519
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6472 4146 6500 6326
rect 6564 4826 6592 6831
rect 6656 6186 6684 7103
rect 6840 7041 6868 11183
rect 6932 10538 6960 12786
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7024 11626 7052 12174
rect 7116 11898 7144 13670
rect 7208 12322 7236 15574
rect 7288 15564 7340 15570
rect 7392 15552 7420 16050
rect 7340 15524 7420 15552
rect 7288 15506 7340 15512
rect 7392 15026 7420 15524
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7484 14906 7512 17070
rect 7668 16794 7696 19200
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7760 17338 7788 17478
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 8036 17270 8064 19200
rect 8404 17898 8432 19200
rect 8312 17870 8432 17898
rect 8312 17338 8340 17870
rect 8772 17626 8800 19200
rect 8772 17598 8892 17626
rect 8452 17436 8748 17456
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8530 17382 8532 17434
rect 8594 17382 8606 17434
rect 8668 17382 8670 17434
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8452 17360 8748 17380
rect 8864 17338 8892 17598
rect 9140 17338 9168 19200
rect 8300 17332 8352 17338
rect 8852 17332 8904 17338
rect 8300 17274 8352 17280
rect 8404 17292 8708 17320
rect 8024 17264 8076 17270
rect 8024 17206 8076 17212
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7944 16946 7972 17138
rect 8404 17134 8432 17292
rect 8680 17134 8708 17292
rect 8852 17274 8904 17280
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7760 16674 7788 16934
rect 7944 16918 8064 16946
rect 7576 16658 7788 16674
rect 7564 16652 7788 16658
rect 7616 16646 7788 16652
rect 7564 16594 7616 16600
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7760 16250 7788 16526
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7760 15502 7788 15982
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7392 14878 7512 14906
rect 7392 14278 7420 14878
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7484 13870 7512 14758
rect 7656 14476 7708 14482
rect 7760 14464 7788 15438
rect 7932 15428 7984 15434
rect 7932 15370 7984 15376
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7852 15026 7880 15302
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7852 14550 7880 14962
rect 7944 14822 7972 15370
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 8036 14634 8064 16918
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 7944 14606 8064 14634
rect 7840 14544 7892 14550
rect 7840 14486 7892 14492
rect 7708 14436 7788 14464
rect 7656 14418 7708 14424
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7392 13190 7420 13738
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12850 7420 13126
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7378 12744 7434 12753
rect 7378 12679 7380 12688
rect 7432 12679 7434 12688
rect 7380 12650 7432 12656
rect 7392 12442 7420 12650
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7208 12294 7512 12322
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7300 11694 7328 12038
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 7116 10810 7144 11630
rect 7196 11076 7248 11082
rect 7196 11018 7248 11024
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 7208 10470 7236 11018
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7300 10606 7328 10950
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6932 9994 6960 10202
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6932 9081 6960 9930
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6918 9072 6974 9081
rect 6918 9007 6974 9016
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 6932 7954 6960 8502
rect 7024 7993 7052 9862
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7116 8974 7144 9386
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7102 8800 7158 8809
rect 7102 8735 7158 8744
rect 7010 7984 7066 7993
rect 6920 7948 6972 7954
rect 7010 7919 7066 7928
rect 6920 7890 6972 7896
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6826 7032 6882 7041
rect 6932 7002 6960 7346
rect 6826 6967 6882 6976
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7024 6866 7052 7346
rect 7116 7342 7144 8735
rect 7208 8634 7236 10066
rect 7286 9888 7342 9897
rect 7286 9823 7342 9832
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7300 7342 7328 9823
rect 7392 9110 7420 10406
rect 7484 10062 7512 12294
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7484 8294 7512 9998
rect 7576 9926 7604 12242
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7668 11354 7696 11494
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7564 9920 7616 9926
rect 7668 9897 7696 10202
rect 7564 9862 7616 9868
rect 7654 9888 7710 9897
rect 7654 9823 7710 9832
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7472 8288 7524 8294
rect 7564 8288 7616 8294
rect 7472 8230 7524 8236
rect 7562 8256 7564 8265
rect 7616 8256 7618 8265
rect 7562 8191 7618 8200
rect 7576 7732 7604 8191
rect 7668 7834 7696 9318
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7760 8634 7788 8910
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 8129 7788 8230
rect 7746 8120 7802 8129
rect 7746 8055 7802 8064
rect 7668 7806 7788 7834
rect 7656 7744 7708 7750
rect 7576 7704 7656 7732
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 5920 1550 6316 1578
rect 5920 800 5948 1550
rect 6380 1442 6408 4014
rect 6472 3670 6500 4082
rect 6564 3942 6592 4762
rect 6656 4690 6684 6122
rect 6840 5914 6868 6802
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6828 5296 6880 5302
rect 6826 5264 6828 5273
rect 6880 5264 6882 5273
rect 6736 5228 6788 5234
rect 6826 5199 6882 5208
rect 6736 5170 6788 5176
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6748 4146 6776 5170
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6840 4162 6868 5102
rect 6932 5098 6960 5646
rect 7024 5642 7052 6802
rect 7116 6458 7144 7278
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7392 6934 7420 7210
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7116 6254 7144 6394
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7024 4570 7052 4966
rect 7024 4542 7144 4570
rect 6736 4140 6788 4146
rect 6840 4134 7052 4162
rect 6736 4082 6788 4088
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6564 3482 6592 3878
rect 6472 3454 6592 3482
rect 6472 3194 6500 3454
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6458 3088 6514 3097
rect 6458 3023 6460 3032
rect 6512 3023 6514 3032
rect 6460 2994 6512 3000
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 6472 2650 6500 2858
rect 6564 2689 6592 3334
rect 6642 3088 6698 3097
rect 6642 3023 6698 3032
rect 6550 2680 6606 2689
rect 6460 2644 6512 2650
rect 6550 2615 6606 2624
rect 6460 2586 6512 2592
rect 6288 1414 6408 1442
rect 6288 800 6316 1414
rect 6656 800 6684 3023
rect 6748 2990 6776 4082
rect 7024 3534 7052 4134
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6748 2825 6776 2926
rect 6840 2854 6868 3130
rect 6918 2952 6974 2961
rect 7024 2922 7052 3470
rect 6918 2887 6974 2896
rect 7012 2916 7064 2922
rect 6828 2848 6880 2854
rect 6734 2816 6790 2825
rect 6828 2790 6880 2796
rect 6734 2751 6790 2760
rect 6932 2650 6960 2887
rect 7012 2858 7064 2864
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 6932 800 6960 2450
rect 7116 1834 7144 4542
rect 7208 3942 7236 6054
rect 7300 4826 7328 6054
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7392 4826 7420 5714
rect 7484 5710 7512 6258
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7484 5370 7512 5646
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7380 4072 7432 4078
rect 7484 4060 7512 4558
rect 7432 4032 7512 4060
rect 7380 4014 7432 4020
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7208 3346 7236 3538
rect 7300 3466 7328 3878
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7484 3466 7512 3606
rect 7288 3460 7340 3466
rect 7288 3402 7340 3408
rect 7472 3460 7524 3466
rect 7472 3402 7524 3408
rect 7380 3392 7432 3398
rect 7208 3318 7328 3346
rect 7380 3334 7432 3340
rect 7300 2961 7328 3318
rect 7392 2990 7420 3334
rect 7380 2984 7432 2990
rect 7286 2952 7342 2961
rect 7196 2916 7248 2922
rect 7380 2926 7432 2932
rect 7286 2887 7342 2896
rect 7196 2858 7248 2864
rect 7104 1828 7156 1834
rect 7104 1770 7156 1776
rect 7208 1562 7236 2858
rect 7196 1556 7248 1562
rect 7196 1498 7248 1504
rect 7300 800 7328 2887
rect 7576 1902 7604 7704
rect 7656 7686 7708 7692
rect 7760 7342 7788 7806
rect 7748 7336 7800 7342
rect 7668 7296 7748 7324
rect 7668 6662 7696 7296
rect 7748 7278 7800 7284
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7760 6118 7788 7142
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 5574 7788 6054
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 7668 4214 7696 4490
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 7760 4060 7788 5510
rect 7852 4690 7880 11222
rect 7944 8514 7972 14606
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8036 8616 8064 13806
rect 8128 11286 8156 16594
rect 8496 16538 8524 17070
rect 8944 17060 8996 17066
rect 8944 17002 8996 17008
rect 8956 16969 8984 17002
rect 9404 16992 9456 16998
rect 8942 16960 8998 16969
rect 9404 16934 9456 16940
rect 8942 16895 8998 16904
rect 8220 16510 8524 16538
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8220 15638 8248 16510
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8312 16046 8340 16390
rect 8452 16348 8748 16368
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8530 16294 8532 16346
rect 8594 16294 8606 16346
rect 8668 16294 8670 16346
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8452 16272 8748 16292
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8452 15260 8748 15280
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8530 15206 8532 15258
rect 8594 15206 8606 15258
rect 8668 15206 8670 15258
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8452 15184 8748 15204
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8772 14550 8800 14758
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8864 14498 8892 16186
rect 8956 15706 8984 16526
rect 9036 15972 9088 15978
rect 9036 15914 9088 15920
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 15065 8984 15302
rect 8942 15056 8998 15065
rect 9048 15026 9076 15914
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9140 15162 9168 15438
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 8942 14991 8998 15000
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 9048 14618 9076 14962
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 8864 14470 9076 14498
rect 8452 14172 8748 14192
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8530 14118 8532 14170
rect 8594 14118 8606 14170
rect 8668 14118 8670 14170
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8452 14096 8748 14116
rect 8852 14068 8904 14074
rect 8852 14010 8904 14016
rect 8864 13802 8892 14010
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8220 12850 8248 13330
rect 8852 13252 8904 13258
rect 8852 13194 8904 13200
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8312 12782 8340 13126
rect 8452 13084 8748 13104
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8530 13030 8532 13082
rect 8594 13030 8606 13082
rect 8668 13030 8670 13082
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8452 13008 8748 13028
rect 8864 12866 8892 13194
rect 8680 12838 8892 12866
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8390 12472 8446 12481
rect 8680 12442 8708 12838
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8772 12442 8800 12650
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8390 12407 8446 12416
rect 8668 12436 8720 12442
rect 8404 12374 8432 12407
rect 8668 12378 8720 12384
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8392 12368 8444 12374
rect 8298 12336 8354 12345
rect 8208 12300 8260 12306
rect 8392 12310 8444 12316
rect 8298 12271 8354 12280
rect 8208 12242 8260 12248
rect 8220 11830 8248 12242
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 8312 11626 8340 12271
rect 8452 11996 8748 12016
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8530 11942 8532 11994
rect 8594 11942 8606 11994
rect 8668 11942 8670 11994
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8452 11920 8748 11940
rect 8864 11898 8892 12582
rect 8956 12374 8984 13874
rect 9048 12918 9076 14470
rect 9232 13530 9260 15506
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 9126 12880 9182 12889
rect 9126 12815 9182 12824
rect 9140 12714 9168 12815
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8956 11694 8984 12310
rect 9048 12186 9076 12378
rect 9048 12158 9168 12186
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8944 11688 8996 11694
rect 8864 11648 8944 11676
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8116 11280 8168 11286
rect 8300 11280 8352 11286
rect 8116 11222 8168 11228
rect 8298 11248 8300 11257
rect 8352 11248 8354 11257
rect 8298 11183 8354 11192
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8128 9722 8156 9930
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8128 8974 8156 9318
rect 8220 9042 8248 10610
rect 8312 10606 8340 10950
rect 8452 10908 8748 10928
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8530 10854 8532 10906
rect 8594 10854 8606 10906
rect 8668 10854 8670 10906
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8452 10832 8748 10852
rect 8300 10600 8352 10606
rect 8864 10554 8892 11648
rect 8944 11630 8996 11636
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8300 10542 8352 10548
rect 8772 10526 8892 10554
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 9654 8340 10406
rect 8772 10266 8800 10526
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8772 9994 8800 10202
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8452 9820 8748 9840
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8530 9766 8532 9818
rect 8594 9766 8606 9818
rect 8668 9766 8670 9818
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8452 9744 8748 9764
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8772 9466 8800 9590
rect 8864 9586 8892 10406
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8392 9444 8444 9450
rect 8772 9438 8892 9466
rect 8392 9386 8444 9392
rect 8404 9178 8432 9386
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8452 8732 8748 8752
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8530 8678 8532 8730
rect 8594 8678 8606 8730
rect 8668 8678 8670 8730
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8452 8656 8748 8676
rect 8864 8616 8892 9438
rect 8036 8588 8432 8616
rect 7944 8486 8248 8514
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7944 7342 7972 8026
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8128 7002 8156 8366
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8220 6458 8248 8486
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8312 8022 8340 8434
rect 8404 8294 8432 8588
rect 8772 8588 8892 8616
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8666 8528 8722 8537
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8300 8016 8352 8022
rect 8404 7993 8432 8230
rect 8496 8090 8524 8502
rect 8666 8463 8722 8472
rect 8680 8430 8708 8463
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8772 8022 8800 8588
rect 8956 8242 8984 11086
rect 9048 11014 9076 12038
rect 9140 11626 9168 12158
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9232 11286 9260 13466
rect 9416 13326 9444 16934
rect 9508 16810 9536 19200
rect 9508 16782 9628 16810
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9508 15162 9536 16594
rect 9600 15910 9628 16782
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 9692 16590 9720 16662
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9692 16028 9720 16526
rect 9772 16040 9824 16046
rect 9692 16000 9772 16028
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9324 13002 9352 13262
rect 9416 13190 9444 13262
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9324 12974 9444 13002
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 8864 8214 8984 8242
rect 8760 8016 8812 8022
rect 8300 7958 8352 7964
rect 8390 7984 8446 7993
rect 8760 7958 8812 7964
rect 8390 7919 8446 7928
rect 8404 7868 8432 7919
rect 8312 7840 8432 7868
rect 8312 7177 8340 7840
rect 8452 7644 8748 7664
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8530 7590 8532 7642
rect 8594 7590 8606 7642
rect 8668 7590 8670 7642
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8452 7568 8748 7588
rect 8298 7168 8354 7177
rect 8298 7103 8354 7112
rect 8298 7032 8354 7041
rect 8298 6967 8300 6976
rect 8352 6967 8354 6976
rect 8300 6938 8352 6944
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 7932 5840 7984 5846
rect 7932 5782 7984 5788
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7668 4032 7788 4060
rect 7668 3670 7696 4032
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7668 3233 7696 3402
rect 7654 3224 7710 3233
rect 7654 3159 7710 3168
rect 7564 1896 7616 1902
rect 7564 1838 7616 1844
rect 7668 800 7696 3159
rect 7760 2650 7788 3878
rect 7852 3777 7880 4626
rect 7944 4486 7972 5782
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7838 3768 7894 3777
rect 7838 3703 7894 3712
rect 7932 3732 7984 3738
rect 7932 3674 7984 3680
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7852 3398 7880 3470
rect 7840 3392 7892 3398
rect 7944 3369 7972 3674
rect 7840 3334 7892 3340
rect 7930 3360 7986 3369
rect 7852 3058 7880 3334
rect 7930 3295 7986 3304
rect 8036 3194 8064 6394
rect 8312 6390 8340 6938
rect 8452 6556 8748 6576
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8530 6502 8532 6554
rect 8594 6502 8606 6554
rect 8668 6502 8670 6554
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8452 6480 8748 6500
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 8220 5098 8248 5578
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 8312 4826 8340 6054
rect 8772 5914 8800 6326
rect 8760 5908 8812 5914
rect 8864 5896 8892 8214
rect 8942 8120 8998 8129
rect 8942 8055 8944 8064
rect 8996 8055 8998 8064
rect 8944 8026 8996 8032
rect 8942 7984 8998 7993
rect 8942 7919 8944 7928
rect 8996 7919 8998 7928
rect 8944 7890 8996 7896
rect 8944 6248 8996 6254
rect 8942 6216 8944 6225
rect 8996 6216 8998 6225
rect 8942 6151 8998 6160
rect 8864 5868 8984 5896
rect 8760 5850 8812 5856
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8452 5468 8748 5488
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8530 5414 8532 5466
rect 8594 5414 8606 5466
rect 8668 5414 8670 5466
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8452 5392 8748 5412
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8298 4720 8354 4729
rect 8298 4655 8354 4664
rect 8312 4264 8340 4655
rect 8588 4622 8616 4966
rect 8864 4826 8892 5714
rect 8956 5370 8984 5868
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 8452 4380 8748 4400
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8530 4326 8532 4378
rect 8594 4326 8606 4378
rect 8668 4326 8670 4378
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8452 4304 8748 4324
rect 9048 4298 9076 10542
rect 9140 10538 9168 11086
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9140 9926 9168 10474
rect 9232 10441 9260 10950
rect 9218 10432 9274 10441
rect 9218 10367 9274 10376
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9140 9586 9168 9862
rect 9232 9654 9260 10367
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9140 8498 9168 9522
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 9140 6866 9168 7958
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9140 5778 9168 6802
rect 9232 6254 9260 9454
rect 9324 8362 9352 12854
rect 9416 12782 9444 12974
rect 9404 12776 9456 12782
rect 9508 12753 9536 13330
rect 9404 12718 9456 12724
rect 9494 12744 9550 12753
rect 9600 12730 9628 15574
rect 9692 15434 9720 16000
rect 9772 15982 9824 15988
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14618 9720 14758
rect 9784 14618 9812 15030
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9770 14104 9826 14113
rect 9770 14039 9772 14048
rect 9824 14039 9826 14048
rect 9772 14010 9824 14016
rect 9876 13870 9904 19200
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9968 16250 9996 16594
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9968 15502 9996 15914
rect 10060 15570 10088 17478
rect 10140 16788 10192 16794
rect 10140 16730 10192 16736
rect 10152 15910 10180 16730
rect 10244 16726 10272 19200
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10232 16720 10284 16726
rect 10232 16662 10284 16668
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10244 15638 10272 16118
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 10140 15496 10192 15502
rect 10192 15444 10272 15450
rect 10140 15438 10272 15444
rect 9968 15026 9996 15438
rect 10048 15428 10100 15434
rect 10152 15422 10272 15438
rect 10048 15370 10100 15376
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9864 13864 9916 13870
rect 9784 13824 9864 13852
rect 9600 12714 9720 12730
rect 9600 12708 9732 12714
rect 9600 12702 9680 12708
rect 9494 12679 9550 12688
rect 9680 12650 9732 12656
rect 9402 12472 9458 12481
rect 9402 12407 9404 12416
rect 9456 12407 9458 12416
rect 9404 12378 9456 12384
rect 9588 12368 9640 12374
rect 9588 12310 9640 12316
rect 9600 12050 9628 12310
rect 9784 12102 9812 13824
rect 9864 13806 9916 13812
rect 9954 12880 10010 12889
rect 9954 12815 10010 12824
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9876 12374 9904 12650
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9968 12306 9996 12815
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9416 12022 9628 12050
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9416 10198 9444 12022
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9494 11792 9550 11801
rect 9494 11727 9550 11736
rect 9508 11694 9536 11727
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9416 9382 9444 10134
rect 9508 10130 9536 11630
rect 9784 11626 9812 11834
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9586 10976 9642 10985
rect 9642 10934 9720 10962
rect 9586 10911 9642 10920
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9508 9518 9536 10066
rect 9692 10010 9720 10934
rect 9600 9982 9720 10010
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9324 8090 9352 8298
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9416 7886 9444 9318
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9508 8634 9536 9046
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9600 8242 9628 9982
rect 9784 9722 9812 11562
rect 9968 11506 9996 12242
rect 9876 11478 9996 11506
rect 9876 11354 9904 11478
rect 10060 11370 10088 15370
rect 10244 15094 10272 15422
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10152 14074 10180 14894
rect 10336 14482 10364 16934
rect 10612 16640 10640 19200
rect 10980 17105 11008 19200
rect 10966 17096 11022 17105
rect 10966 17031 11022 17040
rect 10950 16892 11246 16912
rect 11006 16890 11030 16892
rect 11086 16890 11110 16892
rect 11166 16890 11190 16892
rect 11028 16838 11030 16890
rect 11092 16838 11104 16890
rect 11166 16838 11168 16890
rect 11006 16836 11030 16838
rect 11086 16836 11110 16838
rect 11166 16836 11190 16838
rect 10950 16816 11246 16836
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 10428 16612 10640 16640
rect 10428 15706 10456 16612
rect 11164 16590 11192 16662
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10336 14226 10364 14418
rect 10428 14346 10456 14758
rect 10416 14340 10468 14346
rect 10416 14282 10468 14288
rect 10336 14198 10456 14226
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10428 13870 10456 14198
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10152 12102 10180 12242
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10152 11762 10180 12038
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9968 11342 10088 11370
rect 9876 10810 9904 11290
rect 9968 11150 9996 11342
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9876 10674 9904 10746
rect 9864 10668 9916 10674
rect 9916 10628 9996 10656
rect 9864 10610 9916 10616
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9508 8214 9628 8242
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9508 7732 9536 8214
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9416 7704 9536 7732
rect 9416 7313 9444 7704
rect 9402 7304 9458 7313
rect 9312 7268 9364 7274
rect 9402 7239 9458 7248
rect 9312 7210 9364 7216
rect 9324 6798 9352 7210
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9140 5574 9168 5714
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 8864 4270 9076 4298
rect 8312 4236 8432 4264
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8128 3194 8156 3878
rect 8220 3670 8248 4082
rect 8300 3936 8352 3942
rect 8404 3913 8432 4236
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8300 3878 8352 3884
rect 8390 3904 8446 3913
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 7852 2446 7880 2994
rect 8036 2938 8064 3130
rect 8220 3126 8248 3606
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8036 2910 8156 2938
rect 8128 2530 8156 2910
rect 8206 2816 8262 2825
rect 8206 2751 8262 2760
rect 8220 2650 8248 2751
rect 8208 2644 8260 2650
rect 8312 2632 8340 3878
rect 8390 3839 8446 3848
rect 8772 3738 8800 4150
rect 8864 3738 8892 4270
rect 9036 4072 9088 4078
rect 9140 4060 9168 5510
rect 9232 4826 9260 6190
rect 9324 5710 9352 6258
rect 9416 5778 9444 7239
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9324 5166 9352 5646
rect 9508 5574 9536 6054
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9088 4032 9168 4060
rect 9036 4014 9088 4020
rect 9232 3942 9260 4762
rect 9324 4622 9352 5102
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9416 4486 9444 5034
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8452 3292 8748 3312
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8530 3238 8532 3290
rect 8594 3238 8606 3290
rect 8668 3238 8670 3290
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8452 3216 8748 3236
rect 8576 3120 8628 3126
rect 8864 3074 8892 3674
rect 8576 3062 8628 3068
rect 8588 2650 8616 3062
rect 8772 3046 8892 3074
rect 8772 2938 8800 3046
rect 8680 2922 8800 2938
rect 8668 2916 8800 2922
rect 8720 2910 8800 2916
rect 8852 2916 8904 2922
rect 8668 2858 8720 2864
rect 8852 2858 8904 2864
rect 8680 2825 8708 2858
rect 8760 2848 8812 2854
rect 8666 2816 8722 2825
rect 8760 2790 8812 2796
rect 8666 2751 8722 2760
rect 8772 2689 8800 2790
rect 8758 2680 8814 2689
rect 8576 2644 8628 2650
rect 8312 2604 8432 2632
rect 8208 2586 8260 2592
rect 8128 2502 8340 2530
rect 8404 2514 8432 2604
rect 8758 2615 8814 2624
rect 8576 2586 8628 2592
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8024 2032 8076 2038
rect 8024 1974 8076 1980
rect 8036 800 8064 1974
rect 8312 800 8340 2502
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 8864 2378 8892 2858
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 8956 2310 8984 3878
rect 9048 3126 9076 3878
rect 9126 3768 9182 3777
rect 9126 3703 9182 3712
rect 9140 3194 9168 3703
rect 9232 3398 9260 3878
rect 9416 3602 9444 4422
rect 9508 3670 9536 5306
rect 9600 4826 9628 8026
rect 9692 6746 9720 9386
rect 9784 9382 9812 9658
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9784 9110 9812 9318
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9876 9042 9904 10406
rect 9968 10130 9996 10628
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9968 8634 9996 9930
rect 10060 9654 10088 11154
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10060 9081 10088 9318
rect 10152 9178 10180 11086
rect 10244 9382 10272 13262
rect 10324 13184 10376 13190
rect 10324 13126 10376 13132
rect 10336 12986 10364 13126
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10322 11792 10378 11801
rect 10322 11727 10324 11736
rect 10376 11727 10378 11736
rect 10324 11698 10376 11704
rect 10428 9738 10456 13806
rect 10520 11898 10548 15846
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10600 15632 10652 15638
rect 10600 15574 10652 15580
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10612 11830 10640 15574
rect 10704 14890 10732 15642
rect 10692 14884 10744 14890
rect 10692 14826 10744 14832
rect 10796 13938 10824 16050
rect 10888 15434 10916 16186
rect 11164 16046 11192 16526
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11348 15858 11376 19200
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11428 16516 11480 16522
rect 11624 16504 11652 16662
rect 11480 16476 11652 16504
rect 11428 16458 11480 16464
rect 11624 16114 11652 16476
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11348 15830 11560 15858
rect 10950 15804 11246 15824
rect 11006 15802 11030 15804
rect 11086 15802 11110 15804
rect 11166 15802 11190 15804
rect 11028 15750 11030 15802
rect 11092 15750 11104 15802
rect 11166 15750 11168 15802
rect 11006 15748 11030 15750
rect 11086 15748 11110 15750
rect 11166 15748 11190 15750
rect 10950 15728 11246 15748
rect 11334 15600 11390 15609
rect 11334 15535 11336 15544
rect 11388 15535 11390 15544
rect 11336 15506 11388 15512
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10980 15314 11008 15438
rect 10888 15286 11008 15314
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10888 13818 10916 15286
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 10950 14716 11246 14736
rect 11006 14714 11030 14716
rect 11086 14714 11110 14716
rect 11166 14714 11190 14716
rect 11028 14662 11030 14714
rect 11092 14662 11104 14714
rect 11166 14662 11168 14714
rect 11006 14660 11030 14662
rect 11086 14660 11110 14662
rect 11166 14660 11190 14662
rect 10950 14640 11246 14660
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11164 14074 11192 14418
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 10704 13790 10916 13818
rect 11072 13802 11100 13942
rect 11348 13870 11376 15030
rect 11440 15026 11468 15302
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11336 13864 11388 13870
rect 11336 13806 11388 13812
rect 11060 13796 11112 13802
rect 10704 12458 10732 13790
rect 11060 13738 11112 13744
rect 10950 13628 11246 13648
rect 11006 13626 11030 13628
rect 11086 13626 11110 13628
rect 11166 13626 11190 13628
rect 11028 13574 11030 13626
rect 11092 13574 11104 13626
rect 11166 13574 11168 13626
rect 11006 13572 11030 13574
rect 11086 13572 11110 13574
rect 11166 13572 11190 13574
rect 10950 13552 11246 13572
rect 11440 13530 11468 14554
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10796 12986 10824 13262
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10888 12646 10916 13262
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10950 12540 11246 12560
rect 11006 12538 11030 12540
rect 11086 12538 11110 12540
rect 11166 12538 11190 12540
rect 11028 12486 11030 12538
rect 11092 12486 11104 12538
rect 11166 12486 11168 12538
rect 11006 12484 11030 12486
rect 11086 12484 11110 12486
rect 11166 12484 11190 12486
rect 10950 12464 11246 12484
rect 10704 12430 10916 12458
rect 11348 12442 11376 13330
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10796 10606 10824 11086
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10428 9710 10640 9738
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10046 9072 10102 9081
rect 10046 9007 10102 9016
rect 10140 9036 10192 9042
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9784 8022 9812 8502
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 10060 8242 10088 9007
rect 10140 8978 10192 8984
rect 10152 8838 10180 8978
rect 10244 8945 10272 9318
rect 10336 9178 10364 9522
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10416 8968 10468 8974
rect 10230 8936 10286 8945
rect 10416 8910 10468 8916
rect 10230 8871 10286 8880
rect 10140 8832 10192 8838
rect 10140 8774 10192 8780
rect 10152 8498 10180 8774
rect 10428 8673 10456 8910
rect 10414 8664 10470 8673
rect 10520 8634 10548 9318
rect 10414 8599 10470 8608
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10336 8294 10364 8366
rect 10324 8288 10376 8294
rect 9968 8090 9996 8230
rect 10060 8214 10272 8242
rect 10324 8230 10376 8236
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 9956 8084 10008 8090
rect 10008 8044 10088 8072
rect 9956 8026 10008 8032
rect 9772 8016 9824 8022
rect 9772 7958 9824 7964
rect 9784 7342 9812 7958
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9784 6866 9812 7278
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9876 6866 9904 7142
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9692 6718 9812 6746
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6322 9720 6598
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9692 5273 9720 5306
rect 9678 5264 9734 5273
rect 9678 5199 9734 5208
rect 9588 4820 9640 4826
rect 9640 4780 9720 4808
rect 9588 4762 9640 4768
rect 9588 4616 9640 4622
rect 9586 4584 9588 4593
rect 9640 4584 9642 4593
rect 9586 4519 9642 4528
rect 9586 4176 9642 4185
rect 9586 4111 9642 4120
rect 9496 3664 9548 3670
rect 9496 3606 9548 3612
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 9034 2544 9090 2553
rect 9034 2479 9090 2488
rect 9140 2496 9168 3130
rect 9416 3058 9444 3538
rect 9600 3534 9628 4111
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9508 2922 9536 3334
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9600 2650 9628 3470
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9220 2508 9272 2514
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8452 2204 8748 2224
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8530 2150 8532 2202
rect 8594 2150 8606 2202
rect 8668 2150 8670 2202
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8452 2128 8748 2148
rect 8668 1828 8720 1834
rect 8668 1770 8720 1776
rect 8680 800 8708 1770
rect 9048 800 9076 2479
rect 9140 2468 9220 2496
rect 9220 2450 9272 2456
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9140 2106 9168 2246
rect 9128 2100 9180 2106
rect 9128 2042 9180 2048
rect 9508 2038 9536 2450
rect 9496 2032 9548 2038
rect 9496 1974 9548 1980
rect 9312 1760 9364 1766
rect 9312 1702 9364 1708
rect 9324 800 9352 1702
rect 9692 800 9720 4780
rect 9784 3602 9812 6718
rect 9876 6322 9904 6802
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9876 4060 9904 5714
rect 9968 4690 9996 6598
rect 10060 5914 10088 8044
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10152 7478 10180 7754
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10140 6928 10192 6934
rect 10140 6870 10192 6876
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10060 5166 10088 5714
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10152 5012 10180 6870
rect 10244 6474 10272 8214
rect 10428 7993 10456 8230
rect 10414 7984 10470 7993
rect 10414 7919 10470 7928
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10336 7546 10364 7686
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10520 6662 10548 8366
rect 10612 8362 10640 9710
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10704 9110 10732 9522
rect 10782 9480 10838 9489
rect 10782 9415 10838 9424
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10704 8974 10732 9046
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10796 8090 10824 9415
rect 10888 9160 10916 12430
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11440 12170 11468 12786
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 10950 11452 11246 11472
rect 11006 11450 11030 11452
rect 11086 11450 11110 11452
rect 11166 11450 11190 11452
rect 11028 11398 11030 11450
rect 11092 11398 11104 11450
rect 11166 11398 11168 11450
rect 11006 11396 11030 11398
rect 11086 11396 11110 11398
rect 11166 11396 11190 11398
rect 10950 11376 11246 11396
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11072 10674 11100 11018
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10950 10364 11246 10384
rect 11006 10362 11030 10364
rect 11086 10362 11110 10364
rect 11166 10362 11190 10364
rect 11028 10310 11030 10362
rect 11092 10310 11104 10362
rect 11166 10310 11168 10362
rect 11006 10308 11030 10310
rect 11086 10308 11110 10310
rect 11166 10308 11190 10310
rect 10950 10288 11246 10308
rect 11348 10198 11376 10678
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11440 9625 11468 10406
rect 11426 9616 11482 9625
rect 11426 9551 11482 9560
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11428 9444 11480 9450
rect 11428 9386 11480 9392
rect 10950 9276 11246 9296
rect 11006 9274 11030 9276
rect 11086 9274 11110 9276
rect 11166 9274 11190 9276
rect 11028 9222 11030 9274
rect 11092 9222 11104 9274
rect 11166 9222 11168 9274
rect 11006 9220 11030 9222
rect 11086 9220 11110 9222
rect 11166 9220 11190 9222
rect 10950 9200 11246 9220
rect 10888 9132 11008 9160
rect 10980 8276 11008 9132
rect 11348 9081 11376 9386
rect 11334 9072 11390 9081
rect 11244 9036 11296 9042
rect 11334 9007 11390 9016
rect 11244 8978 11296 8984
rect 11256 8566 11284 8978
rect 11440 8945 11468 9386
rect 11426 8936 11482 8945
rect 11336 8900 11388 8906
rect 11426 8871 11482 8880
rect 11336 8842 11388 8848
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 10888 8248 11008 8276
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10692 7948 10744 7954
rect 10692 7890 10744 7896
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10612 7342 10640 7822
rect 10704 7546 10732 7890
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10244 6446 10548 6474
rect 10322 6216 10378 6225
rect 10322 6151 10378 6160
rect 10336 5846 10364 6151
rect 10324 5840 10376 5846
rect 10060 4984 10180 5012
rect 10244 5800 10324 5828
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9956 4072 10008 4078
rect 9876 4032 9956 4060
rect 9956 4014 10008 4020
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9770 2952 9826 2961
rect 9770 2887 9772 2896
rect 9824 2887 9826 2896
rect 9772 2858 9824 2864
rect 9876 2514 9904 3334
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9968 2650 9996 2926
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 10060 800 10088 4984
rect 10140 4752 10192 4758
rect 10140 4694 10192 4700
rect 10152 3738 10180 4694
rect 10244 4214 10272 5800
rect 10324 5782 10376 5788
rect 10324 5092 10376 5098
rect 10324 5034 10376 5040
rect 10336 4758 10364 5034
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10414 4720 10470 4729
rect 10414 4655 10470 4664
rect 10428 4622 10456 4655
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10140 3732 10192 3738
rect 10192 3692 10272 3720
rect 10140 3674 10192 3680
rect 10244 2854 10272 3692
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10336 1834 10364 4490
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10428 4146 10456 4422
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10520 3942 10548 6446
rect 10612 6254 10640 7142
rect 10704 6934 10732 7210
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10704 6100 10732 6870
rect 10796 6458 10824 7822
rect 10888 7274 10916 8248
rect 10950 8188 11246 8208
rect 11006 8186 11030 8188
rect 11086 8186 11110 8188
rect 11166 8186 11190 8188
rect 11028 8134 11030 8186
rect 11092 8134 11104 8186
rect 11166 8134 11168 8186
rect 11006 8132 11030 8134
rect 11086 8132 11110 8134
rect 11166 8132 11190 8134
rect 10950 8112 11246 8132
rect 11348 8090 11376 8842
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11440 8090 11468 8434
rect 11532 8129 11560 15830
rect 11624 15502 11652 16050
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11624 14550 11652 14962
rect 11716 14804 11744 16934
rect 11808 15638 11836 19200
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11796 15496 11848 15502
rect 11794 15464 11796 15473
rect 11848 15464 11850 15473
rect 11794 15399 11850 15408
rect 11796 14816 11848 14822
rect 11716 14776 11796 14804
rect 11796 14758 11848 14764
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11624 13530 11652 13942
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11808 12646 11836 14758
rect 11900 14482 11928 15982
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11612 12232 11664 12238
rect 11664 12180 11744 12186
rect 11612 12174 11744 12180
rect 11624 12158 11744 12174
rect 11716 12102 11744 12158
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11610 11792 11666 11801
rect 11610 11727 11666 11736
rect 11624 9722 11652 11727
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11624 9518 11652 9658
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11518 8120 11574 8129
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11428 8084 11480 8090
rect 11518 8055 11574 8064
rect 11428 8026 11480 8032
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11348 7410 11376 7890
rect 11624 7868 11652 9454
rect 11615 7857 11652 7868
rect 11610 7848 11666 7857
rect 11610 7783 11666 7792
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 10950 7100 11246 7120
rect 11006 7098 11030 7100
rect 11086 7098 11110 7100
rect 11166 7098 11190 7100
rect 11028 7046 11030 7098
rect 11092 7046 11104 7098
rect 11166 7046 11168 7098
rect 11006 7044 11030 7046
rect 11086 7044 11110 7046
rect 11166 7044 11190 7046
rect 10950 7024 11246 7044
rect 11348 6984 11376 7346
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11440 7002 11468 7278
rect 11164 6956 11376 6984
rect 11428 6996 11480 7002
rect 11164 6662 11192 6956
rect 11428 6938 11480 6944
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 11164 6322 11192 6598
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 10612 6072 10732 6100
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10414 3496 10470 3505
rect 10612 3482 10640 6072
rect 10950 6012 11246 6032
rect 11006 6010 11030 6012
rect 11086 6010 11110 6012
rect 11166 6010 11190 6012
rect 11028 5958 11030 6010
rect 11092 5958 11104 6010
rect 11166 5958 11168 6010
rect 11006 5956 11030 5958
rect 11086 5956 11110 5958
rect 11166 5956 11190 5958
rect 10950 5936 11246 5956
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10704 5030 10732 5782
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10704 4214 10732 4966
rect 10950 4924 11246 4944
rect 11006 4922 11030 4924
rect 11086 4922 11110 4924
rect 11166 4922 11190 4924
rect 11028 4870 11030 4922
rect 11092 4870 11104 4922
rect 11166 4870 11168 4922
rect 11006 4868 11030 4870
rect 11086 4868 11110 4870
rect 11166 4868 11190 4870
rect 10950 4848 11246 4868
rect 11348 4690 11376 5102
rect 11440 4826 11468 6938
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 10796 4282 10824 4626
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10782 3904 10838 3913
rect 10470 3454 10640 3482
rect 10414 3431 10470 3440
rect 10324 1828 10376 1834
rect 10324 1770 10376 1776
rect 10428 800 10456 3431
rect 10704 2106 10732 3878
rect 10782 3839 10838 3848
rect 10796 2553 10824 3839
rect 10888 3738 10916 4558
rect 10950 3836 11246 3856
rect 11006 3834 11030 3836
rect 11086 3834 11110 3836
rect 11166 3834 11190 3836
rect 11028 3782 11030 3834
rect 11092 3782 11104 3834
rect 11166 3782 11168 3834
rect 11006 3780 11030 3782
rect 11086 3780 11110 3782
rect 11166 3780 11190 3782
rect 10950 3760 11246 3780
rect 11348 3738 11376 4626
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 10888 2632 10916 3538
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10980 3194 11008 3470
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10950 2748 11246 2768
rect 11006 2746 11030 2748
rect 11086 2746 11110 2748
rect 11166 2746 11190 2748
rect 11028 2694 11030 2746
rect 11092 2694 11104 2746
rect 11166 2694 11168 2746
rect 11006 2692 11030 2694
rect 11086 2692 11110 2694
rect 11166 2692 11190 2694
rect 10950 2672 11246 2692
rect 11348 2650 11376 3538
rect 11440 3534 11468 4082
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11532 3194 11560 3878
rect 11624 3738 11652 7783
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11624 3058 11652 3538
rect 11716 3398 11744 12038
rect 11808 9761 11836 12582
rect 11794 9752 11850 9761
rect 11794 9687 11850 9696
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11808 6934 11836 8366
rect 11900 7342 11928 14418
rect 11992 13682 12020 17614
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 12084 14346 12112 16594
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 12084 13870 12112 14282
rect 12176 14113 12204 19200
rect 12256 16176 12308 16182
rect 12256 16118 12308 16124
rect 12268 15502 12296 16118
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12268 14278 12296 14962
rect 12348 14884 12400 14890
rect 12348 14826 12400 14832
rect 12360 14618 12388 14826
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12162 14104 12218 14113
rect 12268 14074 12296 14214
rect 12162 14039 12218 14048
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12268 13938 12296 14010
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 11992 13654 12204 13682
rect 11980 10192 12032 10198
rect 11980 10134 12032 10140
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11900 7002 11928 7142
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11336 2644 11388 2650
rect 10888 2604 11100 2632
rect 10782 2544 10838 2553
rect 10782 2479 10838 2488
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 10796 1970 10824 2246
rect 10784 1964 10836 1970
rect 10784 1906 10836 1912
rect 10690 912 10746 921
rect 10690 847 10746 856
rect 10704 800 10732 847
rect 11072 800 11100 2604
rect 11336 2586 11388 2592
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11256 2310 11284 2382
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11256 2106 11284 2246
rect 11244 2100 11296 2106
rect 11244 2042 11296 2048
rect 11440 800 11468 2586
rect 11624 2446 11652 2994
rect 11808 2514 11836 3674
rect 11992 2582 12020 10134
rect 12072 9512 12124 9518
rect 12070 9480 12072 9489
rect 12124 9480 12126 9489
rect 12070 9415 12126 9424
rect 12176 8634 12204 13654
rect 12452 13462 12480 14758
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12452 10198 12480 12922
rect 12440 10192 12492 10198
rect 12440 10134 12492 10140
rect 12544 10146 12572 19200
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12636 13734 12664 15846
rect 12820 15706 12848 15846
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12912 15094 12940 19200
rect 13280 16776 13308 19200
rect 13648 17898 13676 19200
rect 14016 17898 14044 19200
rect 13188 16748 13308 16776
rect 13372 17870 13676 17898
rect 13832 17870 14044 17898
rect 12992 16516 13044 16522
rect 12992 16458 13044 16464
rect 13004 16114 13032 16458
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12900 15088 12952 15094
rect 12900 15030 12952 15036
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12820 14618 12848 14758
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12900 14544 12952 14550
rect 12900 14486 12952 14492
rect 12716 14476 12768 14482
rect 12768 14436 12848 14464
rect 12716 14418 12768 14424
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12728 12442 12756 14282
rect 12820 14278 12848 14436
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12728 12102 12756 12378
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10674 12756 10950
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12820 10554 12848 14214
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12728 10526 12848 10554
rect 12636 10266 12664 10474
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12544 10118 12664 10146
rect 12636 9874 12664 10118
rect 12452 9846 12664 9874
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12084 7993 12112 8366
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12070 7984 12126 7993
rect 12070 7919 12126 7928
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 12084 6866 12112 7278
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12084 6662 12112 6802
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 12084 5370 12112 6598
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 12084 3942 12112 4014
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12084 2650 12112 3878
rect 12176 2922 12204 8026
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 11980 2576 12032 2582
rect 11980 2518 12032 2524
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 12070 2408 12126 2417
rect 12070 2343 12126 2352
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 11716 1306 11744 1974
rect 11992 1902 12020 2246
rect 11980 1896 12032 1902
rect 11980 1838 12032 1844
rect 11716 1278 11836 1306
rect 11808 800 11836 1278
rect 12084 800 12112 2343
rect 12176 1766 12204 2858
rect 12268 2854 12296 9114
rect 12348 8560 12400 8566
rect 12346 8528 12348 8537
rect 12400 8528 12402 8537
rect 12346 8463 12402 8472
rect 12452 8294 12480 9846
rect 12728 9738 12756 10526
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12820 10266 12848 10406
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12808 9988 12860 9994
rect 12808 9930 12860 9936
rect 12636 9710 12756 9738
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12440 7268 12492 7274
rect 12440 7210 12492 7216
rect 12452 7002 12480 7210
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12544 6882 12572 9114
rect 12452 6854 12572 6882
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12360 4690 12388 5170
rect 12452 5166 12480 6854
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12360 4146 12388 4626
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12360 3738 12388 4082
rect 12544 4049 12572 6734
rect 12636 5114 12664 9710
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12728 9042 12756 9522
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12728 8498 12756 8978
rect 12820 8922 12848 9930
rect 12912 9178 12940 14486
rect 13004 14482 13032 16050
rect 13188 15570 13216 16748
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 13004 10062 13032 11154
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13004 9178 13032 9998
rect 13096 9518 13124 15030
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12820 8894 13124 8922
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 12806 8664 12862 8673
rect 12806 8599 12862 8608
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12728 8090 12756 8434
rect 12820 8430 12848 8599
rect 13004 8498 13032 8774
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12808 8288 12860 8294
rect 12860 8248 13032 8276
rect 12808 8230 12860 8236
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12820 6322 12848 6802
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12900 5160 12952 5166
rect 12636 5086 12756 5114
rect 12900 5102 12952 5108
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12530 4040 12586 4049
rect 12636 4010 12664 4966
rect 12728 4826 12756 5086
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12808 4752 12860 4758
rect 12806 4720 12808 4729
rect 12860 4720 12862 4729
rect 12716 4684 12768 4690
rect 12806 4655 12862 4664
rect 12716 4626 12768 4632
rect 12728 4486 12756 4626
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12728 4214 12756 4422
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 12820 4146 12848 4422
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12530 3975 12586 3984
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12452 2650 12480 2790
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12452 2378 12480 2586
rect 12440 2372 12492 2378
rect 12440 2314 12492 2320
rect 12440 1828 12492 1834
rect 12440 1770 12492 1776
rect 12164 1760 12216 1766
rect 12164 1702 12216 1708
rect 12452 800 12480 1770
rect 12636 1714 12664 3606
rect 12806 3088 12862 3097
rect 12806 3023 12862 3032
rect 12820 2650 12848 3023
rect 12912 2650 12940 5102
rect 13004 2854 13032 8248
rect 13096 3670 13124 8894
rect 13188 8362 13216 15098
rect 13280 14278 13308 16594
rect 13372 16046 13400 17870
rect 13449 17436 13745 17456
rect 13505 17434 13529 17436
rect 13585 17434 13609 17436
rect 13665 17434 13689 17436
rect 13527 17382 13529 17434
rect 13591 17382 13603 17434
rect 13665 17382 13667 17434
rect 13505 17380 13529 17382
rect 13585 17380 13609 17382
rect 13665 17380 13689 17382
rect 13449 17360 13745 17380
rect 13449 16348 13745 16368
rect 13505 16346 13529 16348
rect 13585 16346 13609 16348
rect 13665 16346 13689 16348
rect 13527 16294 13529 16346
rect 13591 16294 13603 16346
rect 13665 16294 13667 16346
rect 13505 16292 13529 16294
rect 13585 16292 13609 16294
rect 13665 16292 13689 16294
rect 13449 16272 13745 16292
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13449 15260 13745 15280
rect 13505 15258 13529 15260
rect 13585 15258 13609 15260
rect 13665 15258 13689 15260
rect 13527 15206 13529 15258
rect 13591 15206 13603 15258
rect 13665 15206 13667 15258
rect 13505 15204 13529 15206
rect 13585 15204 13609 15206
rect 13665 15204 13689 15206
rect 13449 15184 13745 15204
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 14618 13584 14758
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13449 14172 13745 14192
rect 13505 14170 13529 14172
rect 13585 14170 13609 14172
rect 13665 14170 13689 14172
rect 13527 14118 13529 14170
rect 13591 14118 13603 14170
rect 13665 14118 13667 14170
rect 13505 14116 13529 14118
rect 13585 14116 13609 14118
rect 13665 14116 13689 14118
rect 13449 14096 13745 14116
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13280 13326 13308 13670
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13176 6928 13228 6934
rect 13176 6870 13228 6876
rect 13188 6662 13216 6870
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12900 2644 12952 2650
rect 12900 2586 12952 2592
rect 12636 1686 12848 1714
rect 12820 800 12848 1686
rect 13188 800 13216 6598
rect 13280 3641 13308 13262
rect 13449 13084 13745 13104
rect 13505 13082 13529 13084
rect 13585 13082 13609 13084
rect 13665 13082 13689 13084
rect 13527 13030 13529 13082
rect 13591 13030 13603 13082
rect 13665 13030 13667 13082
rect 13505 13028 13529 13030
rect 13585 13028 13609 13030
rect 13665 13028 13689 13030
rect 13449 13008 13745 13028
rect 13832 12986 13860 17870
rect 14384 17762 14412 19200
rect 13924 17734 14412 17762
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13449 11996 13745 12016
rect 13505 11994 13529 11996
rect 13585 11994 13609 11996
rect 13665 11994 13689 11996
rect 13527 11942 13529 11994
rect 13591 11942 13603 11994
rect 13665 11942 13667 11994
rect 13505 11940 13529 11942
rect 13585 11940 13609 11942
rect 13665 11940 13689 11942
rect 13449 11920 13745 11940
rect 13449 10908 13745 10928
rect 13505 10906 13529 10908
rect 13585 10906 13609 10908
rect 13665 10906 13689 10908
rect 13527 10854 13529 10906
rect 13591 10854 13603 10906
rect 13665 10854 13667 10906
rect 13505 10852 13529 10854
rect 13585 10852 13609 10854
rect 13665 10852 13689 10854
rect 13449 10832 13745 10852
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13372 10266 13400 10406
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13449 9820 13745 9840
rect 13505 9818 13529 9820
rect 13585 9818 13609 9820
rect 13665 9818 13689 9820
rect 13527 9766 13529 9818
rect 13591 9766 13603 9818
rect 13665 9766 13667 9818
rect 13505 9764 13529 9766
rect 13585 9764 13609 9766
rect 13665 9764 13689 9766
rect 13449 9744 13745 9764
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13449 8732 13745 8752
rect 13505 8730 13529 8732
rect 13585 8730 13609 8732
rect 13665 8730 13689 8732
rect 13527 8678 13529 8730
rect 13591 8678 13603 8730
rect 13665 8678 13667 8730
rect 13505 8676 13529 8678
rect 13585 8676 13609 8678
rect 13665 8676 13689 8678
rect 13449 8656 13745 8676
rect 13360 8356 13412 8362
rect 13360 8298 13412 8304
rect 13372 6866 13400 8298
rect 13449 7644 13745 7664
rect 13505 7642 13529 7644
rect 13585 7642 13609 7644
rect 13665 7642 13689 7644
rect 13527 7590 13529 7642
rect 13591 7590 13603 7642
rect 13665 7590 13667 7642
rect 13505 7588 13529 7590
rect 13585 7588 13609 7590
rect 13665 7588 13689 7590
rect 13449 7568 13745 7588
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13449 6556 13745 6576
rect 13505 6554 13529 6556
rect 13585 6554 13609 6556
rect 13665 6554 13689 6556
rect 13527 6502 13529 6554
rect 13591 6502 13603 6554
rect 13665 6502 13667 6554
rect 13505 6500 13529 6502
rect 13585 6500 13609 6502
rect 13665 6500 13689 6502
rect 13449 6480 13745 6500
rect 13449 5468 13745 5488
rect 13505 5466 13529 5468
rect 13585 5466 13609 5468
rect 13665 5466 13689 5468
rect 13527 5414 13529 5466
rect 13591 5414 13603 5466
rect 13665 5414 13667 5466
rect 13505 5412 13529 5414
rect 13585 5412 13609 5414
rect 13665 5412 13689 5414
rect 13449 5392 13745 5412
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13372 4622 13400 5170
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13464 4554 13492 4762
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13266 3632 13322 3641
rect 13266 3567 13322 3576
rect 13372 3482 13400 4422
rect 13449 4380 13745 4400
rect 13505 4378 13529 4380
rect 13585 4378 13609 4380
rect 13665 4378 13689 4380
rect 13527 4326 13529 4378
rect 13591 4326 13603 4378
rect 13665 4326 13667 4378
rect 13505 4324 13529 4326
rect 13585 4324 13609 4326
rect 13665 4324 13689 4326
rect 13449 4304 13745 4324
rect 13280 3454 13400 3482
rect 13280 1986 13308 3454
rect 13449 3292 13745 3312
rect 13505 3290 13529 3292
rect 13585 3290 13609 3292
rect 13665 3290 13689 3292
rect 13527 3238 13529 3290
rect 13591 3238 13603 3290
rect 13665 3238 13667 3290
rect 13505 3236 13529 3238
rect 13585 3236 13609 3238
rect 13665 3236 13689 3238
rect 13449 3216 13745 3236
rect 13449 2204 13745 2224
rect 13505 2202 13529 2204
rect 13585 2202 13609 2204
rect 13665 2202 13689 2204
rect 13527 2150 13529 2202
rect 13591 2150 13603 2202
rect 13665 2150 13667 2202
rect 13505 2148 13529 2150
rect 13585 2148 13609 2150
rect 13665 2148 13689 2150
rect 13449 2128 13745 2148
rect 13280 1958 13492 1986
rect 13464 800 13492 1958
rect 13832 800 13860 9318
rect 13924 8430 13952 17734
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 14108 2650 14136 16594
rect 14292 2990 14320 17070
rect 14660 16658 14688 17546
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 14370 16008 14426 16017
rect 14370 15943 14426 15952
rect 14384 15638 14412 15943
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 14752 4826 14780 19200
rect 15016 17740 15068 17746
rect 15016 17682 15068 17688
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14844 16561 14872 17002
rect 14830 16552 14886 16561
rect 14830 16487 14886 16496
rect 14924 15360 14976 15366
rect 14924 15302 14976 15308
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 14844 5370 14872 7414
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14844 5166 14872 5306
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14936 4706 14964 15302
rect 15028 9518 15056 17682
rect 15120 16250 15148 19200
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15488 14346 15516 19200
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15856 13394 15884 19200
rect 16224 13802 16252 19200
rect 16592 15162 16620 19200
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16960 14550 16988 19200
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 16224 10266 16252 13738
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 15290 10024 15346 10033
rect 15290 9959 15346 9968
rect 15304 9586 15332 9959
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 14568 4678 14964 4706
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14568 2972 14596 4678
rect 14648 2984 14700 2990
rect 14568 2944 14648 2972
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 14108 2514 14136 2586
rect 14186 2544 14242 2553
rect 14096 2508 14148 2514
rect 14186 2479 14242 2488
rect 14096 2450 14148 2456
rect 14200 800 14228 2479
rect 14568 800 14596 2944
rect 14648 2926 14700 2932
rect 15936 2916 15988 2922
rect 15936 2858 15988 2864
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 14646 2544 14702 2553
rect 14646 2479 14648 2488
rect 14700 2479 14702 2488
rect 14648 2450 14700 2456
rect 14844 800 14872 2586
rect 15212 800 15240 2790
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15580 800 15608 2382
rect 15948 800 15976 2858
rect 16224 800 16252 5034
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 16592 800 16620 2518
rect 16960 800 16988 2994
rect 1490 504 1546 513
rect 1490 439 1546 448
rect 1766 0 1822 800
rect 2134 0 2190 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
<< via2 >>
rect 1950 19352 2006 19408
rect 1674 18400 1730 18456
rect 570 15952 626 16008
rect 1766 16496 1822 16552
rect 1766 16360 1822 16416
rect 1674 15444 1676 15464
rect 1676 15444 1728 15464
rect 1728 15444 1730 15464
rect 1674 15408 1730 15444
rect 1674 14356 1676 14376
rect 1676 14356 1728 14376
rect 1728 14356 1730 14376
rect 1674 14320 1730 14356
rect 1858 13368 1914 13424
rect 1766 12416 1822 12472
rect 1766 11328 1822 11384
rect 1490 9560 1546 9616
rect 1766 8336 1822 8392
rect 1674 7404 1730 7440
rect 1674 7384 1676 7404
rect 1676 7384 1728 7404
rect 1728 7384 1730 7404
rect 1674 6432 1730 6488
rect 2226 5344 2282 5400
rect 3454 17434 3510 17436
rect 3534 17434 3590 17436
rect 3614 17434 3670 17436
rect 3694 17434 3750 17436
rect 3454 17382 3480 17434
rect 3480 17382 3510 17434
rect 3534 17382 3544 17434
rect 3544 17382 3590 17434
rect 3614 17382 3660 17434
rect 3660 17382 3670 17434
rect 3694 17382 3724 17434
rect 3724 17382 3750 17434
rect 3454 17380 3510 17382
rect 3534 17380 3590 17382
rect 3614 17380 3670 17382
rect 3694 17380 3750 17382
rect 3422 16652 3478 16688
rect 3422 16632 3424 16652
rect 3424 16632 3476 16652
rect 3476 16632 3478 16652
rect 3454 16346 3510 16348
rect 3534 16346 3590 16348
rect 3614 16346 3670 16348
rect 3694 16346 3750 16348
rect 3454 16294 3480 16346
rect 3480 16294 3510 16346
rect 3534 16294 3544 16346
rect 3544 16294 3590 16346
rect 3614 16294 3660 16346
rect 3660 16294 3670 16346
rect 3694 16294 3724 16346
rect 3724 16294 3750 16346
rect 3454 16292 3510 16294
rect 3534 16292 3590 16294
rect 3614 16292 3670 16294
rect 3694 16292 3750 16294
rect 3454 15258 3510 15260
rect 3534 15258 3590 15260
rect 3614 15258 3670 15260
rect 3694 15258 3750 15260
rect 3454 15206 3480 15258
rect 3480 15206 3510 15258
rect 3534 15206 3544 15258
rect 3544 15206 3590 15258
rect 3614 15206 3660 15258
rect 3660 15206 3670 15258
rect 3694 15206 3724 15258
rect 3724 15206 3750 15258
rect 3454 15204 3510 15206
rect 3534 15204 3590 15206
rect 3614 15204 3670 15206
rect 3694 15204 3750 15206
rect 3974 16632 4030 16688
rect 3454 14170 3510 14172
rect 3534 14170 3590 14172
rect 3614 14170 3670 14172
rect 3694 14170 3750 14172
rect 3454 14118 3480 14170
rect 3480 14118 3510 14170
rect 3534 14118 3544 14170
rect 3544 14118 3590 14170
rect 3614 14118 3660 14170
rect 3660 14118 3670 14170
rect 3694 14118 3724 14170
rect 3724 14118 3750 14170
rect 3454 14116 3510 14118
rect 3534 14116 3590 14118
rect 3614 14116 3670 14118
rect 3694 14116 3750 14118
rect 3454 13082 3510 13084
rect 3534 13082 3590 13084
rect 3614 13082 3670 13084
rect 3694 13082 3750 13084
rect 3454 13030 3480 13082
rect 3480 13030 3510 13082
rect 3534 13030 3544 13082
rect 3544 13030 3590 13082
rect 3614 13030 3660 13082
rect 3660 13030 3670 13082
rect 3694 13030 3724 13082
rect 3724 13030 3750 13082
rect 3454 13028 3510 13030
rect 3534 13028 3590 13030
rect 3614 13028 3670 13030
rect 3694 13028 3750 13030
rect 3454 11994 3510 11996
rect 3534 11994 3590 11996
rect 3614 11994 3670 11996
rect 3694 11994 3750 11996
rect 3454 11942 3480 11994
rect 3480 11942 3510 11994
rect 3534 11942 3544 11994
rect 3544 11942 3590 11994
rect 3614 11942 3660 11994
rect 3660 11942 3670 11994
rect 3694 11942 3724 11994
rect 3724 11942 3750 11994
rect 3454 11940 3510 11942
rect 3534 11940 3590 11942
rect 3614 11940 3670 11942
rect 3694 11940 3750 11942
rect 2778 10376 2834 10432
rect 3454 10906 3510 10908
rect 3534 10906 3590 10908
rect 3614 10906 3670 10908
rect 3694 10906 3750 10908
rect 3454 10854 3480 10906
rect 3480 10854 3510 10906
rect 3534 10854 3544 10906
rect 3544 10854 3590 10906
rect 3614 10854 3660 10906
rect 3660 10854 3670 10906
rect 3694 10854 3724 10906
rect 3724 10854 3750 10906
rect 3454 10852 3510 10854
rect 3534 10852 3590 10854
rect 3614 10852 3670 10854
rect 3694 10852 3750 10854
rect 2502 9016 2558 9072
rect 2318 4664 2374 4720
rect 1766 4392 1822 4448
rect 2778 8880 2834 8936
rect 3454 9818 3510 9820
rect 3534 9818 3590 9820
rect 3614 9818 3670 9820
rect 3694 9818 3750 9820
rect 3454 9766 3480 9818
rect 3480 9766 3510 9818
rect 3534 9766 3544 9818
rect 3544 9766 3590 9818
rect 3614 9766 3660 9818
rect 3660 9766 3670 9818
rect 3694 9766 3724 9818
rect 3724 9766 3750 9818
rect 3454 9764 3510 9766
rect 3534 9764 3590 9766
rect 3614 9764 3670 9766
rect 3694 9764 3750 9766
rect 3698 9424 3754 9480
rect 3454 8730 3510 8732
rect 3534 8730 3590 8732
rect 3614 8730 3670 8732
rect 3694 8730 3750 8732
rect 3454 8678 3480 8730
rect 3480 8678 3510 8730
rect 3534 8678 3544 8730
rect 3544 8678 3590 8730
rect 3614 8678 3660 8730
rect 3660 8678 3670 8730
rect 3694 8678 3724 8730
rect 3724 8678 3750 8730
rect 3454 8676 3510 8678
rect 3534 8676 3590 8678
rect 3614 8676 3670 8678
rect 3694 8676 3750 8678
rect 2778 6740 2780 6760
rect 2780 6740 2832 6760
rect 2832 6740 2834 6760
rect 2778 6704 2834 6740
rect 3146 7384 3202 7440
rect 3454 7642 3510 7644
rect 3534 7642 3590 7644
rect 3614 7642 3670 7644
rect 3694 7642 3750 7644
rect 3454 7590 3480 7642
rect 3480 7590 3510 7642
rect 3534 7590 3544 7642
rect 3544 7590 3590 7642
rect 3614 7590 3660 7642
rect 3660 7590 3670 7642
rect 3694 7590 3724 7642
rect 3724 7590 3750 7642
rect 3454 7588 3510 7590
rect 3534 7588 3590 7590
rect 3614 7588 3670 7590
rect 3694 7588 3750 7590
rect 3974 8472 4030 8528
rect 4986 15000 5042 15056
rect 5953 16890 6009 16892
rect 6033 16890 6089 16892
rect 6113 16890 6169 16892
rect 6193 16890 6249 16892
rect 5953 16838 5979 16890
rect 5979 16838 6009 16890
rect 6033 16838 6043 16890
rect 6043 16838 6089 16890
rect 6113 16838 6159 16890
rect 6159 16838 6169 16890
rect 6193 16838 6223 16890
rect 6223 16838 6249 16890
rect 5953 16836 6009 16838
rect 6033 16836 6089 16838
rect 6113 16836 6169 16838
rect 6193 16836 6249 16838
rect 5953 15802 6009 15804
rect 6033 15802 6089 15804
rect 6113 15802 6169 15804
rect 6193 15802 6249 15804
rect 5953 15750 5979 15802
rect 5979 15750 6009 15802
rect 6033 15750 6043 15802
rect 6043 15750 6089 15802
rect 6113 15750 6159 15802
rect 6159 15750 6169 15802
rect 6193 15750 6223 15802
rect 6223 15750 6249 15802
rect 5953 15748 6009 15750
rect 6033 15748 6089 15750
rect 6113 15748 6169 15750
rect 6193 15748 6249 15750
rect 6458 15544 6514 15600
rect 5953 14714 6009 14716
rect 6033 14714 6089 14716
rect 6113 14714 6169 14716
rect 6193 14714 6249 14716
rect 5953 14662 5979 14714
rect 5979 14662 6009 14714
rect 6033 14662 6043 14714
rect 6043 14662 6089 14714
rect 6113 14662 6159 14714
rect 6159 14662 6169 14714
rect 6193 14662 6223 14714
rect 6223 14662 6249 14714
rect 5953 14660 6009 14662
rect 6033 14660 6089 14662
rect 6113 14660 6169 14662
rect 6193 14660 6249 14662
rect 2594 4120 2650 4176
rect 1674 3476 1676 3496
rect 1676 3476 1728 3496
rect 1728 3476 1730 3496
rect 1674 3440 1730 3476
rect 2410 3440 2466 3496
rect 1858 2896 1914 2952
rect 1582 2760 1638 2816
rect 3454 6554 3510 6556
rect 3534 6554 3590 6556
rect 3614 6554 3670 6556
rect 3694 6554 3750 6556
rect 3454 6502 3480 6554
rect 3480 6502 3510 6554
rect 3534 6502 3544 6554
rect 3544 6502 3590 6554
rect 3614 6502 3660 6554
rect 3660 6502 3670 6554
rect 3694 6502 3724 6554
rect 3724 6502 3750 6554
rect 3454 6500 3510 6502
rect 3534 6500 3590 6502
rect 3614 6500 3670 6502
rect 3694 6500 3750 6502
rect 4526 8880 4582 8936
rect 4434 8472 4490 8528
rect 3454 5466 3510 5468
rect 3534 5466 3590 5468
rect 3614 5466 3670 5468
rect 3694 5466 3750 5468
rect 3454 5414 3480 5466
rect 3480 5414 3510 5466
rect 3534 5414 3544 5466
rect 3544 5414 3590 5466
rect 3614 5414 3660 5466
rect 3660 5414 3670 5466
rect 3694 5414 3724 5466
rect 3724 5414 3750 5466
rect 3454 5412 3510 5414
rect 3534 5412 3590 5414
rect 3614 5412 3670 5414
rect 3694 5412 3750 5414
rect 3454 4378 3510 4380
rect 3534 4378 3590 4380
rect 3614 4378 3670 4380
rect 3694 4378 3750 4380
rect 3454 4326 3480 4378
rect 3480 4326 3510 4378
rect 3534 4326 3544 4378
rect 3544 4326 3590 4378
rect 3614 4326 3660 4378
rect 3660 4326 3670 4378
rect 3694 4326 3724 4378
rect 3724 4326 3750 4378
rect 3454 4324 3510 4326
rect 3534 4324 3590 4326
rect 3614 4324 3670 4326
rect 3694 4324 3750 4326
rect 3330 4020 3332 4040
rect 3332 4020 3384 4040
rect 3384 4020 3386 4040
rect 3330 3984 3386 4020
rect 3454 3290 3510 3292
rect 3534 3290 3590 3292
rect 3614 3290 3670 3292
rect 3694 3290 3750 3292
rect 3454 3238 3480 3290
rect 3480 3238 3510 3290
rect 3534 3238 3544 3290
rect 3544 3238 3590 3290
rect 3614 3238 3660 3290
rect 3660 3238 3670 3290
rect 3694 3238 3724 3290
rect 3724 3238 3750 3290
rect 3454 3236 3510 3238
rect 3534 3236 3590 3238
rect 3614 3236 3670 3238
rect 3694 3236 3750 3238
rect 2962 2352 3018 2408
rect 2870 1400 2926 1456
rect 5078 9868 5080 9888
rect 5080 9868 5132 9888
rect 5132 9868 5134 9888
rect 5078 9832 5134 9868
rect 4894 8880 4950 8936
rect 4986 7656 5042 7712
rect 7102 16632 7158 16688
rect 5953 13626 6009 13628
rect 6033 13626 6089 13628
rect 6113 13626 6169 13628
rect 6193 13626 6249 13628
rect 5953 13574 5979 13626
rect 5979 13574 6009 13626
rect 6033 13574 6043 13626
rect 6043 13574 6089 13626
rect 6113 13574 6159 13626
rect 6159 13574 6169 13626
rect 6193 13574 6223 13626
rect 6223 13574 6249 13626
rect 5953 13572 6009 13574
rect 6033 13572 6089 13574
rect 6113 13572 6169 13574
rect 6193 13572 6249 13574
rect 5953 12538 6009 12540
rect 6033 12538 6089 12540
rect 6113 12538 6169 12540
rect 6193 12538 6249 12540
rect 5953 12486 5979 12538
rect 5979 12486 6009 12538
rect 6033 12486 6043 12538
rect 6043 12486 6089 12538
rect 6113 12486 6159 12538
rect 6159 12486 6169 12538
rect 6193 12486 6223 12538
rect 6223 12486 6249 12538
rect 5953 12484 6009 12486
rect 6033 12484 6089 12486
rect 6113 12484 6169 12486
rect 6193 12484 6249 12486
rect 5630 11192 5686 11248
rect 5953 11450 6009 11452
rect 6033 11450 6089 11452
rect 6113 11450 6169 11452
rect 6193 11450 6249 11452
rect 5953 11398 5979 11450
rect 5979 11398 6009 11450
rect 6033 11398 6043 11450
rect 6043 11398 6089 11450
rect 6113 11398 6159 11450
rect 6159 11398 6169 11450
rect 6193 11398 6223 11450
rect 6223 11398 6249 11450
rect 5953 11396 6009 11398
rect 6033 11396 6089 11398
rect 6113 11396 6169 11398
rect 6193 11396 6249 11398
rect 5814 10648 5870 10704
rect 4894 6704 4950 6760
rect 4802 5208 4858 5264
rect 5953 10362 6009 10364
rect 6033 10362 6089 10364
rect 6113 10362 6169 10364
rect 6193 10362 6249 10364
rect 5953 10310 5979 10362
rect 5979 10310 6009 10362
rect 6033 10310 6043 10362
rect 6043 10310 6089 10362
rect 6113 10310 6159 10362
rect 6159 10310 6169 10362
rect 6193 10310 6223 10362
rect 6223 10310 6249 10362
rect 5953 10308 6009 10310
rect 6033 10308 6089 10310
rect 6113 10308 6169 10310
rect 6193 10308 6249 10310
rect 6458 10412 6460 10432
rect 6460 10412 6512 10432
rect 6512 10412 6514 10432
rect 6458 10376 6514 10412
rect 7286 15852 7288 15872
rect 7288 15852 7340 15872
rect 7340 15852 7342 15872
rect 7286 15816 7342 15852
rect 5953 9274 6009 9276
rect 6033 9274 6089 9276
rect 6113 9274 6169 9276
rect 6193 9274 6249 9276
rect 5953 9222 5979 9274
rect 5979 9222 6009 9274
rect 6033 9222 6043 9274
rect 6043 9222 6089 9274
rect 6113 9222 6159 9274
rect 6159 9222 6169 9274
rect 6193 9222 6223 9274
rect 6223 9222 6249 9274
rect 5953 9220 6009 9222
rect 6033 9220 6089 9222
rect 6113 9220 6169 9222
rect 6193 9220 6249 9222
rect 5814 9016 5870 9072
rect 5953 8186 6009 8188
rect 6033 8186 6089 8188
rect 6113 8186 6169 8188
rect 6193 8186 6249 8188
rect 5953 8134 5979 8186
rect 5979 8134 6009 8186
rect 6033 8134 6043 8186
rect 6043 8134 6089 8186
rect 6113 8134 6159 8186
rect 6159 8134 6169 8186
rect 6193 8134 6223 8186
rect 6223 8134 6249 8186
rect 5953 8132 6009 8134
rect 6033 8132 6089 8134
rect 6113 8132 6169 8134
rect 6193 8132 6249 8134
rect 5630 7284 5632 7304
rect 5632 7284 5684 7304
rect 5684 7284 5686 7304
rect 5630 7248 5686 7284
rect 6090 7828 6092 7848
rect 6092 7828 6144 7848
rect 6144 7828 6146 7848
rect 6090 7792 6146 7828
rect 5953 7098 6009 7100
rect 6033 7098 6089 7100
rect 6113 7098 6169 7100
rect 6193 7098 6249 7100
rect 5953 7046 5979 7098
rect 5979 7046 6009 7098
rect 6033 7046 6043 7098
rect 6043 7046 6089 7098
rect 6113 7046 6159 7098
rect 6159 7046 6169 7098
rect 6193 7046 6223 7098
rect 6223 7046 6249 7098
rect 5953 7044 6009 7046
rect 6033 7044 6089 7046
rect 6113 7044 6169 7046
rect 6193 7044 6249 7046
rect 6826 11192 6882 11248
rect 6734 10648 6790 10704
rect 6550 8336 6606 8392
rect 6550 7948 6606 7984
rect 6550 7928 6552 7948
rect 6552 7928 6604 7948
rect 6604 7928 6606 7948
rect 6550 7656 6606 7712
rect 6550 7384 6606 7440
rect 6642 7112 6698 7168
rect 6550 6840 6606 6896
rect 5953 6010 6009 6012
rect 6033 6010 6089 6012
rect 6113 6010 6169 6012
rect 6193 6010 6249 6012
rect 5953 5958 5979 6010
rect 5979 5958 6009 6010
rect 6033 5958 6043 6010
rect 6043 5958 6089 6010
rect 6113 5958 6159 6010
rect 6159 5958 6169 6010
rect 6193 5958 6223 6010
rect 6223 5958 6249 6010
rect 5953 5956 6009 5958
rect 6033 5956 6089 5958
rect 6113 5956 6169 5958
rect 6193 5956 6249 5958
rect 4802 3440 4858 3496
rect 4526 3168 4582 3224
rect 3454 2202 3510 2204
rect 3534 2202 3590 2204
rect 3614 2202 3670 2204
rect 3694 2202 3750 2204
rect 3454 2150 3480 2202
rect 3480 2150 3510 2202
rect 3534 2150 3544 2202
rect 3544 2150 3590 2202
rect 3614 2150 3660 2202
rect 3660 2150 3670 2202
rect 3694 2150 3724 2202
rect 3724 2150 3750 2202
rect 3454 2148 3510 2150
rect 3534 2148 3590 2150
rect 3614 2148 3670 2150
rect 3694 2148 3750 2150
rect 4802 2796 4804 2816
rect 4804 2796 4856 2816
rect 4856 2796 4858 2816
rect 4802 2760 4858 2796
rect 5170 3168 5226 3224
rect 5953 4922 6009 4924
rect 6033 4922 6089 4924
rect 6113 4922 6169 4924
rect 6193 4922 6249 4924
rect 5953 4870 5979 4922
rect 5979 4870 6009 4922
rect 6033 4870 6043 4922
rect 6043 4870 6089 4922
rect 6113 4870 6159 4922
rect 6159 4870 6169 4922
rect 6193 4870 6223 4922
rect 6223 4870 6249 4922
rect 5953 4868 6009 4870
rect 6033 4868 6089 4870
rect 6113 4868 6169 4870
rect 6193 4868 6249 4870
rect 6366 4528 6422 4584
rect 5538 4020 5540 4040
rect 5540 4020 5592 4040
rect 5592 4020 5594 4040
rect 5538 3984 5594 4020
rect 5446 3304 5502 3360
rect 5953 3834 6009 3836
rect 6033 3834 6089 3836
rect 6113 3834 6169 3836
rect 6193 3834 6249 3836
rect 5953 3782 5979 3834
rect 5979 3782 6009 3834
rect 6033 3782 6043 3834
rect 6043 3782 6089 3834
rect 6113 3782 6159 3834
rect 6159 3782 6169 3834
rect 6193 3782 6223 3834
rect 6223 3782 6249 3834
rect 5953 3780 6009 3782
rect 6033 3780 6089 3782
rect 6113 3780 6169 3782
rect 6193 3780 6249 3782
rect 6182 3032 6238 3088
rect 5953 2746 6009 2748
rect 6033 2746 6089 2748
rect 6113 2746 6169 2748
rect 6193 2746 6249 2748
rect 5953 2694 5979 2746
rect 5979 2694 6009 2746
rect 6033 2694 6043 2746
rect 6043 2694 6089 2746
rect 6113 2694 6159 2746
rect 6159 2694 6169 2746
rect 6193 2694 6223 2746
rect 6223 2694 6249 2746
rect 5953 2692 6009 2694
rect 6033 2692 6089 2694
rect 6113 2692 6169 2694
rect 6193 2692 6249 2694
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8478 17434
rect 8478 17382 8508 17434
rect 8532 17382 8542 17434
rect 8542 17382 8588 17434
rect 8612 17382 8658 17434
rect 8658 17382 8668 17434
rect 8692 17382 8722 17434
rect 8722 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 7378 12708 7434 12744
rect 7378 12688 7380 12708
rect 7380 12688 7432 12708
rect 7432 12688 7434 12708
rect 6918 9016 6974 9072
rect 7102 8744 7158 8800
rect 7010 7928 7066 7984
rect 6826 6976 6882 7032
rect 7286 9832 7342 9888
rect 7654 9832 7710 9888
rect 7562 8236 7564 8256
rect 7564 8236 7616 8256
rect 7616 8236 7618 8256
rect 7562 8200 7618 8236
rect 7746 8064 7802 8120
rect 6826 5244 6828 5264
rect 6828 5244 6880 5264
rect 6880 5244 6882 5264
rect 6826 5208 6882 5244
rect 6458 3052 6514 3088
rect 6458 3032 6460 3052
rect 6460 3032 6512 3052
rect 6512 3032 6514 3052
rect 6642 3032 6698 3088
rect 6550 2624 6606 2680
rect 6918 2896 6974 2952
rect 6734 2760 6790 2816
rect 7286 2896 7342 2952
rect 8942 16904 8998 16960
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8478 16346
rect 8478 16294 8508 16346
rect 8532 16294 8542 16346
rect 8542 16294 8588 16346
rect 8612 16294 8658 16346
rect 8658 16294 8668 16346
rect 8692 16294 8722 16346
rect 8722 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8478 15258
rect 8478 15206 8508 15258
rect 8532 15206 8542 15258
rect 8542 15206 8588 15258
rect 8612 15206 8658 15258
rect 8658 15206 8668 15258
rect 8692 15206 8722 15258
rect 8722 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8942 15000 8998 15056
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8478 14170
rect 8478 14118 8508 14170
rect 8532 14118 8542 14170
rect 8542 14118 8588 14170
rect 8612 14118 8658 14170
rect 8658 14118 8668 14170
rect 8692 14118 8722 14170
rect 8722 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8478 13082
rect 8478 13030 8508 13082
rect 8532 13030 8542 13082
rect 8542 13030 8588 13082
rect 8612 13030 8658 13082
rect 8658 13030 8668 13082
rect 8692 13030 8722 13082
rect 8722 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 8390 12416 8446 12472
rect 8298 12280 8354 12336
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8478 11994
rect 8478 11942 8508 11994
rect 8532 11942 8542 11994
rect 8542 11942 8588 11994
rect 8612 11942 8658 11994
rect 8658 11942 8668 11994
rect 8692 11942 8722 11994
rect 8722 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 9126 12824 9182 12880
rect 8298 11228 8300 11248
rect 8300 11228 8352 11248
rect 8352 11228 8354 11248
rect 8298 11192 8354 11228
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8478 10906
rect 8478 10854 8508 10906
rect 8532 10854 8542 10906
rect 8542 10854 8588 10906
rect 8612 10854 8658 10906
rect 8658 10854 8668 10906
rect 8692 10854 8722 10906
rect 8722 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8478 9818
rect 8478 9766 8508 9818
rect 8532 9766 8542 9818
rect 8542 9766 8588 9818
rect 8612 9766 8658 9818
rect 8658 9766 8668 9818
rect 8692 9766 8722 9818
rect 8722 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8478 8730
rect 8478 8678 8508 8730
rect 8532 8678 8542 8730
rect 8542 8678 8588 8730
rect 8612 8678 8658 8730
rect 8658 8678 8668 8730
rect 8692 8678 8722 8730
rect 8722 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8666 8472 8722 8528
rect 8390 7928 8446 7984
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8478 7642
rect 8478 7590 8508 7642
rect 8532 7590 8542 7642
rect 8542 7590 8588 7642
rect 8612 7590 8658 7642
rect 8658 7590 8668 7642
rect 8692 7590 8722 7642
rect 8722 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8298 7112 8354 7168
rect 8298 6996 8354 7032
rect 8298 6976 8300 6996
rect 8300 6976 8352 6996
rect 8352 6976 8354 6996
rect 7654 3168 7710 3224
rect 7838 3712 7894 3768
rect 7930 3304 7986 3360
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8478 6554
rect 8478 6502 8508 6554
rect 8532 6502 8542 6554
rect 8542 6502 8588 6554
rect 8612 6502 8658 6554
rect 8658 6502 8668 6554
rect 8692 6502 8722 6554
rect 8722 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 8942 8084 8998 8120
rect 8942 8064 8944 8084
rect 8944 8064 8996 8084
rect 8996 8064 8998 8084
rect 8942 7948 8998 7984
rect 8942 7928 8944 7948
rect 8944 7928 8996 7948
rect 8996 7928 8998 7948
rect 8942 6196 8944 6216
rect 8944 6196 8996 6216
rect 8996 6196 8998 6216
rect 8942 6160 8998 6196
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8478 5466
rect 8478 5414 8508 5466
rect 8532 5414 8542 5466
rect 8542 5414 8588 5466
rect 8612 5414 8658 5466
rect 8658 5414 8668 5466
rect 8692 5414 8722 5466
rect 8722 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8298 4664 8354 4720
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8478 4378
rect 8478 4326 8508 4378
rect 8532 4326 8542 4378
rect 8542 4326 8588 4378
rect 8612 4326 8658 4378
rect 8658 4326 8668 4378
rect 8692 4326 8722 4378
rect 8722 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 9218 10376 9274 10432
rect 9494 12688 9550 12744
rect 9770 14068 9826 14104
rect 9770 14048 9772 14068
rect 9772 14048 9824 14068
rect 9824 14048 9826 14068
rect 9402 12436 9458 12472
rect 9402 12416 9404 12436
rect 9404 12416 9456 12436
rect 9456 12416 9458 12436
rect 9954 12824 10010 12880
rect 9494 11736 9550 11792
rect 9586 10920 9642 10976
rect 10966 17040 11022 17096
rect 10950 16890 11006 16892
rect 11030 16890 11086 16892
rect 11110 16890 11166 16892
rect 11190 16890 11246 16892
rect 10950 16838 10976 16890
rect 10976 16838 11006 16890
rect 11030 16838 11040 16890
rect 11040 16838 11086 16890
rect 11110 16838 11156 16890
rect 11156 16838 11166 16890
rect 11190 16838 11220 16890
rect 11220 16838 11246 16890
rect 10950 16836 11006 16838
rect 11030 16836 11086 16838
rect 11110 16836 11166 16838
rect 11190 16836 11246 16838
rect 9402 7248 9458 7304
rect 8206 2760 8262 2816
rect 8390 3848 8446 3904
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8478 3290
rect 8478 3238 8508 3290
rect 8532 3238 8542 3290
rect 8542 3238 8588 3290
rect 8612 3238 8658 3290
rect 8658 3238 8668 3290
rect 8692 3238 8722 3290
rect 8722 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8666 2760 8722 2816
rect 8758 2624 8814 2680
rect 9126 3712 9182 3768
rect 10322 11756 10378 11792
rect 10322 11736 10324 11756
rect 10324 11736 10376 11756
rect 10376 11736 10378 11756
rect 10950 15802 11006 15804
rect 11030 15802 11086 15804
rect 11110 15802 11166 15804
rect 11190 15802 11246 15804
rect 10950 15750 10976 15802
rect 10976 15750 11006 15802
rect 11030 15750 11040 15802
rect 11040 15750 11086 15802
rect 11110 15750 11156 15802
rect 11156 15750 11166 15802
rect 11190 15750 11220 15802
rect 11220 15750 11246 15802
rect 10950 15748 11006 15750
rect 11030 15748 11086 15750
rect 11110 15748 11166 15750
rect 11190 15748 11246 15750
rect 11334 15564 11390 15600
rect 11334 15544 11336 15564
rect 11336 15544 11388 15564
rect 11388 15544 11390 15564
rect 10950 14714 11006 14716
rect 11030 14714 11086 14716
rect 11110 14714 11166 14716
rect 11190 14714 11246 14716
rect 10950 14662 10976 14714
rect 10976 14662 11006 14714
rect 11030 14662 11040 14714
rect 11040 14662 11086 14714
rect 11110 14662 11156 14714
rect 11156 14662 11166 14714
rect 11190 14662 11220 14714
rect 11220 14662 11246 14714
rect 10950 14660 11006 14662
rect 11030 14660 11086 14662
rect 11110 14660 11166 14662
rect 11190 14660 11246 14662
rect 10950 13626 11006 13628
rect 11030 13626 11086 13628
rect 11110 13626 11166 13628
rect 11190 13626 11246 13628
rect 10950 13574 10976 13626
rect 10976 13574 11006 13626
rect 11030 13574 11040 13626
rect 11040 13574 11086 13626
rect 11110 13574 11156 13626
rect 11156 13574 11166 13626
rect 11190 13574 11220 13626
rect 11220 13574 11246 13626
rect 10950 13572 11006 13574
rect 11030 13572 11086 13574
rect 11110 13572 11166 13574
rect 11190 13572 11246 13574
rect 10950 12538 11006 12540
rect 11030 12538 11086 12540
rect 11110 12538 11166 12540
rect 11190 12538 11246 12540
rect 10950 12486 10976 12538
rect 10976 12486 11006 12538
rect 11030 12486 11040 12538
rect 11040 12486 11086 12538
rect 11110 12486 11156 12538
rect 11156 12486 11166 12538
rect 11190 12486 11220 12538
rect 11220 12486 11246 12538
rect 10950 12484 11006 12486
rect 11030 12484 11086 12486
rect 11110 12484 11166 12486
rect 11190 12484 11246 12486
rect 10046 9016 10102 9072
rect 10230 8880 10286 8936
rect 10414 8608 10470 8664
rect 9678 5208 9734 5264
rect 9586 4564 9588 4584
rect 9588 4564 9640 4584
rect 9640 4564 9642 4584
rect 9586 4528 9642 4564
rect 9586 4120 9642 4176
rect 9034 2488 9090 2544
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8478 2202
rect 8478 2150 8508 2202
rect 8532 2150 8542 2202
rect 8542 2150 8588 2202
rect 8612 2150 8658 2202
rect 8658 2150 8668 2202
rect 8692 2150 8722 2202
rect 8722 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 10414 7928 10470 7984
rect 10782 9424 10838 9480
rect 10950 11450 11006 11452
rect 11030 11450 11086 11452
rect 11110 11450 11166 11452
rect 11190 11450 11246 11452
rect 10950 11398 10976 11450
rect 10976 11398 11006 11450
rect 11030 11398 11040 11450
rect 11040 11398 11086 11450
rect 11110 11398 11156 11450
rect 11156 11398 11166 11450
rect 11190 11398 11220 11450
rect 11220 11398 11246 11450
rect 10950 11396 11006 11398
rect 11030 11396 11086 11398
rect 11110 11396 11166 11398
rect 11190 11396 11246 11398
rect 10950 10362 11006 10364
rect 11030 10362 11086 10364
rect 11110 10362 11166 10364
rect 11190 10362 11246 10364
rect 10950 10310 10976 10362
rect 10976 10310 11006 10362
rect 11030 10310 11040 10362
rect 11040 10310 11086 10362
rect 11110 10310 11156 10362
rect 11156 10310 11166 10362
rect 11190 10310 11220 10362
rect 11220 10310 11246 10362
rect 10950 10308 11006 10310
rect 11030 10308 11086 10310
rect 11110 10308 11166 10310
rect 11190 10308 11246 10310
rect 11426 9560 11482 9616
rect 10950 9274 11006 9276
rect 11030 9274 11086 9276
rect 11110 9274 11166 9276
rect 11190 9274 11246 9276
rect 10950 9222 10976 9274
rect 10976 9222 11006 9274
rect 11030 9222 11040 9274
rect 11040 9222 11086 9274
rect 11110 9222 11156 9274
rect 11156 9222 11166 9274
rect 11190 9222 11220 9274
rect 11220 9222 11246 9274
rect 10950 9220 11006 9222
rect 11030 9220 11086 9222
rect 11110 9220 11166 9222
rect 11190 9220 11246 9222
rect 11334 9016 11390 9072
rect 11426 8880 11482 8936
rect 10322 6160 10378 6216
rect 9770 2916 9826 2952
rect 9770 2896 9772 2916
rect 9772 2896 9824 2916
rect 9824 2896 9826 2916
rect 10414 4664 10470 4720
rect 10950 8186 11006 8188
rect 11030 8186 11086 8188
rect 11110 8186 11166 8188
rect 11190 8186 11246 8188
rect 10950 8134 10976 8186
rect 10976 8134 11006 8186
rect 11030 8134 11040 8186
rect 11040 8134 11086 8186
rect 11110 8134 11156 8186
rect 11156 8134 11166 8186
rect 11190 8134 11220 8186
rect 11220 8134 11246 8186
rect 10950 8132 11006 8134
rect 11030 8132 11086 8134
rect 11110 8132 11166 8134
rect 11190 8132 11246 8134
rect 11794 15444 11796 15464
rect 11796 15444 11848 15464
rect 11848 15444 11850 15464
rect 11794 15408 11850 15444
rect 11610 11736 11666 11792
rect 11518 8064 11574 8120
rect 11610 7792 11666 7848
rect 10950 7098 11006 7100
rect 11030 7098 11086 7100
rect 11110 7098 11166 7100
rect 11190 7098 11246 7100
rect 10950 7046 10976 7098
rect 10976 7046 11006 7098
rect 11030 7046 11040 7098
rect 11040 7046 11086 7098
rect 11110 7046 11156 7098
rect 11156 7046 11166 7098
rect 11190 7046 11220 7098
rect 11220 7046 11246 7098
rect 10950 7044 11006 7046
rect 11030 7044 11086 7046
rect 11110 7044 11166 7046
rect 11190 7044 11246 7046
rect 10414 3440 10470 3496
rect 10950 6010 11006 6012
rect 11030 6010 11086 6012
rect 11110 6010 11166 6012
rect 11190 6010 11246 6012
rect 10950 5958 10976 6010
rect 10976 5958 11006 6010
rect 11030 5958 11040 6010
rect 11040 5958 11086 6010
rect 11110 5958 11156 6010
rect 11156 5958 11166 6010
rect 11190 5958 11220 6010
rect 11220 5958 11246 6010
rect 10950 5956 11006 5958
rect 11030 5956 11086 5958
rect 11110 5956 11166 5958
rect 11190 5956 11246 5958
rect 10950 4922 11006 4924
rect 11030 4922 11086 4924
rect 11110 4922 11166 4924
rect 11190 4922 11246 4924
rect 10950 4870 10976 4922
rect 10976 4870 11006 4922
rect 11030 4870 11040 4922
rect 11040 4870 11086 4922
rect 11110 4870 11156 4922
rect 11156 4870 11166 4922
rect 11190 4870 11220 4922
rect 11220 4870 11246 4922
rect 10950 4868 11006 4870
rect 11030 4868 11086 4870
rect 11110 4868 11166 4870
rect 11190 4868 11246 4870
rect 10782 3848 10838 3904
rect 10950 3834 11006 3836
rect 11030 3834 11086 3836
rect 11110 3834 11166 3836
rect 11190 3834 11246 3836
rect 10950 3782 10976 3834
rect 10976 3782 11006 3834
rect 11030 3782 11040 3834
rect 11040 3782 11086 3834
rect 11110 3782 11156 3834
rect 11156 3782 11166 3834
rect 11190 3782 11220 3834
rect 11220 3782 11246 3834
rect 10950 3780 11006 3782
rect 11030 3780 11086 3782
rect 11110 3780 11166 3782
rect 11190 3780 11246 3782
rect 10950 2746 11006 2748
rect 11030 2746 11086 2748
rect 11110 2746 11166 2748
rect 11190 2746 11246 2748
rect 10950 2694 10976 2746
rect 10976 2694 11006 2746
rect 11030 2694 11040 2746
rect 11040 2694 11086 2746
rect 11110 2694 11156 2746
rect 11156 2694 11166 2746
rect 11190 2694 11220 2746
rect 11220 2694 11246 2746
rect 10950 2692 11006 2694
rect 11030 2692 11086 2694
rect 11110 2692 11166 2694
rect 11190 2692 11246 2694
rect 11794 9696 11850 9752
rect 12162 14048 12218 14104
rect 10782 2488 10838 2544
rect 10690 856 10746 912
rect 12070 9460 12072 9480
rect 12072 9460 12124 9480
rect 12124 9460 12126 9480
rect 12070 9424 12126 9460
rect 12070 7928 12126 7984
rect 12070 2352 12126 2408
rect 12346 8508 12348 8528
rect 12348 8508 12400 8528
rect 12400 8508 12402 8528
rect 12346 8472 12402 8508
rect 12806 8608 12862 8664
rect 12530 3984 12586 4040
rect 12806 4700 12808 4720
rect 12808 4700 12860 4720
rect 12860 4700 12862 4720
rect 12806 4664 12862 4700
rect 12806 3032 12862 3088
rect 13449 17434 13505 17436
rect 13529 17434 13585 17436
rect 13609 17434 13665 17436
rect 13689 17434 13745 17436
rect 13449 17382 13475 17434
rect 13475 17382 13505 17434
rect 13529 17382 13539 17434
rect 13539 17382 13585 17434
rect 13609 17382 13655 17434
rect 13655 17382 13665 17434
rect 13689 17382 13719 17434
rect 13719 17382 13745 17434
rect 13449 17380 13505 17382
rect 13529 17380 13585 17382
rect 13609 17380 13665 17382
rect 13689 17380 13745 17382
rect 13449 16346 13505 16348
rect 13529 16346 13585 16348
rect 13609 16346 13665 16348
rect 13689 16346 13745 16348
rect 13449 16294 13475 16346
rect 13475 16294 13505 16346
rect 13529 16294 13539 16346
rect 13539 16294 13585 16346
rect 13609 16294 13655 16346
rect 13655 16294 13665 16346
rect 13689 16294 13719 16346
rect 13719 16294 13745 16346
rect 13449 16292 13505 16294
rect 13529 16292 13585 16294
rect 13609 16292 13665 16294
rect 13689 16292 13745 16294
rect 13449 15258 13505 15260
rect 13529 15258 13585 15260
rect 13609 15258 13665 15260
rect 13689 15258 13745 15260
rect 13449 15206 13475 15258
rect 13475 15206 13505 15258
rect 13529 15206 13539 15258
rect 13539 15206 13585 15258
rect 13609 15206 13655 15258
rect 13655 15206 13665 15258
rect 13689 15206 13719 15258
rect 13719 15206 13745 15258
rect 13449 15204 13505 15206
rect 13529 15204 13585 15206
rect 13609 15204 13665 15206
rect 13689 15204 13745 15206
rect 13449 14170 13505 14172
rect 13529 14170 13585 14172
rect 13609 14170 13665 14172
rect 13689 14170 13745 14172
rect 13449 14118 13475 14170
rect 13475 14118 13505 14170
rect 13529 14118 13539 14170
rect 13539 14118 13585 14170
rect 13609 14118 13655 14170
rect 13655 14118 13665 14170
rect 13689 14118 13719 14170
rect 13719 14118 13745 14170
rect 13449 14116 13505 14118
rect 13529 14116 13585 14118
rect 13609 14116 13665 14118
rect 13689 14116 13745 14118
rect 13449 13082 13505 13084
rect 13529 13082 13585 13084
rect 13609 13082 13665 13084
rect 13689 13082 13745 13084
rect 13449 13030 13475 13082
rect 13475 13030 13505 13082
rect 13529 13030 13539 13082
rect 13539 13030 13585 13082
rect 13609 13030 13655 13082
rect 13655 13030 13665 13082
rect 13689 13030 13719 13082
rect 13719 13030 13745 13082
rect 13449 13028 13505 13030
rect 13529 13028 13585 13030
rect 13609 13028 13665 13030
rect 13689 13028 13745 13030
rect 13449 11994 13505 11996
rect 13529 11994 13585 11996
rect 13609 11994 13665 11996
rect 13689 11994 13745 11996
rect 13449 11942 13475 11994
rect 13475 11942 13505 11994
rect 13529 11942 13539 11994
rect 13539 11942 13585 11994
rect 13609 11942 13655 11994
rect 13655 11942 13665 11994
rect 13689 11942 13719 11994
rect 13719 11942 13745 11994
rect 13449 11940 13505 11942
rect 13529 11940 13585 11942
rect 13609 11940 13665 11942
rect 13689 11940 13745 11942
rect 13449 10906 13505 10908
rect 13529 10906 13585 10908
rect 13609 10906 13665 10908
rect 13689 10906 13745 10908
rect 13449 10854 13475 10906
rect 13475 10854 13505 10906
rect 13529 10854 13539 10906
rect 13539 10854 13585 10906
rect 13609 10854 13655 10906
rect 13655 10854 13665 10906
rect 13689 10854 13719 10906
rect 13719 10854 13745 10906
rect 13449 10852 13505 10854
rect 13529 10852 13585 10854
rect 13609 10852 13665 10854
rect 13689 10852 13745 10854
rect 13449 9818 13505 9820
rect 13529 9818 13585 9820
rect 13609 9818 13665 9820
rect 13689 9818 13745 9820
rect 13449 9766 13475 9818
rect 13475 9766 13505 9818
rect 13529 9766 13539 9818
rect 13539 9766 13585 9818
rect 13609 9766 13655 9818
rect 13655 9766 13665 9818
rect 13689 9766 13719 9818
rect 13719 9766 13745 9818
rect 13449 9764 13505 9766
rect 13529 9764 13585 9766
rect 13609 9764 13665 9766
rect 13689 9764 13745 9766
rect 13449 8730 13505 8732
rect 13529 8730 13585 8732
rect 13609 8730 13665 8732
rect 13689 8730 13745 8732
rect 13449 8678 13475 8730
rect 13475 8678 13505 8730
rect 13529 8678 13539 8730
rect 13539 8678 13585 8730
rect 13609 8678 13655 8730
rect 13655 8678 13665 8730
rect 13689 8678 13719 8730
rect 13719 8678 13745 8730
rect 13449 8676 13505 8678
rect 13529 8676 13585 8678
rect 13609 8676 13665 8678
rect 13689 8676 13745 8678
rect 13449 7642 13505 7644
rect 13529 7642 13585 7644
rect 13609 7642 13665 7644
rect 13689 7642 13745 7644
rect 13449 7590 13475 7642
rect 13475 7590 13505 7642
rect 13529 7590 13539 7642
rect 13539 7590 13585 7642
rect 13609 7590 13655 7642
rect 13655 7590 13665 7642
rect 13689 7590 13719 7642
rect 13719 7590 13745 7642
rect 13449 7588 13505 7590
rect 13529 7588 13585 7590
rect 13609 7588 13665 7590
rect 13689 7588 13745 7590
rect 13449 6554 13505 6556
rect 13529 6554 13585 6556
rect 13609 6554 13665 6556
rect 13689 6554 13745 6556
rect 13449 6502 13475 6554
rect 13475 6502 13505 6554
rect 13529 6502 13539 6554
rect 13539 6502 13585 6554
rect 13609 6502 13655 6554
rect 13655 6502 13665 6554
rect 13689 6502 13719 6554
rect 13719 6502 13745 6554
rect 13449 6500 13505 6502
rect 13529 6500 13585 6502
rect 13609 6500 13665 6502
rect 13689 6500 13745 6502
rect 13449 5466 13505 5468
rect 13529 5466 13585 5468
rect 13609 5466 13665 5468
rect 13689 5466 13745 5468
rect 13449 5414 13475 5466
rect 13475 5414 13505 5466
rect 13529 5414 13539 5466
rect 13539 5414 13585 5466
rect 13609 5414 13655 5466
rect 13655 5414 13665 5466
rect 13689 5414 13719 5466
rect 13719 5414 13745 5466
rect 13449 5412 13505 5414
rect 13529 5412 13585 5414
rect 13609 5412 13665 5414
rect 13689 5412 13745 5414
rect 13266 3576 13322 3632
rect 13449 4378 13505 4380
rect 13529 4378 13585 4380
rect 13609 4378 13665 4380
rect 13689 4378 13745 4380
rect 13449 4326 13475 4378
rect 13475 4326 13505 4378
rect 13529 4326 13539 4378
rect 13539 4326 13585 4378
rect 13609 4326 13655 4378
rect 13655 4326 13665 4378
rect 13689 4326 13719 4378
rect 13719 4326 13745 4378
rect 13449 4324 13505 4326
rect 13529 4324 13585 4326
rect 13609 4324 13665 4326
rect 13689 4324 13745 4326
rect 13449 3290 13505 3292
rect 13529 3290 13585 3292
rect 13609 3290 13665 3292
rect 13689 3290 13745 3292
rect 13449 3238 13475 3290
rect 13475 3238 13505 3290
rect 13529 3238 13539 3290
rect 13539 3238 13585 3290
rect 13609 3238 13655 3290
rect 13655 3238 13665 3290
rect 13689 3238 13719 3290
rect 13719 3238 13745 3290
rect 13449 3236 13505 3238
rect 13529 3236 13585 3238
rect 13609 3236 13665 3238
rect 13689 3236 13745 3238
rect 13449 2202 13505 2204
rect 13529 2202 13585 2204
rect 13609 2202 13665 2204
rect 13689 2202 13745 2204
rect 13449 2150 13475 2202
rect 13475 2150 13505 2202
rect 13529 2150 13539 2202
rect 13539 2150 13585 2202
rect 13609 2150 13655 2202
rect 13655 2150 13665 2202
rect 13689 2150 13719 2202
rect 13719 2150 13745 2202
rect 13449 2148 13505 2150
rect 13529 2148 13585 2150
rect 13609 2148 13665 2150
rect 13689 2148 13745 2150
rect 14370 15952 14426 16008
rect 14830 16496 14886 16552
rect 15290 9968 15346 10024
rect 14186 2488 14242 2544
rect 14646 2508 14702 2544
rect 14646 2488 14648 2508
rect 14648 2488 14700 2508
rect 14700 2488 14702 2508
rect 1490 448 1546 504
<< metal3 >>
rect 0 19410 800 19440
rect 1945 19410 2011 19413
rect 0 19408 2011 19410
rect 0 19352 1950 19408
rect 2006 19352 2011 19408
rect 0 19350 2011 19352
rect 0 19320 800 19350
rect 1945 19347 2011 19350
rect 0 18458 800 18488
rect 1669 18458 1735 18461
rect 0 18456 1735 18458
rect 0 18400 1674 18456
rect 1730 18400 1735 18456
rect 0 18398 1735 18400
rect 0 18368 800 18398
rect 1669 18395 1735 18398
rect 3442 17440 3762 17441
rect 0 17280 800 17400
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3762 17440
rect 3442 17375 3762 17376
rect 8440 17440 8760 17441
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 17375 8760 17376
rect 13437 17440 13757 17441
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 13437 17375 13757 17376
rect 10961 17098 11027 17101
rect 11462 17098 11468 17100
rect 10961 17096 11468 17098
rect 10961 17040 10966 17096
rect 11022 17040 11468 17096
rect 10961 17038 11468 17040
rect 10961 17035 11027 17038
rect 11462 17036 11468 17038
rect 11532 17036 11538 17100
rect 8937 16962 9003 16965
rect 9070 16962 9076 16964
rect 8937 16960 9076 16962
rect 8937 16904 8942 16960
rect 8998 16904 9076 16960
rect 8937 16902 9076 16904
rect 8937 16899 9003 16902
rect 9070 16900 9076 16902
rect 9140 16900 9146 16964
rect 5941 16896 6261 16897
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 16831 6261 16832
rect 10938 16896 11258 16897
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11258 16896
rect 10938 16831 11258 16832
rect 3417 16690 3483 16693
rect 3969 16690 4035 16693
rect 7097 16690 7163 16693
rect 3417 16688 7163 16690
rect 3417 16632 3422 16688
rect 3478 16632 3974 16688
rect 4030 16632 7102 16688
rect 7158 16632 7163 16688
rect 3417 16630 7163 16632
rect 3417 16627 3483 16630
rect 3969 16627 4035 16630
rect 7097 16627 7163 16630
rect 16400 16600 17200 16720
rect 1761 16554 1827 16557
rect 14825 16554 14891 16557
rect 1761 16552 14891 16554
rect 1761 16496 1766 16552
rect 1822 16496 14830 16552
rect 14886 16496 14891 16552
rect 1761 16494 14891 16496
rect 1761 16491 1827 16494
rect 14825 16491 14891 16494
rect 0 16418 800 16448
rect 1761 16418 1827 16421
rect 0 16416 1827 16418
rect 0 16360 1766 16416
rect 1822 16360 1827 16416
rect 0 16358 1827 16360
rect 0 16328 800 16358
rect 1761 16355 1827 16358
rect 3442 16352 3762 16353
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3762 16352
rect 3442 16287 3762 16288
rect 8440 16352 8760 16353
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 16287 8760 16288
rect 13437 16352 13757 16353
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 13437 16287 13757 16288
rect 565 16010 631 16013
rect 14365 16010 14431 16013
rect 565 16008 14431 16010
rect 565 15952 570 16008
rect 626 15952 14370 16008
rect 14426 15952 14431 16008
rect 565 15950 14431 15952
rect 565 15947 631 15950
rect 14365 15947 14431 15950
rect 7281 15874 7347 15877
rect 7414 15874 7420 15876
rect 7281 15872 7420 15874
rect 7281 15816 7286 15872
rect 7342 15816 7420 15872
rect 7281 15814 7420 15816
rect 7281 15811 7347 15814
rect 7414 15812 7420 15814
rect 7484 15812 7490 15876
rect 5941 15808 6261 15809
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 15743 6261 15744
rect 10938 15808 11258 15809
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11258 15808
rect 10938 15743 11258 15744
rect 6453 15604 6519 15605
rect 6453 15602 6500 15604
rect 6408 15600 6500 15602
rect 6408 15544 6458 15600
rect 6408 15542 6500 15544
rect 6453 15540 6500 15542
rect 6564 15540 6570 15604
rect 11329 15602 11395 15605
rect 11462 15602 11468 15604
rect 11329 15600 11468 15602
rect 11329 15544 11334 15600
rect 11390 15544 11468 15600
rect 11329 15542 11468 15544
rect 6453 15539 6519 15540
rect 11329 15539 11395 15542
rect 11462 15540 11468 15542
rect 11532 15540 11538 15604
rect 0 15466 800 15496
rect 1669 15466 1735 15469
rect 0 15464 1735 15466
rect 0 15408 1674 15464
rect 1730 15408 1735 15464
rect 0 15406 1735 15408
rect 0 15376 800 15406
rect 1669 15403 1735 15406
rect 7414 15404 7420 15468
rect 7484 15466 7490 15468
rect 11789 15466 11855 15469
rect 7484 15464 11855 15466
rect 7484 15408 11794 15464
rect 11850 15408 11855 15464
rect 7484 15406 11855 15408
rect 7484 15404 7490 15406
rect 11789 15403 11855 15406
rect 3442 15264 3762 15265
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3762 15264
rect 3442 15199 3762 15200
rect 8440 15264 8760 15265
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 15199 8760 15200
rect 13437 15264 13757 15265
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 15199 13757 15200
rect 4981 15058 5047 15061
rect 8937 15058 9003 15061
rect 9438 15058 9444 15060
rect 4981 15056 9444 15058
rect 4981 15000 4986 15056
rect 5042 15000 8942 15056
rect 8998 15000 9444 15056
rect 4981 14998 9444 15000
rect 4981 14995 5047 14998
rect 8937 14995 9003 14998
rect 9438 14996 9444 14998
rect 9508 14996 9514 15060
rect 5941 14720 6261 14721
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5941 14655 6261 14656
rect 10938 14720 11258 14721
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11258 14720
rect 10938 14655 11258 14656
rect 0 14378 800 14408
rect 1669 14378 1735 14381
rect 0 14376 1735 14378
rect 0 14320 1674 14376
rect 1730 14320 1735 14376
rect 0 14318 1735 14320
rect 0 14288 800 14318
rect 1669 14315 1735 14318
rect 3442 14176 3762 14177
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3762 14176
rect 3442 14111 3762 14112
rect 8440 14176 8760 14177
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 14111 8760 14112
rect 13437 14176 13757 14177
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 13437 14111 13757 14112
rect 9765 14106 9831 14109
rect 12157 14106 12223 14109
rect 9765 14104 12223 14106
rect 9765 14048 9770 14104
rect 9826 14048 12162 14104
rect 12218 14048 12223 14104
rect 9765 14046 12223 14048
rect 9765 14043 9831 14046
rect 12157 14043 12223 14046
rect 5941 13632 6261 13633
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 13567 6261 13568
rect 10938 13632 11258 13633
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11258 13632
rect 10938 13567 11258 13568
rect 0 13426 800 13456
rect 1853 13426 1919 13429
rect 0 13424 1919 13426
rect 0 13368 1858 13424
rect 1914 13368 1919 13424
rect 0 13366 1919 13368
rect 0 13336 800 13366
rect 1853 13363 1919 13366
rect 3442 13088 3762 13089
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3762 13088
rect 3442 13023 3762 13024
rect 8440 13088 8760 13089
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 13023 8760 13024
rect 13437 13088 13757 13089
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 13437 13023 13757 13024
rect 9121 12882 9187 12885
rect 9949 12882 10015 12885
rect 9121 12880 10015 12882
rect 9121 12824 9126 12880
rect 9182 12824 9954 12880
rect 10010 12824 10015 12880
rect 9121 12822 10015 12824
rect 9121 12819 9187 12822
rect 9949 12819 10015 12822
rect 7373 12746 7439 12749
rect 9489 12746 9555 12749
rect 7373 12744 9555 12746
rect 7373 12688 7378 12744
rect 7434 12688 9494 12744
rect 9550 12688 9555 12744
rect 7373 12686 9555 12688
rect 7373 12683 7439 12686
rect 9489 12683 9555 12686
rect 5941 12544 6261 12545
rect 0 12474 800 12504
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 12479 6261 12480
rect 10938 12544 11258 12545
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11258 12544
rect 10938 12479 11258 12480
rect 1761 12474 1827 12477
rect 0 12472 1827 12474
rect 0 12416 1766 12472
rect 1822 12416 1827 12472
rect 0 12414 1827 12416
rect 0 12384 800 12414
rect 1761 12411 1827 12414
rect 8385 12474 8451 12477
rect 9397 12474 9463 12477
rect 8385 12472 9463 12474
rect 8385 12416 8390 12472
rect 8446 12416 9402 12472
rect 9458 12416 9463 12472
rect 8385 12414 9463 12416
rect 8385 12411 8451 12414
rect 9397 12411 9463 12414
rect 6494 12276 6500 12340
rect 6564 12338 6570 12340
rect 8293 12338 8359 12341
rect 6564 12336 8359 12338
rect 6564 12280 8298 12336
rect 8354 12280 8359 12336
rect 6564 12278 8359 12280
rect 6564 12276 6570 12278
rect 8293 12275 8359 12278
rect 3442 12000 3762 12001
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3762 12000
rect 3442 11935 3762 11936
rect 8440 12000 8760 12001
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 11935 8760 11936
rect 13437 12000 13757 12001
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 13437 11935 13757 11936
rect 9489 11796 9555 11797
rect 9438 11794 9444 11796
rect 9398 11734 9444 11794
rect 9508 11792 9555 11796
rect 9550 11736 9555 11792
rect 9438 11732 9444 11734
rect 9508 11732 9555 11736
rect 9489 11731 9555 11732
rect 10317 11794 10383 11797
rect 11462 11794 11468 11796
rect 10317 11792 11468 11794
rect 10317 11736 10322 11792
rect 10378 11736 11468 11792
rect 10317 11734 11468 11736
rect 10317 11731 10383 11734
rect 11462 11732 11468 11734
rect 11532 11794 11538 11796
rect 11605 11794 11671 11797
rect 11532 11792 11671 11794
rect 11532 11736 11610 11792
rect 11666 11736 11671 11792
rect 11532 11734 11671 11736
rect 11532 11732 11538 11734
rect 11605 11731 11671 11734
rect 5941 11456 6261 11457
rect 0 11386 800 11416
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 11391 6261 11392
rect 10938 11456 11258 11457
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11258 11456
rect 10938 11391 11258 11392
rect 1761 11386 1827 11389
rect 0 11384 1827 11386
rect 0 11328 1766 11384
rect 1822 11328 1827 11384
rect 0 11326 1827 11328
rect 0 11296 800 11326
rect 1761 11323 1827 11326
rect 5625 11250 5691 11253
rect 6821 11250 6887 11253
rect 8293 11250 8359 11253
rect 5625 11248 8359 11250
rect 5625 11192 5630 11248
rect 5686 11192 6826 11248
rect 6882 11192 8298 11248
rect 8354 11192 8359 11248
rect 5625 11190 8359 11192
rect 5625 11187 5691 11190
rect 6821 11187 6887 11190
rect 8293 11187 8359 11190
rect 9070 10916 9076 10980
rect 9140 10978 9146 10980
rect 9581 10978 9647 10981
rect 9140 10976 9647 10978
rect 9140 10920 9586 10976
rect 9642 10920 9647 10976
rect 9140 10918 9647 10920
rect 9140 10916 9146 10918
rect 9581 10915 9647 10918
rect 3442 10912 3762 10913
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3762 10912
rect 3442 10847 3762 10848
rect 8440 10912 8760 10913
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 10847 8760 10848
rect 13437 10912 13757 10913
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13437 10847 13757 10848
rect 5809 10706 5875 10709
rect 6729 10706 6795 10709
rect 5809 10704 6795 10706
rect 5809 10648 5814 10704
rect 5870 10648 6734 10704
rect 6790 10648 6795 10704
rect 5809 10646 6795 10648
rect 5809 10643 5875 10646
rect 6729 10643 6795 10646
rect 0 10434 800 10464
rect 2773 10434 2839 10437
rect 0 10432 2839 10434
rect 0 10376 2778 10432
rect 2834 10376 2839 10432
rect 0 10374 2839 10376
rect 0 10344 800 10374
rect 2773 10371 2839 10374
rect 6453 10434 6519 10437
rect 9213 10434 9279 10437
rect 6453 10432 9279 10434
rect 6453 10376 6458 10432
rect 6514 10376 9218 10432
rect 9274 10376 9279 10432
rect 6453 10374 9279 10376
rect 6453 10371 6519 10374
rect 9213 10371 9279 10374
rect 5941 10368 6261 10369
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5941 10303 6261 10304
rect 10938 10368 11258 10369
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11258 10368
rect 10938 10303 11258 10304
rect 15285 10026 15351 10029
rect 16400 10026 17200 10056
rect 15285 10024 17200 10026
rect 15285 9968 15290 10024
rect 15346 9968 17200 10024
rect 15285 9966 17200 9968
rect 15285 9963 15351 9966
rect 16400 9936 17200 9966
rect 5073 9890 5139 9893
rect 7281 9890 7347 9893
rect 7649 9890 7715 9893
rect 5073 9888 7715 9890
rect 5073 9832 5078 9888
rect 5134 9832 7286 9888
rect 7342 9832 7654 9888
rect 7710 9832 7715 9888
rect 5073 9830 7715 9832
rect 5073 9827 5139 9830
rect 7281 9827 7347 9830
rect 7649 9827 7715 9830
rect 3442 9824 3762 9825
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3762 9824
rect 3442 9759 3762 9760
rect 8440 9824 8760 9825
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 9759 8760 9760
rect 13437 9824 13757 9825
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 13437 9759 13757 9760
rect 11789 9754 11855 9757
rect 11654 9752 11855 9754
rect 11654 9696 11794 9752
rect 11850 9696 11855 9752
rect 11654 9694 11855 9696
rect 1485 9618 1551 9621
rect 11421 9618 11487 9621
rect 11654 9620 11714 9694
rect 11789 9691 11855 9694
rect 1485 9616 11487 9618
rect 1485 9560 1490 9616
rect 1546 9560 11426 9616
rect 11482 9560 11487 9616
rect 1485 9558 11487 9560
rect 1485 9555 1551 9558
rect 11421 9555 11487 9558
rect 11646 9556 11652 9620
rect 11716 9556 11722 9620
rect 0 9482 800 9512
rect 3693 9482 3759 9485
rect 0 9480 3759 9482
rect 0 9424 3698 9480
rect 3754 9424 3759 9480
rect 0 9422 3759 9424
rect 0 9392 800 9422
rect 3693 9419 3759 9422
rect 10777 9482 10843 9485
rect 12065 9482 12131 9485
rect 10777 9480 12131 9482
rect 10777 9424 10782 9480
rect 10838 9424 12070 9480
rect 12126 9424 12131 9480
rect 10777 9422 12131 9424
rect 10777 9419 10843 9422
rect 12065 9419 12131 9422
rect 5941 9280 6261 9281
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 9215 6261 9216
rect 10938 9280 11258 9281
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11258 9280
rect 10938 9215 11258 9216
rect 2497 9074 2563 9077
rect 5809 9074 5875 9077
rect 2497 9072 5875 9074
rect 2497 9016 2502 9072
rect 2558 9016 5814 9072
rect 5870 9016 5875 9072
rect 2497 9014 5875 9016
rect 2497 9011 2563 9014
rect 5809 9011 5875 9014
rect 6913 9074 6979 9077
rect 10041 9074 10107 9077
rect 11329 9074 11395 9077
rect 6913 9072 7114 9074
rect 6913 9016 6918 9072
rect 6974 9016 7114 9072
rect 6913 9014 7114 9016
rect 6913 9011 6979 9014
rect 2773 8938 2839 8941
rect 4521 8938 4587 8941
rect 4889 8938 4955 8941
rect 2773 8936 4955 8938
rect 2773 8880 2778 8936
rect 2834 8880 4526 8936
rect 4582 8880 4894 8936
rect 4950 8880 4955 8936
rect 2773 8878 4955 8880
rect 2773 8875 2839 8878
rect 4521 8875 4587 8878
rect 4889 8875 4955 8878
rect 7054 8805 7114 9014
rect 10041 9072 11395 9074
rect 10041 9016 10046 9072
rect 10102 9016 11334 9072
rect 11390 9016 11395 9072
rect 10041 9014 11395 9016
rect 10041 9011 10107 9014
rect 11329 9011 11395 9014
rect 10225 8938 10291 8941
rect 10358 8938 10364 8940
rect 10225 8936 10364 8938
rect 10225 8880 10230 8936
rect 10286 8880 10364 8936
rect 10225 8878 10364 8880
rect 10225 8875 10291 8878
rect 10358 8876 10364 8878
rect 10428 8938 10434 8940
rect 11421 8938 11487 8941
rect 10428 8936 11487 8938
rect 10428 8880 11426 8936
rect 11482 8880 11487 8936
rect 10428 8878 11487 8880
rect 10428 8876 10434 8878
rect 11421 8875 11487 8878
rect 7054 8800 7163 8805
rect 7054 8744 7102 8800
rect 7158 8744 7163 8800
rect 7054 8742 7163 8744
rect 7097 8739 7163 8742
rect 3442 8736 3762 8737
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3762 8736
rect 3442 8671 3762 8672
rect 8440 8736 8760 8737
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 8671 8760 8672
rect 13437 8736 13757 8737
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13437 8671 13757 8672
rect 10409 8666 10475 8669
rect 12801 8666 12867 8669
rect 10409 8664 12867 8666
rect 10409 8608 10414 8664
rect 10470 8608 12806 8664
rect 12862 8608 12867 8664
rect 10409 8606 12867 8608
rect 10409 8603 10475 8606
rect 12801 8603 12867 8606
rect 3969 8530 4035 8533
rect 4429 8530 4495 8533
rect 8661 8530 8727 8533
rect 12341 8530 12407 8533
rect 3969 8528 8727 8530
rect 3969 8472 3974 8528
rect 4030 8472 4434 8528
rect 4490 8472 8666 8528
rect 8722 8472 8727 8528
rect 3969 8470 8727 8472
rect 3969 8467 4035 8470
rect 4429 8467 4495 8470
rect 8661 8467 8727 8470
rect 11102 8528 12407 8530
rect 11102 8472 12346 8528
rect 12402 8472 12407 8528
rect 11102 8470 12407 8472
rect 0 8394 800 8424
rect 1761 8394 1827 8397
rect 0 8392 1827 8394
rect 0 8336 1766 8392
rect 1822 8336 1827 8392
rect 0 8334 1827 8336
rect 0 8304 800 8334
rect 1761 8331 1827 8334
rect 6545 8394 6611 8397
rect 11102 8394 11162 8470
rect 12341 8467 12407 8470
rect 6545 8392 11162 8394
rect 6545 8336 6550 8392
rect 6606 8336 11162 8392
rect 6545 8334 11162 8336
rect 6545 8331 6611 8334
rect 7414 8196 7420 8260
rect 7484 8258 7490 8260
rect 7557 8258 7623 8261
rect 7484 8256 7623 8258
rect 7484 8200 7562 8256
rect 7618 8200 7623 8256
rect 7484 8198 7623 8200
rect 7484 8196 7490 8198
rect 7557 8195 7623 8198
rect 5941 8192 6261 8193
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5941 8127 6261 8128
rect 10938 8192 11258 8193
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11258 8192
rect 10938 8127 11258 8128
rect 7741 8122 7807 8125
rect 8937 8122 9003 8125
rect 11513 8124 11579 8125
rect 11462 8122 11468 8124
rect 7741 8120 9003 8122
rect 7741 8064 7746 8120
rect 7802 8064 8942 8120
rect 8998 8064 9003 8120
rect 7741 8062 9003 8064
rect 11422 8062 11468 8122
rect 11532 8120 11579 8124
rect 11574 8064 11579 8120
rect 7741 8059 7807 8062
rect 8937 8059 9003 8062
rect 11462 8060 11468 8062
rect 11532 8060 11579 8064
rect 11513 8059 11579 8060
rect 6545 7986 6611 7989
rect 7005 7986 7071 7989
rect 6545 7984 7071 7986
rect 6545 7928 6550 7984
rect 6606 7928 7010 7984
rect 7066 7928 7071 7984
rect 6545 7926 7071 7928
rect 6545 7923 6611 7926
rect 7005 7923 7071 7926
rect 8385 7986 8451 7989
rect 8937 7986 9003 7989
rect 8385 7984 9003 7986
rect 8385 7928 8390 7984
rect 8446 7928 8942 7984
rect 8998 7928 9003 7984
rect 8385 7926 9003 7928
rect 8385 7923 8451 7926
rect 8937 7923 9003 7926
rect 10409 7986 10475 7989
rect 12065 7986 12131 7989
rect 10409 7984 12131 7986
rect 10409 7928 10414 7984
rect 10470 7928 12070 7984
rect 12126 7928 12131 7984
rect 10409 7926 12131 7928
rect 10409 7923 10475 7926
rect 12065 7923 12131 7926
rect 6085 7850 6151 7853
rect 11605 7850 11671 7853
rect 6085 7848 11671 7850
rect 6085 7792 6090 7848
rect 6146 7792 11610 7848
rect 11666 7792 11671 7848
rect 6085 7790 11671 7792
rect 6085 7787 6151 7790
rect 11605 7787 11671 7790
rect 4981 7714 5047 7717
rect 6545 7714 6611 7717
rect 4981 7712 6611 7714
rect 4981 7656 4986 7712
rect 5042 7656 6550 7712
rect 6606 7656 6611 7712
rect 4981 7654 6611 7656
rect 4981 7651 5047 7654
rect 6545 7651 6611 7654
rect 3442 7648 3762 7649
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3762 7648
rect 3442 7583 3762 7584
rect 8440 7648 8760 7649
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 7583 8760 7584
rect 13437 7648 13757 7649
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 7583 13757 7584
rect 0 7442 800 7472
rect 1669 7442 1735 7445
rect 0 7440 1735 7442
rect 0 7384 1674 7440
rect 1730 7384 1735 7440
rect 0 7382 1735 7384
rect 0 7352 800 7382
rect 1669 7379 1735 7382
rect 3141 7442 3207 7445
rect 6545 7442 6611 7445
rect 3141 7440 6611 7442
rect 3141 7384 3146 7440
rect 3202 7384 6550 7440
rect 6606 7384 6611 7440
rect 3141 7382 6611 7384
rect 3141 7379 3207 7382
rect 6545 7379 6611 7382
rect 5625 7306 5691 7309
rect 9397 7306 9463 7309
rect 5625 7304 9463 7306
rect 5625 7248 5630 7304
rect 5686 7248 9402 7304
rect 9458 7248 9463 7304
rect 5625 7246 9463 7248
rect 5625 7243 5691 7246
rect 9397 7243 9463 7246
rect 6637 7170 6703 7173
rect 8293 7170 8359 7173
rect 6637 7168 8359 7170
rect 6637 7112 6642 7168
rect 6698 7112 8298 7168
rect 8354 7112 8359 7168
rect 6637 7110 8359 7112
rect 6637 7107 6703 7110
rect 8293 7107 8359 7110
rect 5941 7104 6261 7105
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 7039 6261 7040
rect 10938 7104 11258 7105
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11258 7104
rect 10938 7039 11258 7040
rect 6821 7034 6887 7037
rect 8293 7034 8359 7037
rect 6548 7032 8359 7034
rect 6548 6976 6826 7032
rect 6882 6976 8298 7032
rect 8354 6976 8359 7032
rect 6548 6974 8359 6976
rect 6548 6901 6608 6974
rect 6821 6971 6887 6974
rect 8293 6971 8359 6974
rect 6545 6896 6611 6901
rect 6545 6840 6550 6896
rect 6606 6840 6611 6896
rect 6545 6835 6611 6840
rect 2773 6762 2839 6765
rect 4889 6762 4955 6765
rect 2773 6760 4955 6762
rect 2773 6704 2778 6760
rect 2834 6704 4894 6760
rect 4950 6704 4955 6760
rect 2773 6702 4955 6704
rect 2773 6699 2839 6702
rect 4889 6699 4955 6702
rect 3442 6560 3762 6561
rect 0 6490 800 6520
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3762 6560
rect 3442 6495 3762 6496
rect 8440 6560 8760 6561
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 6495 8760 6496
rect 13437 6560 13757 6561
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 6495 13757 6496
rect 1669 6490 1735 6493
rect 0 6488 1735 6490
rect 0 6432 1674 6488
rect 1730 6432 1735 6488
rect 0 6430 1735 6432
rect 0 6400 800 6430
rect 1669 6427 1735 6430
rect 8937 6218 9003 6221
rect 10317 6218 10383 6221
rect 11462 6218 11468 6220
rect 8937 6216 11468 6218
rect 8937 6160 8942 6216
rect 8998 6160 10322 6216
rect 10378 6160 11468 6216
rect 8937 6158 11468 6160
rect 8937 6155 9003 6158
rect 10317 6155 10383 6158
rect 11462 6156 11468 6158
rect 11532 6156 11538 6220
rect 5941 6016 6261 6017
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 5951 6261 5952
rect 10938 6016 11258 6017
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11258 6016
rect 10938 5951 11258 5952
rect 3442 5472 3762 5473
rect 0 5402 800 5432
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3762 5472
rect 3442 5407 3762 5408
rect 8440 5472 8760 5473
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 5407 8760 5408
rect 13437 5472 13757 5473
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 13437 5407 13757 5408
rect 2221 5402 2287 5405
rect 0 5400 2287 5402
rect 0 5344 2226 5400
rect 2282 5344 2287 5400
rect 0 5342 2287 5344
rect 0 5312 800 5342
rect 2221 5339 2287 5342
rect 4797 5266 4863 5269
rect 6821 5266 6887 5269
rect 9673 5266 9739 5269
rect 4797 5264 9739 5266
rect 4797 5208 4802 5264
rect 4858 5208 6826 5264
rect 6882 5208 9678 5264
rect 9734 5208 9739 5264
rect 4797 5206 9739 5208
rect 4797 5203 4863 5206
rect 6821 5203 6887 5206
rect 9673 5203 9739 5206
rect 5941 4928 6261 4929
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 5941 4863 6261 4864
rect 10938 4928 11258 4929
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11258 4928
rect 10938 4863 11258 4864
rect 2313 4722 2379 4725
rect 8293 4722 8359 4725
rect 2313 4720 8359 4722
rect 2313 4664 2318 4720
rect 2374 4664 8298 4720
rect 8354 4664 8359 4720
rect 2313 4662 8359 4664
rect 2313 4659 2379 4662
rect 8293 4659 8359 4662
rect 10409 4722 10475 4725
rect 12801 4722 12867 4725
rect 10409 4720 12867 4722
rect 10409 4664 10414 4720
rect 10470 4664 12806 4720
rect 12862 4664 12867 4720
rect 10409 4662 12867 4664
rect 10409 4659 10475 4662
rect 12801 4659 12867 4662
rect 6361 4586 6427 4589
rect 9581 4586 9647 4589
rect 6361 4584 9647 4586
rect 6361 4528 6366 4584
rect 6422 4528 9586 4584
rect 9642 4528 9647 4584
rect 6361 4526 9647 4528
rect 6361 4523 6427 4526
rect 9581 4523 9647 4526
rect 0 4450 800 4480
rect 1761 4450 1827 4453
rect 0 4448 1827 4450
rect 0 4392 1766 4448
rect 1822 4392 1827 4448
rect 0 4390 1827 4392
rect 0 4360 800 4390
rect 1761 4387 1827 4390
rect 3442 4384 3762 4385
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3762 4384
rect 3442 4319 3762 4320
rect 8440 4384 8760 4385
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 4319 8760 4320
rect 13437 4384 13757 4385
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 13437 4319 13757 4320
rect 2589 4178 2655 4181
rect 9581 4178 9647 4181
rect 2589 4176 9647 4178
rect 2589 4120 2594 4176
rect 2650 4120 9586 4176
rect 9642 4120 9647 4176
rect 2589 4118 9647 4120
rect 2589 4115 2655 4118
rect 9581 4115 9647 4118
rect 3325 4042 3391 4045
rect 5533 4042 5599 4045
rect 12525 4042 12591 4045
rect 3325 4040 12591 4042
rect 3325 3984 3330 4040
rect 3386 3984 5538 4040
rect 5594 3984 12530 4040
rect 12586 3984 12591 4040
rect 3325 3982 12591 3984
rect 3325 3979 3391 3982
rect 5533 3979 5599 3982
rect 12525 3979 12591 3982
rect 8385 3906 8451 3909
rect 10777 3906 10843 3909
rect 8385 3904 10843 3906
rect 8385 3848 8390 3904
rect 8446 3848 10782 3904
rect 10838 3848 10843 3904
rect 8385 3846 10843 3848
rect 8385 3843 8451 3846
rect 10777 3843 10843 3846
rect 5941 3840 6261 3841
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 3775 6261 3776
rect 10938 3840 11258 3841
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11258 3840
rect 10938 3775 11258 3776
rect 7833 3770 7899 3773
rect 9121 3770 9187 3773
rect 7833 3768 9187 3770
rect 7833 3712 7838 3768
rect 7894 3712 9126 3768
rect 9182 3712 9187 3768
rect 7833 3710 9187 3712
rect 7833 3707 7899 3710
rect 9121 3707 9187 3710
rect 13261 3634 13327 3637
rect 13261 3632 14658 3634
rect 13261 3576 13266 3632
rect 13322 3576 14658 3632
rect 13261 3574 14658 3576
rect 13261 3571 13327 3574
rect 0 3498 800 3528
rect 1669 3498 1735 3501
rect 0 3496 1735 3498
rect 0 3440 1674 3496
rect 1730 3440 1735 3496
rect 0 3438 1735 3440
rect 0 3408 800 3438
rect 1669 3435 1735 3438
rect 2405 3498 2471 3501
rect 4797 3498 4863 3501
rect 10409 3498 10475 3501
rect 2405 3496 3986 3498
rect 2405 3440 2410 3496
rect 2466 3440 3986 3496
rect 2405 3438 3986 3440
rect 2405 3435 2471 3438
rect 3926 3362 3986 3438
rect 4797 3496 10475 3498
rect 4797 3440 4802 3496
rect 4858 3440 10414 3496
rect 10470 3440 10475 3496
rect 4797 3438 10475 3440
rect 4797 3435 4863 3438
rect 10409 3435 10475 3438
rect 5441 3362 5507 3365
rect 7925 3362 7991 3365
rect 3926 3360 7991 3362
rect 3926 3304 5446 3360
rect 5502 3304 7930 3360
rect 7986 3304 7991 3360
rect 3926 3302 7991 3304
rect 14598 3362 14658 3574
rect 16400 3362 17200 3392
rect 14598 3302 17200 3362
rect 5441 3299 5507 3302
rect 7925 3299 7991 3302
rect 3442 3296 3762 3297
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3762 3296
rect 3442 3231 3762 3232
rect 8440 3296 8760 3297
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 3231 8760 3232
rect 13437 3296 13757 3297
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 16400 3272 17200 3302
rect 13437 3231 13757 3232
rect 4521 3226 4587 3229
rect 5165 3226 5231 3229
rect 7649 3226 7715 3229
rect 4521 3224 7715 3226
rect 4521 3168 4526 3224
rect 4582 3168 5170 3224
rect 5226 3168 7654 3224
rect 7710 3168 7715 3224
rect 4521 3166 7715 3168
rect 4521 3163 4587 3166
rect 5165 3163 5231 3166
rect 7649 3163 7715 3166
rect 6177 3090 6243 3093
rect 6453 3090 6519 3093
rect 6177 3088 6519 3090
rect 6177 3032 6182 3088
rect 6238 3032 6458 3088
rect 6514 3032 6519 3088
rect 6177 3030 6519 3032
rect 6177 3027 6243 3030
rect 6453 3027 6519 3030
rect 6637 3090 6703 3093
rect 12801 3090 12867 3093
rect 6637 3088 12867 3090
rect 6637 3032 6642 3088
rect 6698 3032 12806 3088
rect 12862 3032 12867 3088
rect 6637 3030 12867 3032
rect 6637 3027 6703 3030
rect 12801 3027 12867 3030
rect 1853 2954 1919 2957
rect 6913 2954 6979 2957
rect 1853 2952 6979 2954
rect 1853 2896 1858 2952
rect 1914 2896 6918 2952
rect 6974 2896 6979 2952
rect 1853 2894 6979 2896
rect 1853 2891 1919 2894
rect 6913 2891 6979 2894
rect 7281 2954 7347 2957
rect 9765 2954 9831 2957
rect 7281 2952 9831 2954
rect 7281 2896 7286 2952
rect 7342 2896 9770 2952
rect 9826 2896 9831 2952
rect 7281 2894 9831 2896
rect 7281 2891 7347 2894
rect 9765 2891 9831 2894
rect 1577 2818 1643 2821
rect 4797 2818 4863 2821
rect 1577 2816 4863 2818
rect 1577 2760 1582 2816
rect 1638 2760 4802 2816
rect 4858 2760 4863 2816
rect 1577 2758 4863 2760
rect 1577 2755 1643 2758
rect 4797 2755 4863 2758
rect 6729 2818 6795 2821
rect 8201 2818 8267 2821
rect 6729 2816 8267 2818
rect 6729 2760 6734 2816
rect 6790 2760 8206 2816
rect 8262 2760 8267 2816
rect 6729 2758 8267 2760
rect 6729 2755 6795 2758
rect 8201 2755 8267 2758
rect 8661 2818 8727 2821
rect 8661 2816 9138 2818
rect 8661 2760 8666 2816
rect 8722 2760 9138 2816
rect 8661 2758 9138 2760
rect 8661 2755 8727 2758
rect 5941 2752 6261 2753
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 5941 2687 6261 2688
rect 6545 2682 6611 2685
rect 8753 2682 8819 2685
rect 6545 2680 8819 2682
rect 6545 2624 6550 2680
rect 6606 2624 8758 2680
rect 8814 2624 8819 2680
rect 6545 2622 8819 2624
rect 6545 2619 6611 2622
rect 8753 2619 8819 2622
rect 9078 2549 9138 2758
rect 10938 2752 11258 2753
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11258 2752
rect 10938 2687 11258 2688
rect 9029 2544 9138 2549
rect 9029 2488 9034 2544
rect 9090 2488 9138 2544
rect 9029 2486 9138 2488
rect 10777 2546 10843 2549
rect 14181 2546 14247 2549
rect 14641 2546 14707 2549
rect 10777 2544 14707 2546
rect 10777 2488 10782 2544
rect 10838 2488 14186 2544
rect 14242 2488 14646 2544
rect 14702 2488 14707 2544
rect 10777 2486 14707 2488
rect 9029 2483 9095 2486
rect 10777 2483 10843 2486
rect 14181 2483 14247 2486
rect 14641 2483 14707 2486
rect 0 2410 800 2440
rect 2957 2410 3023 2413
rect 0 2408 3023 2410
rect 0 2352 2962 2408
rect 3018 2352 3023 2408
rect 0 2350 3023 2352
rect 0 2320 800 2350
rect 2957 2347 3023 2350
rect 11646 2348 11652 2412
rect 11716 2410 11722 2412
rect 12065 2410 12131 2413
rect 11716 2408 12131 2410
rect 11716 2352 12070 2408
rect 12126 2352 12131 2408
rect 11716 2350 12131 2352
rect 11716 2348 11722 2350
rect 12065 2347 12131 2350
rect 3442 2208 3762 2209
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3762 2208
rect 3442 2143 3762 2144
rect 8440 2208 8760 2209
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2143 8760 2144
rect 13437 2208 13757 2209
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2143 13757 2144
rect 0 1458 800 1488
rect 2865 1458 2931 1461
rect 0 1456 2931 1458
rect 0 1400 2870 1456
rect 2926 1400 2931 1456
rect 0 1398 2931 1400
rect 0 1368 800 1398
rect 2865 1395 2931 1398
rect 10358 852 10364 916
rect 10428 914 10434 916
rect 10685 914 10751 917
rect 10428 912 10751 914
rect 10428 856 10690 912
rect 10746 856 10751 912
rect 10428 854 10751 856
rect 10428 852 10434 854
rect 10685 851 10751 854
rect 0 506 800 536
rect 1485 506 1551 509
rect 0 504 1551 506
rect 0 448 1490 504
rect 1546 448 1551 504
rect 0 446 1551 448
rect 0 416 800 446
rect 1485 443 1551 446
<< via3 >>
rect 3450 17436 3514 17440
rect 3450 17380 3454 17436
rect 3454 17380 3510 17436
rect 3510 17380 3514 17436
rect 3450 17376 3514 17380
rect 3530 17436 3594 17440
rect 3530 17380 3534 17436
rect 3534 17380 3590 17436
rect 3590 17380 3594 17436
rect 3530 17376 3594 17380
rect 3610 17436 3674 17440
rect 3610 17380 3614 17436
rect 3614 17380 3670 17436
rect 3670 17380 3674 17436
rect 3610 17376 3674 17380
rect 3690 17436 3754 17440
rect 3690 17380 3694 17436
rect 3694 17380 3750 17436
rect 3750 17380 3754 17436
rect 3690 17376 3754 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 13445 17436 13509 17440
rect 13445 17380 13449 17436
rect 13449 17380 13505 17436
rect 13505 17380 13509 17436
rect 13445 17376 13509 17380
rect 13525 17436 13589 17440
rect 13525 17380 13529 17436
rect 13529 17380 13585 17436
rect 13585 17380 13589 17436
rect 13525 17376 13589 17380
rect 13605 17436 13669 17440
rect 13605 17380 13609 17436
rect 13609 17380 13665 17436
rect 13665 17380 13669 17436
rect 13605 17376 13669 17380
rect 13685 17436 13749 17440
rect 13685 17380 13689 17436
rect 13689 17380 13745 17436
rect 13745 17380 13749 17436
rect 13685 17376 13749 17380
rect 11468 17036 11532 17100
rect 9076 16900 9140 16964
rect 5949 16892 6013 16896
rect 5949 16836 5953 16892
rect 5953 16836 6009 16892
rect 6009 16836 6013 16892
rect 5949 16832 6013 16836
rect 6029 16892 6093 16896
rect 6029 16836 6033 16892
rect 6033 16836 6089 16892
rect 6089 16836 6093 16892
rect 6029 16832 6093 16836
rect 6109 16892 6173 16896
rect 6109 16836 6113 16892
rect 6113 16836 6169 16892
rect 6169 16836 6173 16892
rect 6109 16832 6173 16836
rect 6189 16892 6253 16896
rect 6189 16836 6193 16892
rect 6193 16836 6249 16892
rect 6249 16836 6253 16892
rect 6189 16832 6253 16836
rect 10946 16892 11010 16896
rect 10946 16836 10950 16892
rect 10950 16836 11006 16892
rect 11006 16836 11010 16892
rect 10946 16832 11010 16836
rect 11026 16892 11090 16896
rect 11026 16836 11030 16892
rect 11030 16836 11086 16892
rect 11086 16836 11090 16892
rect 11026 16832 11090 16836
rect 11106 16892 11170 16896
rect 11106 16836 11110 16892
rect 11110 16836 11166 16892
rect 11166 16836 11170 16892
rect 11106 16832 11170 16836
rect 11186 16892 11250 16896
rect 11186 16836 11190 16892
rect 11190 16836 11246 16892
rect 11246 16836 11250 16892
rect 11186 16832 11250 16836
rect 3450 16348 3514 16352
rect 3450 16292 3454 16348
rect 3454 16292 3510 16348
rect 3510 16292 3514 16348
rect 3450 16288 3514 16292
rect 3530 16348 3594 16352
rect 3530 16292 3534 16348
rect 3534 16292 3590 16348
rect 3590 16292 3594 16348
rect 3530 16288 3594 16292
rect 3610 16348 3674 16352
rect 3610 16292 3614 16348
rect 3614 16292 3670 16348
rect 3670 16292 3674 16348
rect 3610 16288 3674 16292
rect 3690 16348 3754 16352
rect 3690 16292 3694 16348
rect 3694 16292 3750 16348
rect 3750 16292 3754 16348
rect 3690 16288 3754 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 13445 16348 13509 16352
rect 13445 16292 13449 16348
rect 13449 16292 13505 16348
rect 13505 16292 13509 16348
rect 13445 16288 13509 16292
rect 13525 16348 13589 16352
rect 13525 16292 13529 16348
rect 13529 16292 13585 16348
rect 13585 16292 13589 16348
rect 13525 16288 13589 16292
rect 13605 16348 13669 16352
rect 13605 16292 13609 16348
rect 13609 16292 13665 16348
rect 13665 16292 13669 16348
rect 13605 16288 13669 16292
rect 13685 16348 13749 16352
rect 13685 16292 13689 16348
rect 13689 16292 13745 16348
rect 13745 16292 13749 16348
rect 13685 16288 13749 16292
rect 7420 15812 7484 15876
rect 5949 15804 6013 15808
rect 5949 15748 5953 15804
rect 5953 15748 6009 15804
rect 6009 15748 6013 15804
rect 5949 15744 6013 15748
rect 6029 15804 6093 15808
rect 6029 15748 6033 15804
rect 6033 15748 6089 15804
rect 6089 15748 6093 15804
rect 6029 15744 6093 15748
rect 6109 15804 6173 15808
rect 6109 15748 6113 15804
rect 6113 15748 6169 15804
rect 6169 15748 6173 15804
rect 6109 15744 6173 15748
rect 6189 15804 6253 15808
rect 6189 15748 6193 15804
rect 6193 15748 6249 15804
rect 6249 15748 6253 15804
rect 6189 15744 6253 15748
rect 10946 15804 11010 15808
rect 10946 15748 10950 15804
rect 10950 15748 11006 15804
rect 11006 15748 11010 15804
rect 10946 15744 11010 15748
rect 11026 15804 11090 15808
rect 11026 15748 11030 15804
rect 11030 15748 11086 15804
rect 11086 15748 11090 15804
rect 11026 15744 11090 15748
rect 11106 15804 11170 15808
rect 11106 15748 11110 15804
rect 11110 15748 11166 15804
rect 11166 15748 11170 15804
rect 11106 15744 11170 15748
rect 11186 15804 11250 15808
rect 11186 15748 11190 15804
rect 11190 15748 11246 15804
rect 11246 15748 11250 15804
rect 11186 15744 11250 15748
rect 6500 15600 6564 15604
rect 6500 15544 6514 15600
rect 6514 15544 6564 15600
rect 6500 15540 6564 15544
rect 11468 15540 11532 15604
rect 7420 15404 7484 15468
rect 3450 15260 3514 15264
rect 3450 15204 3454 15260
rect 3454 15204 3510 15260
rect 3510 15204 3514 15260
rect 3450 15200 3514 15204
rect 3530 15260 3594 15264
rect 3530 15204 3534 15260
rect 3534 15204 3590 15260
rect 3590 15204 3594 15260
rect 3530 15200 3594 15204
rect 3610 15260 3674 15264
rect 3610 15204 3614 15260
rect 3614 15204 3670 15260
rect 3670 15204 3674 15260
rect 3610 15200 3674 15204
rect 3690 15260 3754 15264
rect 3690 15204 3694 15260
rect 3694 15204 3750 15260
rect 3750 15204 3754 15260
rect 3690 15200 3754 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 13445 15260 13509 15264
rect 13445 15204 13449 15260
rect 13449 15204 13505 15260
rect 13505 15204 13509 15260
rect 13445 15200 13509 15204
rect 13525 15260 13589 15264
rect 13525 15204 13529 15260
rect 13529 15204 13585 15260
rect 13585 15204 13589 15260
rect 13525 15200 13589 15204
rect 13605 15260 13669 15264
rect 13605 15204 13609 15260
rect 13609 15204 13665 15260
rect 13665 15204 13669 15260
rect 13605 15200 13669 15204
rect 13685 15260 13749 15264
rect 13685 15204 13689 15260
rect 13689 15204 13745 15260
rect 13745 15204 13749 15260
rect 13685 15200 13749 15204
rect 9444 14996 9508 15060
rect 5949 14716 6013 14720
rect 5949 14660 5953 14716
rect 5953 14660 6009 14716
rect 6009 14660 6013 14716
rect 5949 14656 6013 14660
rect 6029 14716 6093 14720
rect 6029 14660 6033 14716
rect 6033 14660 6089 14716
rect 6089 14660 6093 14716
rect 6029 14656 6093 14660
rect 6109 14716 6173 14720
rect 6109 14660 6113 14716
rect 6113 14660 6169 14716
rect 6169 14660 6173 14716
rect 6109 14656 6173 14660
rect 6189 14716 6253 14720
rect 6189 14660 6193 14716
rect 6193 14660 6249 14716
rect 6249 14660 6253 14716
rect 6189 14656 6253 14660
rect 10946 14716 11010 14720
rect 10946 14660 10950 14716
rect 10950 14660 11006 14716
rect 11006 14660 11010 14716
rect 10946 14656 11010 14660
rect 11026 14716 11090 14720
rect 11026 14660 11030 14716
rect 11030 14660 11086 14716
rect 11086 14660 11090 14716
rect 11026 14656 11090 14660
rect 11106 14716 11170 14720
rect 11106 14660 11110 14716
rect 11110 14660 11166 14716
rect 11166 14660 11170 14716
rect 11106 14656 11170 14660
rect 11186 14716 11250 14720
rect 11186 14660 11190 14716
rect 11190 14660 11246 14716
rect 11246 14660 11250 14716
rect 11186 14656 11250 14660
rect 3450 14172 3514 14176
rect 3450 14116 3454 14172
rect 3454 14116 3510 14172
rect 3510 14116 3514 14172
rect 3450 14112 3514 14116
rect 3530 14172 3594 14176
rect 3530 14116 3534 14172
rect 3534 14116 3590 14172
rect 3590 14116 3594 14172
rect 3530 14112 3594 14116
rect 3610 14172 3674 14176
rect 3610 14116 3614 14172
rect 3614 14116 3670 14172
rect 3670 14116 3674 14172
rect 3610 14112 3674 14116
rect 3690 14172 3754 14176
rect 3690 14116 3694 14172
rect 3694 14116 3750 14172
rect 3750 14116 3754 14172
rect 3690 14112 3754 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 13445 14172 13509 14176
rect 13445 14116 13449 14172
rect 13449 14116 13505 14172
rect 13505 14116 13509 14172
rect 13445 14112 13509 14116
rect 13525 14172 13589 14176
rect 13525 14116 13529 14172
rect 13529 14116 13585 14172
rect 13585 14116 13589 14172
rect 13525 14112 13589 14116
rect 13605 14172 13669 14176
rect 13605 14116 13609 14172
rect 13609 14116 13665 14172
rect 13665 14116 13669 14172
rect 13605 14112 13669 14116
rect 13685 14172 13749 14176
rect 13685 14116 13689 14172
rect 13689 14116 13745 14172
rect 13745 14116 13749 14172
rect 13685 14112 13749 14116
rect 5949 13628 6013 13632
rect 5949 13572 5953 13628
rect 5953 13572 6009 13628
rect 6009 13572 6013 13628
rect 5949 13568 6013 13572
rect 6029 13628 6093 13632
rect 6029 13572 6033 13628
rect 6033 13572 6089 13628
rect 6089 13572 6093 13628
rect 6029 13568 6093 13572
rect 6109 13628 6173 13632
rect 6109 13572 6113 13628
rect 6113 13572 6169 13628
rect 6169 13572 6173 13628
rect 6109 13568 6173 13572
rect 6189 13628 6253 13632
rect 6189 13572 6193 13628
rect 6193 13572 6249 13628
rect 6249 13572 6253 13628
rect 6189 13568 6253 13572
rect 10946 13628 11010 13632
rect 10946 13572 10950 13628
rect 10950 13572 11006 13628
rect 11006 13572 11010 13628
rect 10946 13568 11010 13572
rect 11026 13628 11090 13632
rect 11026 13572 11030 13628
rect 11030 13572 11086 13628
rect 11086 13572 11090 13628
rect 11026 13568 11090 13572
rect 11106 13628 11170 13632
rect 11106 13572 11110 13628
rect 11110 13572 11166 13628
rect 11166 13572 11170 13628
rect 11106 13568 11170 13572
rect 11186 13628 11250 13632
rect 11186 13572 11190 13628
rect 11190 13572 11246 13628
rect 11246 13572 11250 13628
rect 11186 13568 11250 13572
rect 3450 13084 3514 13088
rect 3450 13028 3454 13084
rect 3454 13028 3510 13084
rect 3510 13028 3514 13084
rect 3450 13024 3514 13028
rect 3530 13084 3594 13088
rect 3530 13028 3534 13084
rect 3534 13028 3590 13084
rect 3590 13028 3594 13084
rect 3530 13024 3594 13028
rect 3610 13084 3674 13088
rect 3610 13028 3614 13084
rect 3614 13028 3670 13084
rect 3670 13028 3674 13084
rect 3610 13024 3674 13028
rect 3690 13084 3754 13088
rect 3690 13028 3694 13084
rect 3694 13028 3750 13084
rect 3750 13028 3754 13084
rect 3690 13024 3754 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 13445 13084 13509 13088
rect 13445 13028 13449 13084
rect 13449 13028 13505 13084
rect 13505 13028 13509 13084
rect 13445 13024 13509 13028
rect 13525 13084 13589 13088
rect 13525 13028 13529 13084
rect 13529 13028 13585 13084
rect 13585 13028 13589 13084
rect 13525 13024 13589 13028
rect 13605 13084 13669 13088
rect 13605 13028 13609 13084
rect 13609 13028 13665 13084
rect 13665 13028 13669 13084
rect 13605 13024 13669 13028
rect 13685 13084 13749 13088
rect 13685 13028 13689 13084
rect 13689 13028 13745 13084
rect 13745 13028 13749 13084
rect 13685 13024 13749 13028
rect 5949 12540 6013 12544
rect 5949 12484 5953 12540
rect 5953 12484 6009 12540
rect 6009 12484 6013 12540
rect 5949 12480 6013 12484
rect 6029 12540 6093 12544
rect 6029 12484 6033 12540
rect 6033 12484 6089 12540
rect 6089 12484 6093 12540
rect 6029 12480 6093 12484
rect 6109 12540 6173 12544
rect 6109 12484 6113 12540
rect 6113 12484 6169 12540
rect 6169 12484 6173 12540
rect 6109 12480 6173 12484
rect 6189 12540 6253 12544
rect 6189 12484 6193 12540
rect 6193 12484 6249 12540
rect 6249 12484 6253 12540
rect 6189 12480 6253 12484
rect 10946 12540 11010 12544
rect 10946 12484 10950 12540
rect 10950 12484 11006 12540
rect 11006 12484 11010 12540
rect 10946 12480 11010 12484
rect 11026 12540 11090 12544
rect 11026 12484 11030 12540
rect 11030 12484 11086 12540
rect 11086 12484 11090 12540
rect 11026 12480 11090 12484
rect 11106 12540 11170 12544
rect 11106 12484 11110 12540
rect 11110 12484 11166 12540
rect 11166 12484 11170 12540
rect 11106 12480 11170 12484
rect 11186 12540 11250 12544
rect 11186 12484 11190 12540
rect 11190 12484 11246 12540
rect 11246 12484 11250 12540
rect 11186 12480 11250 12484
rect 6500 12276 6564 12340
rect 3450 11996 3514 12000
rect 3450 11940 3454 11996
rect 3454 11940 3510 11996
rect 3510 11940 3514 11996
rect 3450 11936 3514 11940
rect 3530 11996 3594 12000
rect 3530 11940 3534 11996
rect 3534 11940 3590 11996
rect 3590 11940 3594 11996
rect 3530 11936 3594 11940
rect 3610 11996 3674 12000
rect 3610 11940 3614 11996
rect 3614 11940 3670 11996
rect 3670 11940 3674 11996
rect 3610 11936 3674 11940
rect 3690 11996 3754 12000
rect 3690 11940 3694 11996
rect 3694 11940 3750 11996
rect 3750 11940 3754 11996
rect 3690 11936 3754 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 13445 11996 13509 12000
rect 13445 11940 13449 11996
rect 13449 11940 13505 11996
rect 13505 11940 13509 11996
rect 13445 11936 13509 11940
rect 13525 11996 13589 12000
rect 13525 11940 13529 11996
rect 13529 11940 13585 11996
rect 13585 11940 13589 11996
rect 13525 11936 13589 11940
rect 13605 11996 13669 12000
rect 13605 11940 13609 11996
rect 13609 11940 13665 11996
rect 13665 11940 13669 11996
rect 13605 11936 13669 11940
rect 13685 11996 13749 12000
rect 13685 11940 13689 11996
rect 13689 11940 13745 11996
rect 13745 11940 13749 11996
rect 13685 11936 13749 11940
rect 9444 11792 9508 11796
rect 9444 11736 9494 11792
rect 9494 11736 9508 11792
rect 9444 11732 9508 11736
rect 11468 11732 11532 11796
rect 5949 11452 6013 11456
rect 5949 11396 5953 11452
rect 5953 11396 6009 11452
rect 6009 11396 6013 11452
rect 5949 11392 6013 11396
rect 6029 11452 6093 11456
rect 6029 11396 6033 11452
rect 6033 11396 6089 11452
rect 6089 11396 6093 11452
rect 6029 11392 6093 11396
rect 6109 11452 6173 11456
rect 6109 11396 6113 11452
rect 6113 11396 6169 11452
rect 6169 11396 6173 11452
rect 6109 11392 6173 11396
rect 6189 11452 6253 11456
rect 6189 11396 6193 11452
rect 6193 11396 6249 11452
rect 6249 11396 6253 11452
rect 6189 11392 6253 11396
rect 10946 11452 11010 11456
rect 10946 11396 10950 11452
rect 10950 11396 11006 11452
rect 11006 11396 11010 11452
rect 10946 11392 11010 11396
rect 11026 11452 11090 11456
rect 11026 11396 11030 11452
rect 11030 11396 11086 11452
rect 11086 11396 11090 11452
rect 11026 11392 11090 11396
rect 11106 11452 11170 11456
rect 11106 11396 11110 11452
rect 11110 11396 11166 11452
rect 11166 11396 11170 11452
rect 11106 11392 11170 11396
rect 11186 11452 11250 11456
rect 11186 11396 11190 11452
rect 11190 11396 11246 11452
rect 11246 11396 11250 11452
rect 11186 11392 11250 11396
rect 9076 10916 9140 10980
rect 3450 10908 3514 10912
rect 3450 10852 3454 10908
rect 3454 10852 3510 10908
rect 3510 10852 3514 10908
rect 3450 10848 3514 10852
rect 3530 10908 3594 10912
rect 3530 10852 3534 10908
rect 3534 10852 3590 10908
rect 3590 10852 3594 10908
rect 3530 10848 3594 10852
rect 3610 10908 3674 10912
rect 3610 10852 3614 10908
rect 3614 10852 3670 10908
rect 3670 10852 3674 10908
rect 3610 10848 3674 10852
rect 3690 10908 3754 10912
rect 3690 10852 3694 10908
rect 3694 10852 3750 10908
rect 3750 10852 3754 10908
rect 3690 10848 3754 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 13445 10908 13509 10912
rect 13445 10852 13449 10908
rect 13449 10852 13505 10908
rect 13505 10852 13509 10908
rect 13445 10848 13509 10852
rect 13525 10908 13589 10912
rect 13525 10852 13529 10908
rect 13529 10852 13585 10908
rect 13585 10852 13589 10908
rect 13525 10848 13589 10852
rect 13605 10908 13669 10912
rect 13605 10852 13609 10908
rect 13609 10852 13665 10908
rect 13665 10852 13669 10908
rect 13605 10848 13669 10852
rect 13685 10908 13749 10912
rect 13685 10852 13689 10908
rect 13689 10852 13745 10908
rect 13745 10852 13749 10908
rect 13685 10848 13749 10852
rect 5949 10364 6013 10368
rect 5949 10308 5953 10364
rect 5953 10308 6009 10364
rect 6009 10308 6013 10364
rect 5949 10304 6013 10308
rect 6029 10364 6093 10368
rect 6029 10308 6033 10364
rect 6033 10308 6089 10364
rect 6089 10308 6093 10364
rect 6029 10304 6093 10308
rect 6109 10364 6173 10368
rect 6109 10308 6113 10364
rect 6113 10308 6169 10364
rect 6169 10308 6173 10364
rect 6109 10304 6173 10308
rect 6189 10364 6253 10368
rect 6189 10308 6193 10364
rect 6193 10308 6249 10364
rect 6249 10308 6253 10364
rect 6189 10304 6253 10308
rect 10946 10364 11010 10368
rect 10946 10308 10950 10364
rect 10950 10308 11006 10364
rect 11006 10308 11010 10364
rect 10946 10304 11010 10308
rect 11026 10364 11090 10368
rect 11026 10308 11030 10364
rect 11030 10308 11086 10364
rect 11086 10308 11090 10364
rect 11026 10304 11090 10308
rect 11106 10364 11170 10368
rect 11106 10308 11110 10364
rect 11110 10308 11166 10364
rect 11166 10308 11170 10364
rect 11106 10304 11170 10308
rect 11186 10364 11250 10368
rect 11186 10308 11190 10364
rect 11190 10308 11246 10364
rect 11246 10308 11250 10364
rect 11186 10304 11250 10308
rect 3450 9820 3514 9824
rect 3450 9764 3454 9820
rect 3454 9764 3510 9820
rect 3510 9764 3514 9820
rect 3450 9760 3514 9764
rect 3530 9820 3594 9824
rect 3530 9764 3534 9820
rect 3534 9764 3590 9820
rect 3590 9764 3594 9820
rect 3530 9760 3594 9764
rect 3610 9820 3674 9824
rect 3610 9764 3614 9820
rect 3614 9764 3670 9820
rect 3670 9764 3674 9820
rect 3610 9760 3674 9764
rect 3690 9820 3754 9824
rect 3690 9764 3694 9820
rect 3694 9764 3750 9820
rect 3750 9764 3754 9820
rect 3690 9760 3754 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 13445 9820 13509 9824
rect 13445 9764 13449 9820
rect 13449 9764 13505 9820
rect 13505 9764 13509 9820
rect 13445 9760 13509 9764
rect 13525 9820 13589 9824
rect 13525 9764 13529 9820
rect 13529 9764 13585 9820
rect 13585 9764 13589 9820
rect 13525 9760 13589 9764
rect 13605 9820 13669 9824
rect 13605 9764 13609 9820
rect 13609 9764 13665 9820
rect 13665 9764 13669 9820
rect 13605 9760 13669 9764
rect 13685 9820 13749 9824
rect 13685 9764 13689 9820
rect 13689 9764 13745 9820
rect 13745 9764 13749 9820
rect 13685 9760 13749 9764
rect 11652 9556 11716 9620
rect 5949 9276 6013 9280
rect 5949 9220 5953 9276
rect 5953 9220 6009 9276
rect 6009 9220 6013 9276
rect 5949 9216 6013 9220
rect 6029 9276 6093 9280
rect 6029 9220 6033 9276
rect 6033 9220 6089 9276
rect 6089 9220 6093 9276
rect 6029 9216 6093 9220
rect 6109 9276 6173 9280
rect 6109 9220 6113 9276
rect 6113 9220 6169 9276
rect 6169 9220 6173 9276
rect 6109 9216 6173 9220
rect 6189 9276 6253 9280
rect 6189 9220 6193 9276
rect 6193 9220 6249 9276
rect 6249 9220 6253 9276
rect 6189 9216 6253 9220
rect 10946 9276 11010 9280
rect 10946 9220 10950 9276
rect 10950 9220 11006 9276
rect 11006 9220 11010 9276
rect 10946 9216 11010 9220
rect 11026 9276 11090 9280
rect 11026 9220 11030 9276
rect 11030 9220 11086 9276
rect 11086 9220 11090 9276
rect 11026 9216 11090 9220
rect 11106 9276 11170 9280
rect 11106 9220 11110 9276
rect 11110 9220 11166 9276
rect 11166 9220 11170 9276
rect 11106 9216 11170 9220
rect 11186 9276 11250 9280
rect 11186 9220 11190 9276
rect 11190 9220 11246 9276
rect 11246 9220 11250 9276
rect 11186 9216 11250 9220
rect 10364 8876 10428 8940
rect 3450 8732 3514 8736
rect 3450 8676 3454 8732
rect 3454 8676 3510 8732
rect 3510 8676 3514 8732
rect 3450 8672 3514 8676
rect 3530 8732 3594 8736
rect 3530 8676 3534 8732
rect 3534 8676 3590 8732
rect 3590 8676 3594 8732
rect 3530 8672 3594 8676
rect 3610 8732 3674 8736
rect 3610 8676 3614 8732
rect 3614 8676 3670 8732
rect 3670 8676 3674 8732
rect 3610 8672 3674 8676
rect 3690 8732 3754 8736
rect 3690 8676 3694 8732
rect 3694 8676 3750 8732
rect 3750 8676 3754 8732
rect 3690 8672 3754 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 13445 8732 13509 8736
rect 13445 8676 13449 8732
rect 13449 8676 13505 8732
rect 13505 8676 13509 8732
rect 13445 8672 13509 8676
rect 13525 8732 13589 8736
rect 13525 8676 13529 8732
rect 13529 8676 13585 8732
rect 13585 8676 13589 8732
rect 13525 8672 13589 8676
rect 13605 8732 13669 8736
rect 13605 8676 13609 8732
rect 13609 8676 13665 8732
rect 13665 8676 13669 8732
rect 13605 8672 13669 8676
rect 13685 8732 13749 8736
rect 13685 8676 13689 8732
rect 13689 8676 13745 8732
rect 13745 8676 13749 8732
rect 13685 8672 13749 8676
rect 7420 8196 7484 8260
rect 5949 8188 6013 8192
rect 5949 8132 5953 8188
rect 5953 8132 6009 8188
rect 6009 8132 6013 8188
rect 5949 8128 6013 8132
rect 6029 8188 6093 8192
rect 6029 8132 6033 8188
rect 6033 8132 6089 8188
rect 6089 8132 6093 8188
rect 6029 8128 6093 8132
rect 6109 8188 6173 8192
rect 6109 8132 6113 8188
rect 6113 8132 6169 8188
rect 6169 8132 6173 8188
rect 6109 8128 6173 8132
rect 6189 8188 6253 8192
rect 6189 8132 6193 8188
rect 6193 8132 6249 8188
rect 6249 8132 6253 8188
rect 6189 8128 6253 8132
rect 10946 8188 11010 8192
rect 10946 8132 10950 8188
rect 10950 8132 11006 8188
rect 11006 8132 11010 8188
rect 10946 8128 11010 8132
rect 11026 8188 11090 8192
rect 11026 8132 11030 8188
rect 11030 8132 11086 8188
rect 11086 8132 11090 8188
rect 11026 8128 11090 8132
rect 11106 8188 11170 8192
rect 11106 8132 11110 8188
rect 11110 8132 11166 8188
rect 11166 8132 11170 8188
rect 11106 8128 11170 8132
rect 11186 8188 11250 8192
rect 11186 8132 11190 8188
rect 11190 8132 11246 8188
rect 11246 8132 11250 8188
rect 11186 8128 11250 8132
rect 11468 8120 11532 8124
rect 11468 8064 11518 8120
rect 11518 8064 11532 8120
rect 11468 8060 11532 8064
rect 3450 7644 3514 7648
rect 3450 7588 3454 7644
rect 3454 7588 3510 7644
rect 3510 7588 3514 7644
rect 3450 7584 3514 7588
rect 3530 7644 3594 7648
rect 3530 7588 3534 7644
rect 3534 7588 3590 7644
rect 3590 7588 3594 7644
rect 3530 7584 3594 7588
rect 3610 7644 3674 7648
rect 3610 7588 3614 7644
rect 3614 7588 3670 7644
rect 3670 7588 3674 7644
rect 3610 7584 3674 7588
rect 3690 7644 3754 7648
rect 3690 7588 3694 7644
rect 3694 7588 3750 7644
rect 3750 7588 3754 7644
rect 3690 7584 3754 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 13445 7644 13509 7648
rect 13445 7588 13449 7644
rect 13449 7588 13505 7644
rect 13505 7588 13509 7644
rect 13445 7584 13509 7588
rect 13525 7644 13589 7648
rect 13525 7588 13529 7644
rect 13529 7588 13585 7644
rect 13585 7588 13589 7644
rect 13525 7584 13589 7588
rect 13605 7644 13669 7648
rect 13605 7588 13609 7644
rect 13609 7588 13665 7644
rect 13665 7588 13669 7644
rect 13605 7584 13669 7588
rect 13685 7644 13749 7648
rect 13685 7588 13689 7644
rect 13689 7588 13745 7644
rect 13745 7588 13749 7644
rect 13685 7584 13749 7588
rect 5949 7100 6013 7104
rect 5949 7044 5953 7100
rect 5953 7044 6009 7100
rect 6009 7044 6013 7100
rect 5949 7040 6013 7044
rect 6029 7100 6093 7104
rect 6029 7044 6033 7100
rect 6033 7044 6089 7100
rect 6089 7044 6093 7100
rect 6029 7040 6093 7044
rect 6109 7100 6173 7104
rect 6109 7044 6113 7100
rect 6113 7044 6169 7100
rect 6169 7044 6173 7100
rect 6109 7040 6173 7044
rect 6189 7100 6253 7104
rect 6189 7044 6193 7100
rect 6193 7044 6249 7100
rect 6249 7044 6253 7100
rect 6189 7040 6253 7044
rect 10946 7100 11010 7104
rect 10946 7044 10950 7100
rect 10950 7044 11006 7100
rect 11006 7044 11010 7100
rect 10946 7040 11010 7044
rect 11026 7100 11090 7104
rect 11026 7044 11030 7100
rect 11030 7044 11086 7100
rect 11086 7044 11090 7100
rect 11026 7040 11090 7044
rect 11106 7100 11170 7104
rect 11106 7044 11110 7100
rect 11110 7044 11166 7100
rect 11166 7044 11170 7100
rect 11106 7040 11170 7044
rect 11186 7100 11250 7104
rect 11186 7044 11190 7100
rect 11190 7044 11246 7100
rect 11246 7044 11250 7100
rect 11186 7040 11250 7044
rect 3450 6556 3514 6560
rect 3450 6500 3454 6556
rect 3454 6500 3510 6556
rect 3510 6500 3514 6556
rect 3450 6496 3514 6500
rect 3530 6556 3594 6560
rect 3530 6500 3534 6556
rect 3534 6500 3590 6556
rect 3590 6500 3594 6556
rect 3530 6496 3594 6500
rect 3610 6556 3674 6560
rect 3610 6500 3614 6556
rect 3614 6500 3670 6556
rect 3670 6500 3674 6556
rect 3610 6496 3674 6500
rect 3690 6556 3754 6560
rect 3690 6500 3694 6556
rect 3694 6500 3750 6556
rect 3750 6500 3754 6556
rect 3690 6496 3754 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 13445 6556 13509 6560
rect 13445 6500 13449 6556
rect 13449 6500 13505 6556
rect 13505 6500 13509 6556
rect 13445 6496 13509 6500
rect 13525 6556 13589 6560
rect 13525 6500 13529 6556
rect 13529 6500 13585 6556
rect 13585 6500 13589 6556
rect 13525 6496 13589 6500
rect 13605 6556 13669 6560
rect 13605 6500 13609 6556
rect 13609 6500 13665 6556
rect 13665 6500 13669 6556
rect 13605 6496 13669 6500
rect 13685 6556 13749 6560
rect 13685 6500 13689 6556
rect 13689 6500 13745 6556
rect 13745 6500 13749 6556
rect 13685 6496 13749 6500
rect 11468 6156 11532 6220
rect 5949 6012 6013 6016
rect 5949 5956 5953 6012
rect 5953 5956 6009 6012
rect 6009 5956 6013 6012
rect 5949 5952 6013 5956
rect 6029 6012 6093 6016
rect 6029 5956 6033 6012
rect 6033 5956 6089 6012
rect 6089 5956 6093 6012
rect 6029 5952 6093 5956
rect 6109 6012 6173 6016
rect 6109 5956 6113 6012
rect 6113 5956 6169 6012
rect 6169 5956 6173 6012
rect 6109 5952 6173 5956
rect 6189 6012 6253 6016
rect 6189 5956 6193 6012
rect 6193 5956 6249 6012
rect 6249 5956 6253 6012
rect 6189 5952 6253 5956
rect 10946 6012 11010 6016
rect 10946 5956 10950 6012
rect 10950 5956 11006 6012
rect 11006 5956 11010 6012
rect 10946 5952 11010 5956
rect 11026 6012 11090 6016
rect 11026 5956 11030 6012
rect 11030 5956 11086 6012
rect 11086 5956 11090 6012
rect 11026 5952 11090 5956
rect 11106 6012 11170 6016
rect 11106 5956 11110 6012
rect 11110 5956 11166 6012
rect 11166 5956 11170 6012
rect 11106 5952 11170 5956
rect 11186 6012 11250 6016
rect 11186 5956 11190 6012
rect 11190 5956 11246 6012
rect 11246 5956 11250 6012
rect 11186 5952 11250 5956
rect 3450 5468 3514 5472
rect 3450 5412 3454 5468
rect 3454 5412 3510 5468
rect 3510 5412 3514 5468
rect 3450 5408 3514 5412
rect 3530 5468 3594 5472
rect 3530 5412 3534 5468
rect 3534 5412 3590 5468
rect 3590 5412 3594 5468
rect 3530 5408 3594 5412
rect 3610 5468 3674 5472
rect 3610 5412 3614 5468
rect 3614 5412 3670 5468
rect 3670 5412 3674 5468
rect 3610 5408 3674 5412
rect 3690 5468 3754 5472
rect 3690 5412 3694 5468
rect 3694 5412 3750 5468
rect 3750 5412 3754 5468
rect 3690 5408 3754 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 13445 5468 13509 5472
rect 13445 5412 13449 5468
rect 13449 5412 13505 5468
rect 13505 5412 13509 5468
rect 13445 5408 13509 5412
rect 13525 5468 13589 5472
rect 13525 5412 13529 5468
rect 13529 5412 13585 5468
rect 13585 5412 13589 5468
rect 13525 5408 13589 5412
rect 13605 5468 13669 5472
rect 13605 5412 13609 5468
rect 13609 5412 13665 5468
rect 13665 5412 13669 5468
rect 13605 5408 13669 5412
rect 13685 5468 13749 5472
rect 13685 5412 13689 5468
rect 13689 5412 13745 5468
rect 13745 5412 13749 5468
rect 13685 5408 13749 5412
rect 5949 4924 6013 4928
rect 5949 4868 5953 4924
rect 5953 4868 6009 4924
rect 6009 4868 6013 4924
rect 5949 4864 6013 4868
rect 6029 4924 6093 4928
rect 6029 4868 6033 4924
rect 6033 4868 6089 4924
rect 6089 4868 6093 4924
rect 6029 4864 6093 4868
rect 6109 4924 6173 4928
rect 6109 4868 6113 4924
rect 6113 4868 6169 4924
rect 6169 4868 6173 4924
rect 6109 4864 6173 4868
rect 6189 4924 6253 4928
rect 6189 4868 6193 4924
rect 6193 4868 6249 4924
rect 6249 4868 6253 4924
rect 6189 4864 6253 4868
rect 10946 4924 11010 4928
rect 10946 4868 10950 4924
rect 10950 4868 11006 4924
rect 11006 4868 11010 4924
rect 10946 4864 11010 4868
rect 11026 4924 11090 4928
rect 11026 4868 11030 4924
rect 11030 4868 11086 4924
rect 11086 4868 11090 4924
rect 11026 4864 11090 4868
rect 11106 4924 11170 4928
rect 11106 4868 11110 4924
rect 11110 4868 11166 4924
rect 11166 4868 11170 4924
rect 11106 4864 11170 4868
rect 11186 4924 11250 4928
rect 11186 4868 11190 4924
rect 11190 4868 11246 4924
rect 11246 4868 11250 4924
rect 11186 4864 11250 4868
rect 3450 4380 3514 4384
rect 3450 4324 3454 4380
rect 3454 4324 3510 4380
rect 3510 4324 3514 4380
rect 3450 4320 3514 4324
rect 3530 4380 3594 4384
rect 3530 4324 3534 4380
rect 3534 4324 3590 4380
rect 3590 4324 3594 4380
rect 3530 4320 3594 4324
rect 3610 4380 3674 4384
rect 3610 4324 3614 4380
rect 3614 4324 3670 4380
rect 3670 4324 3674 4380
rect 3610 4320 3674 4324
rect 3690 4380 3754 4384
rect 3690 4324 3694 4380
rect 3694 4324 3750 4380
rect 3750 4324 3754 4380
rect 3690 4320 3754 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 13445 4380 13509 4384
rect 13445 4324 13449 4380
rect 13449 4324 13505 4380
rect 13505 4324 13509 4380
rect 13445 4320 13509 4324
rect 13525 4380 13589 4384
rect 13525 4324 13529 4380
rect 13529 4324 13585 4380
rect 13585 4324 13589 4380
rect 13525 4320 13589 4324
rect 13605 4380 13669 4384
rect 13605 4324 13609 4380
rect 13609 4324 13665 4380
rect 13665 4324 13669 4380
rect 13605 4320 13669 4324
rect 13685 4380 13749 4384
rect 13685 4324 13689 4380
rect 13689 4324 13745 4380
rect 13745 4324 13749 4380
rect 13685 4320 13749 4324
rect 5949 3836 6013 3840
rect 5949 3780 5953 3836
rect 5953 3780 6009 3836
rect 6009 3780 6013 3836
rect 5949 3776 6013 3780
rect 6029 3836 6093 3840
rect 6029 3780 6033 3836
rect 6033 3780 6089 3836
rect 6089 3780 6093 3836
rect 6029 3776 6093 3780
rect 6109 3836 6173 3840
rect 6109 3780 6113 3836
rect 6113 3780 6169 3836
rect 6169 3780 6173 3836
rect 6109 3776 6173 3780
rect 6189 3836 6253 3840
rect 6189 3780 6193 3836
rect 6193 3780 6249 3836
rect 6249 3780 6253 3836
rect 6189 3776 6253 3780
rect 10946 3836 11010 3840
rect 10946 3780 10950 3836
rect 10950 3780 11006 3836
rect 11006 3780 11010 3836
rect 10946 3776 11010 3780
rect 11026 3836 11090 3840
rect 11026 3780 11030 3836
rect 11030 3780 11086 3836
rect 11086 3780 11090 3836
rect 11026 3776 11090 3780
rect 11106 3836 11170 3840
rect 11106 3780 11110 3836
rect 11110 3780 11166 3836
rect 11166 3780 11170 3836
rect 11106 3776 11170 3780
rect 11186 3836 11250 3840
rect 11186 3780 11190 3836
rect 11190 3780 11246 3836
rect 11246 3780 11250 3836
rect 11186 3776 11250 3780
rect 3450 3292 3514 3296
rect 3450 3236 3454 3292
rect 3454 3236 3510 3292
rect 3510 3236 3514 3292
rect 3450 3232 3514 3236
rect 3530 3292 3594 3296
rect 3530 3236 3534 3292
rect 3534 3236 3590 3292
rect 3590 3236 3594 3292
rect 3530 3232 3594 3236
rect 3610 3292 3674 3296
rect 3610 3236 3614 3292
rect 3614 3236 3670 3292
rect 3670 3236 3674 3292
rect 3610 3232 3674 3236
rect 3690 3292 3754 3296
rect 3690 3236 3694 3292
rect 3694 3236 3750 3292
rect 3750 3236 3754 3292
rect 3690 3232 3754 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 13445 3292 13509 3296
rect 13445 3236 13449 3292
rect 13449 3236 13505 3292
rect 13505 3236 13509 3292
rect 13445 3232 13509 3236
rect 13525 3292 13589 3296
rect 13525 3236 13529 3292
rect 13529 3236 13585 3292
rect 13585 3236 13589 3292
rect 13525 3232 13589 3236
rect 13605 3292 13669 3296
rect 13605 3236 13609 3292
rect 13609 3236 13665 3292
rect 13665 3236 13669 3292
rect 13605 3232 13669 3236
rect 13685 3292 13749 3296
rect 13685 3236 13689 3292
rect 13689 3236 13745 3292
rect 13745 3236 13749 3292
rect 13685 3232 13749 3236
rect 5949 2748 6013 2752
rect 5949 2692 5953 2748
rect 5953 2692 6009 2748
rect 6009 2692 6013 2748
rect 5949 2688 6013 2692
rect 6029 2748 6093 2752
rect 6029 2692 6033 2748
rect 6033 2692 6089 2748
rect 6089 2692 6093 2748
rect 6029 2688 6093 2692
rect 6109 2748 6173 2752
rect 6109 2692 6113 2748
rect 6113 2692 6169 2748
rect 6169 2692 6173 2748
rect 6109 2688 6173 2692
rect 6189 2748 6253 2752
rect 6189 2692 6193 2748
rect 6193 2692 6249 2748
rect 6249 2692 6253 2748
rect 6189 2688 6253 2692
rect 10946 2748 11010 2752
rect 10946 2692 10950 2748
rect 10950 2692 11006 2748
rect 11006 2692 11010 2748
rect 10946 2688 11010 2692
rect 11026 2748 11090 2752
rect 11026 2692 11030 2748
rect 11030 2692 11086 2748
rect 11086 2692 11090 2748
rect 11026 2688 11090 2692
rect 11106 2748 11170 2752
rect 11106 2692 11110 2748
rect 11110 2692 11166 2748
rect 11166 2692 11170 2748
rect 11106 2688 11170 2692
rect 11186 2748 11250 2752
rect 11186 2692 11190 2748
rect 11190 2692 11246 2748
rect 11246 2692 11250 2748
rect 11186 2688 11250 2692
rect 11652 2348 11716 2412
rect 3450 2204 3514 2208
rect 3450 2148 3454 2204
rect 3454 2148 3510 2204
rect 3510 2148 3514 2204
rect 3450 2144 3514 2148
rect 3530 2204 3594 2208
rect 3530 2148 3534 2204
rect 3534 2148 3590 2204
rect 3590 2148 3594 2204
rect 3530 2144 3594 2148
rect 3610 2204 3674 2208
rect 3610 2148 3614 2204
rect 3614 2148 3670 2204
rect 3670 2148 3674 2204
rect 3610 2144 3674 2148
rect 3690 2204 3754 2208
rect 3690 2148 3694 2204
rect 3694 2148 3750 2204
rect 3750 2148 3754 2204
rect 3690 2144 3754 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 13445 2204 13509 2208
rect 13445 2148 13449 2204
rect 13449 2148 13505 2204
rect 13505 2148 13509 2204
rect 13445 2144 13509 2148
rect 13525 2204 13589 2208
rect 13525 2148 13529 2204
rect 13529 2148 13585 2204
rect 13585 2148 13589 2204
rect 13525 2144 13589 2148
rect 13605 2204 13669 2208
rect 13605 2148 13609 2204
rect 13609 2148 13665 2204
rect 13665 2148 13669 2204
rect 13605 2144 13669 2148
rect 13685 2204 13749 2208
rect 13685 2148 13689 2204
rect 13689 2148 13745 2204
rect 13745 2148 13749 2204
rect 13685 2144 13749 2148
rect 10364 852 10428 916
<< metal4 >>
rect 3442 17440 3763 17456
rect 3442 17376 3450 17440
rect 3514 17376 3530 17440
rect 3594 17376 3610 17440
rect 3674 17376 3690 17440
rect 3754 17376 3763 17440
rect 3442 16352 3763 17376
rect 3442 16288 3450 16352
rect 3514 16288 3530 16352
rect 3594 16288 3610 16352
rect 3674 16288 3690 16352
rect 3754 16288 3763 16352
rect 3442 15264 3763 16288
rect 3442 15200 3450 15264
rect 3514 15200 3530 15264
rect 3594 15200 3610 15264
rect 3674 15200 3690 15264
rect 3754 15200 3763 15264
rect 3442 14176 3763 15200
rect 3442 14112 3450 14176
rect 3514 14112 3530 14176
rect 3594 14112 3610 14176
rect 3674 14112 3690 14176
rect 3754 14112 3763 14176
rect 3442 13088 3763 14112
rect 3442 13024 3450 13088
rect 3514 13024 3530 13088
rect 3594 13024 3610 13088
rect 3674 13024 3690 13088
rect 3754 13024 3763 13088
rect 3442 12000 3763 13024
rect 3442 11936 3450 12000
rect 3514 11936 3530 12000
rect 3594 11936 3610 12000
rect 3674 11936 3690 12000
rect 3754 11936 3763 12000
rect 3442 10912 3763 11936
rect 3442 10848 3450 10912
rect 3514 10848 3530 10912
rect 3594 10848 3610 10912
rect 3674 10848 3690 10912
rect 3754 10848 3763 10912
rect 3442 9824 3763 10848
rect 3442 9760 3450 9824
rect 3514 9760 3530 9824
rect 3594 9760 3610 9824
rect 3674 9760 3690 9824
rect 3754 9760 3763 9824
rect 3442 8736 3763 9760
rect 3442 8672 3450 8736
rect 3514 8672 3530 8736
rect 3594 8672 3610 8736
rect 3674 8672 3690 8736
rect 3754 8672 3763 8736
rect 3442 7648 3763 8672
rect 3442 7584 3450 7648
rect 3514 7584 3530 7648
rect 3594 7584 3610 7648
rect 3674 7584 3690 7648
rect 3754 7584 3763 7648
rect 3442 6560 3763 7584
rect 3442 6496 3450 6560
rect 3514 6496 3530 6560
rect 3594 6496 3610 6560
rect 3674 6496 3690 6560
rect 3754 6496 3763 6560
rect 3442 5472 3763 6496
rect 3442 5408 3450 5472
rect 3514 5408 3530 5472
rect 3594 5408 3610 5472
rect 3674 5408 3690 5472
rect 3754 5408 3763 5472
rect 3442 4384 3763 5408
rect 3442 4320 3450 4384
rect 3514 4320 3530 4384
rect 3594 4320 3610 4384
rect 3674 4320 3690 4384
rect 3754 4320 3763 4384
rect 3442 3296 3763 4320
rect 3442 3232 3450 3296
rect 3514 3232 3530 3296
rect 3594 3232 3610 3296
rect 3674 3232 3690 3296
rect 3754 3232 3763 3296
rect 3442 2208 3763 3232
rect 3442 2144 3450 2208
rect 3514 2144 3530 2208
rect 3594 2144 3610 2208
rect 3674 2144 3690 2208
rect 3754 2144 3763 2208
rect 3442 2128 3763 2144
rect 5941 16896 6261 17456
rect 5941 16832 5949 16896
rect 6013 16832 6029 16896
rect 6093 16832 6109 16896
rect 6173 16832 6189 16896
rect 6253 16832 6261 16896
rect 5941 15808 6261 16832
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 9075 16964 9141 16965
rect 9075 16900 9076 16964
rect 9140 16900 9141 16964
rect 9075 16899 9141 16900
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 7419 15876 7485 15877
rect 7419 15812 7420 15876
rect 7484 15812 7485 15876
rect 7419 15811 7485 15812
rect 5941 15744 5949 15808
rect 6013 15744 6029 15808
rect 6093 15744 6109 15808
rect 6173 15744 6189 15808
rect 6253 15744 6261 15808
rect 5941 14720 6261 15744
rect 6499 15604 6565 15605
rect 6499 15540 6500 15604
rect 6564 15540 6565 15604
rect 6499 15539 6565 15540
rect 5941 14656 5949 14720
rect 6013 14656 6029 14720
rect 6093 14656 6109 14720
rect 6173 14656 6189 14720
rect 6253 14656 6261 14720
rect 5941 13632 6261 14656
rect 5941 13568 5949 13632
rect 6013 13568 6029 13632
rect 6093 13568 6109 13632
rect 6173 13568 6189 13632
rect 6253 13568 6261 13632
rect 5941 12544 6261 13568
rect 5941 12480 5949 12544
rect 6013 12480 6029 12544
rect 6093 12480 6109 12544
rect 6173 12480 6189 12544
rect 6253 12480 6261 12544
rect 5941 11456 6261 12480
rect 6502 12341 6562 15539
rect 7422 15469 7482 15811
rect 7419 15468 7485 15469
rect 7419 15404 7420 15468
rect 7484 15404 7485 15468
rect 7419 15403 7485 15404
rect 6499 12340 6565 12341
rect 6499 12276 6500 12340
rect 6564 12276 6565 12340
rect 6499 12275 6565 12276
rect 5941 11392 5949 11456
rect 6013 11392 6029 11456
rect 6093 11392 6109 11456
rect 6173 11392 6189 11456
rect 6253 11392 6261 11456
rect 5941 10368 6261 11392
rect 5941 10304 5949 10368
rect 6013 10304 6029 10368
rect 6093 10304 6109 10368
rect 6173 10304 6189 10368
rect 6253 10304 6261 10368
rect 5941 9280 6261 10304
rect 5941 9216 5949 9280
rect 6013 9216 6029 9280
rect 6093 9216 6109 9280
rect 6173 9216 6189 9280
rect 6253 9216 6261 9280
rect 5941 8192 6261 9216
rect 7422 8261 7482 15403
rect 8440 15264 8760 16288
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 9078 10981 9138 16899
rect 10938 16896 11259 17456
rect 13437 17440 13757 17456
rect 13437 17376 13445 17440
rect 13509 17376 13525 17440
rect 13589 17376 13605 17440
rect 13669 17376 13685 17440
rect 13749 17376 13757 17440
rect 11467 17100 11533 17101
rect 11467 17036 11468 17100
rect 11532 17036 11533 17100
rect 11467 17035 11533 17036
rect 10938 16832 10946 16896
rect 11010 16832 11026 16896
rect 11090 16832 11106 16896
rect 11170 16832 11186 16896
rect 11250 16832 11259 16896
rect 10938 15808 11259 16832
rect 10938 15744 10946 15808
rect 11010 15744 11026 15808
rect 11090 15744 11106 15808
rect 11170 15744 11186 15808
rect 11250 15744 11259 15808
rect 9443 15060 9509 15061
rect 9443 14996 9444 15060
rect 9508 14996 9509 15060
rect 9443 14995 9509 14996
rect 9446 11797 9506 14995
rect 10938 14720 11259 15744
rect 11470 15605 11530 17035
rect 13437 16352 13757 17376
rect 13437 16288 13445 16352
rect 13509 16288 13525 16352
rect 13589 16288 13605 16352
rect 13669 16288 13685 16352
rect 13749 16288 13757 16352
rect 11467 15604 11533 15605
rect 11467 15540 11468 15604
rect 11532 15540 11533 15604
rect 11467 15539 11533 15540
rect 10938 14656 10946 14720
rect 11010 14656 11026 14720
rect 11090 14656 11106 14720
rect 11170 14656 11186 14720
rect 11250 14656 11259 14720
rect 10938 13632 11259 14656
rect 10938 13568 10946 13632
rect 11010 13568 11026 13632
rect 11090 13568 11106 13632
rect 11170 13568 11186 13632
rect 11250 13568 11259 13632
rect 10938 12544 11259 13568
rect 10938 12480 10946 12544
rect 11010 12480 11026 12544
rect 11090 12480 11106 12544
rect 11170 12480 11186 12544
rect 11250 12480 11259 12544
rect 9443 11796 9509 11797
rect 9443 11732 9444 11796
rect 9508 11732 9509 11796
rect 9443 11731 9509 11732
rect 10938 11456 11259 12480
rect 11470 11797 11530 15539
rect 13437 15264 13757 16288
rect 13437 15200 13445 15264
rect 13509 15200 13525 15264
rect 13589 15200 13605 15264
rect 13669 15200 13685 15264
rect 13749 15200 13757 15264
rect 13437 14176 13757 15200
rect 13437 14112 13445 14176
rect 13509 14112 13525 14176
rect 13589 14112 13605 14176
rect 13669 14112 13685 14176
rect 13749 14112 13757 14176
rect 13437 13088 13757 14112
rect 13437 13024 13445 13088
rect 13509 13024 13525 13088
rect 13589 13024 13605 13088
rect 13669 13024 13685 13088
rect 13749 13024 13757 13088
rect 13437 12000 13757 13024
rect 13437 11936 13445 12000
rect 13509 11936 13525 12000
rect 13589 11936 13605 12000
rect 13669 11936 13685 12000
rect 13749 11936 13757 12000
rect 11467 11796 11533 11797
rect 11467 11732 11468 11796
rect 11532 11732 11533 11796
rect 11467 11731 11533 11732
rect 10938 11392 10946 11456
rect 11010 11392 11026 11456
rect 11090 11392 11106 11456
rect 11170 11392 11186 11456
rect 11250 11392 11259 11456
rect 9075 10980 9141 10981
rect 9075 10916 9076 10980
rect 9140 10916 9141 10980
rect 9075 10915 9141 10916
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 10938 10368 11259 11392
rect 10938 10304 10946 10368
rect 11010 10304 11026 10368
rect 11090 10304 11106 10368
rect 11170 10304 11186 10368
rect 11250 10304 11259 10368
rect 10938 9280 11259 10304
rect 13437 10912 13757 11936
rect 13437 10848 13445 10912
rect 13509 10848 13525 10912
rect 13589 10848 13605 10912
rect 13669 10848 13685 10912
rect 13749 10848 13757 10912
rect 13437 9824 13757 10848
rect 13437 9760 13445 9824
rect 13509 9760 13525 9824
rect 13589 9760 13605 9824
rect 13669 9760 13685 9824
rect 13749 9760 13757 9824
rect 11651 9620 11717 9621
rect 11651 9556 11652 9620
rect 11716 9556 11717 9620
rect 11651 9555 11717 9556
rect 10938 9216 10946 9280
rect 11010 9216 11026 9280
rect 11090 9216 11106 9280
rect 11170 9216 11186 9280
rect 11250 9216 11259 9280
rect 10363 8940 10429 8941
rect 10363 8876 10364 8940
rect 10428 8876 10429 8940
rect 10363 8875 10429 8876
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 7419 8260 7485 8261
rect 7419 8196 7420 8260
rect 7484 8196 7485 8260
rect 7419 8195 7485 8196
rect 5941 8128 5949 8192
rect 6013 8128 6029 8192
rect 6093 8128 6109 8192
rect 6173 8128 6189 8192
rect 6253 8128 6261 8192
rect 5941 7104 6261 8128
rect 5941 7040 5949 7104
rect 6013 7040 6029 7104
rect 6093 7040 6109 7104
rect 6173 7040 6189 7104
rect 6253 7040 6261 7104
rect 5941 6016 6261 7040
rect 5941 5952 5949 6016
rect 6013 5952 6029 6016
rect 6093 5952 6109 6016
rect 6173 5952 6189 6016
rect 6253 5952 6261 6016
rect 5941 4928 6261 5952
rect 5941 4864 5949 4928
rect 6013 4864 6029 4928
rect 6093 4864 6109 4928
rect 6173 4864 6189 4928
rect 6253 4864 6261 4928
rect 5941 3840 6261 4864
rect 5941 3776 5949 3840
rect 6013 3776 6029 3840
rect 6093 3776 6109 3840
rect 6173 3776 6189 3840
rect 6253 3776 6261 3840
rect 5941 2752 6261 3776
rect 5941 2688 5949 2752
rect 6013 2688 6029 2752
rect 6093 2688 6109 2752
rect 6173 2688 6189 2752
rect 6253 2688 6261 2752
rect 5941 2128 6261 2688
rect 8440 7648 8760 8672
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 2208 8760 3232
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 10366 917 10426 8875
rect 10938 8192 11259 9216
rect 10938 8128 10946 8192
rect 11010 8128 11026 8192
rect 11090 8128 11106 8192
rect 11170 8128 11186 8192
rect 11250 8128 11259 8192
rect 10938 7104 11259 8128
rect 11467 8124 11533 8125
rect 11467 8060 11468 8124
rect 11532 8060 11533 8124
rect 11467 8059 11533 8060
rect 10938 7040 10946 7104
rect 11010 7040 11026 7104
rect 11090 7040 11106 7104
rect 11170 7040 11186 7104
rect 11250 7040 11259 7104
rect 10938 6016 11259 7040
rect 11470 6221 11530 8059
rect 11467 6220 11533 6221
rect 11467 6156 11468 6220
rect 11532 6156 11533 6220
rect 11467 6155 11533 6156
rect 10938 5952 10946 6016
rect 11010 5952 11026 6016
rect 11090 5952 11106 6016
rect 11170 5952 11186 6016
rect 11250 5952 11259 6016
rect 10938 4928 11259 5952
rect 10938 4864 10946 4928
rect 11010 4864 11026 4928
rect 11090 4864 11106 4928
rect 11170 4864 11186 4928
rect 11250 4864 11259 4928
rect 10938 3840 11259 4864
rect 10938 3776 10946 3840
rect 11010 3776 11026 3840
rect 11090 3776 11106 3840
rect 11170 3776 11186 3840
rect 11250 3776 11259 3840
rect 10938 2752 11259 3776
rect 10938 2688 10946 2752
rect 11010 2688 11026 2752
rect 11090 2688 11106 2752
rect 11170 2688 11186 2752
rect 11250 2688 11259 2752
rect 10938 2128 11259 2688
rect 11654 2413 11714 9555
rect 13437 8736 13757 9760
rect 13437 8672 13445 8736
rect 13509 8672 13525 8736
rect 13589 8672 13605 8736
rect 13669 8672 13685 8736
rect 13749 8672 13757 8736
rect 13437 7648 13757 8672
rect 13437 7584 13445 7648
rect 13509 7584 13525 7648
rect 13589 7584 13605 7648
rect 13669 7584 13685 7648
rect 13749 7584 13757 7648
rect 13437 6560 13757 7584
rect 13437 6496 13445 6560
rect 13509 6496 13525 6560
rect 13589 6496 13605 6560
rect 13669 6496 13685 6560
rect 13749 6496 13757 6560
rect 13437 5472 13757 6496
rect 13437 5408 13445 5472
rect 13509 5408 13525 5472
rect 13589 5408 13605 5472
rect 13669 5408 13685 5472
rect 13749 5408 13757 5472
rect 13437 4384 13757 5408
rect 13437 4320 13445 4384
rect 13509 4320 13525 4384
rect 13589 4320 13605 4384
rect 13669 4320 13685 4384
rect 13749 4320 13757 4384
rect 13437 3296 13757 4320
rect 13437 3232 13445 3296
rect 13509 3232 13525 3296
rect 13589 3232 13605 3296
rect 13669 3232 13685 3296
rect 13749 3232 13757 3296
rect 11651 2412 11717 2413
rect 11651 2348 11652 2412
rect 11716 2348 11717 2412
rect 11651 2347 11717 2348
rect 13437 2208 13757 3232
rect 13437 2144 13445 2208
rect 13509 2144 13525 2208
rect 13589 2144 13605 2208
rect 13669 2144 13685 2208
rect 13749 2144 13757 2208
rect 13437 2128 13757 2144
rect 10363 916 10429 917
rect 10363 852 10364 916
rect 10428 852 10429 916
rect 10363 851 10429 852
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1564 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _37_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608910539
transform 1 0 2300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1608910539
transform 1 0 1932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1608910539
transform 1 0 1564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21
timestamp 1608910539
transform 1 0 3036 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4508 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3036 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1608910539
transform 1 0 4876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608910539
transform 1 0 3496 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1608910539
transform 1 0 3128 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 5336 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1608910539
transform 1 0 5612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1608910539
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1608910539
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6532 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1608910539
transform 1 0 6164 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608910539
transform 1 0 6164 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1608910539
transform 1 0 7728 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1608910539
transform 1 0 8556 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8280 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_87
timestamp 1608910539
transform 1 0 9108 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9384 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1608910539
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1608910539
transform 1 0 10212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608910539
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _28_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_106
timestamp 1608910539
transform 1 0 10856 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10948 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1608910539
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1608910539
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_142
timestamp 1608910539
transform 1 0 14168 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_134 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 13432 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_133
timestamp 1608910539
transform 1 0 13340 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1608910539
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1608910539
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_S_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14260 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1608910539
transform 1 0 14076 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_S_FTB01
timestamp 1608910539
transform 1 0 14812 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_S_FTB01
timestamp 1608910539
transform 1 0 14628 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_158
timestamp 1608910539
transform 1 0 15640 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_S_FTB01_A
timestamp 1608910539
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_S_FTB01_A
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_S_FTB01_A
timestamp 1608910539
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_S_FTB01_A
timestamp 1608910539
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 16008 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 16008 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_16
timestamp 1608910539
transform 1 0 2576 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1608910539
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1608910539
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1608910539
transform 1 0 2392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1608910539
transform 1 0 2024 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1608910539
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1608910539
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 4416 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1608910539
transform 1 0 3036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5612 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608910539
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7084 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 8096 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_103
timestamp 1608910539
transform 1 0 10580 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1608910539
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10672 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 11500 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1608910539
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_158
timestamp 1608910539
transform 1 0 15640 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1608910539
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1608910539
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2392 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1608910539
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3404 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4416 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608910539
transform 1 0 5520 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1608910539
transform 1 0 5244 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_71
timestamp 1608910539
transform 1 0 7636 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1608910539
transform 1 0 8556 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7728 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1608910539
transform 1 0 9936 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_3_116 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11776 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_144
timestamp 1608910539
transform 1 0 14352 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_132
timestamp 1608910539
transform 1 0 13248 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_156
timestamp 1608910539
transform 1 0 15456 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 16008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1608910539
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1608910539
transform 1 0 2944 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_32
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 4140 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 3128 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4324 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_53
timestamp 1608910539
transform 1 0 5980 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6624 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 5152 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608910539
transform 1 0 6072 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7912 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8740 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608910539
transform 1 0 7452 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_100
timestamp 1608910539
transform 1 0 10304 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10120 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9936 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_right_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10396 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_110
timestamp 1608910539
transform 1 0 11224 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11316 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_4_140
timestamp 1608910539
transform 1 0 13984 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 13616 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1608910539
transform 1 0 12788 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_158
timestamp 1608910539
transform 1 0 15640 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1608910539
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 16008 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_16
timestamp 1608910539
transform 1 0 2576 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2852 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_38
timestamp 1608910539
transform 1 0 4600 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 4692 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1608910539
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1608910539
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_80
timestamp 1608910539
transform 1 0 8464 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 8280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8556 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 10028 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_5_121
timestamp 1608910539
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1608910539
transform 1 0 11500 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1608910539
transform 1 0 13708 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608910539
transform 1 0 13248 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_157 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1608910539
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 16008 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1608910539
transform 1 0 14996 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_10
timestamp 1608910539
transform 1 0 2024 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp 1608910539
transform 1 0 1932 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2024 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_6_28
timestamp 1608910539
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1608910539
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4600 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3128 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1608910539
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_56
timestamp 1608910539
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_45
timestamp 1608910539
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1608910539
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5428 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_6_63
timestamp 1608910539
transform 1 0 6900 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 6992 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7820 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 8372 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8648 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1608910539
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9200 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_6_101
timestamp 1608910539
transform 1 0 10396 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10212 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10488 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_116
timestamp 1608910539
transform 1 0 11776 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_108
timestamp 1608910539
transform 1 0 11040 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_118
timestamp 1608910539
transform 1 0 11960 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1608910539
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1608910539
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_142
timestamp 1608910539
transform 1 0 14168 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_130
timestamp 1608910539
transform 1 0 13064 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1608910539
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_158
timestamp 1608910539
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp 1608910539
transform 1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 16008 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_10
timestamp 1608910539
transform 1 0 2024 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2116 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2944 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 6532 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5520 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6716 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_77
timestamp 1608910539
transform 1 0 8188 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 8464 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9752 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1608910539
transform 1 0 12420 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1608910539
transform 1 0 11592 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_8_138
timestamp 1608910539
transform 1 0 13800 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_158
timestamp 1608910539
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp 1608910539
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 16008 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_16
timestamp 1608910539
transform 1 0 2576 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_10
timestamp 1608910539
transform 1 0 2024 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 2668 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_26
timestamp 1608910539
transform 1 0 3496 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1608910539
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1608910539
transform 1 0 3864 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1608910539
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_50
timestamp 1608910539
transform 1 0 5704 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 5796 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7636 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9108 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1608910539
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1608910539
transform 1 0 11408 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1608910539
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1608910539
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 16008 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_5
timestamp 1608910539
transform 1 0 1564 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1932 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_10_25
timestamp 1608910539
transform 1 0 3404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1608910539
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 6348 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5520 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 6624 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1608910539
transform 1 0 8096 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_97
timestamp 1608910539
transform 1 0 10028 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1608910539
transform 1 0 10304 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1608910539
transform 1 0 8924 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_109
timestamp 1608910539
transform 1 0 11132 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 11224 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_142
timestamp 1608910539
transform 1 0 14168 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12696 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1608910539
transform 1 0 15640 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_150
timestamp 1608910539
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_15
timestamp 1608910539
transform 1 0 2484 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_40
timestamp 1608910539
transform 1 0 4784 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 4508 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 3036 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5060 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1608910539
transform 1 0 8648 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1608910539
transform 1 0 7820 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6992 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 10304 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1608910539
transform 1 0 9476 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10948 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_11_134
timestamp 1608910539
transform 1 0 13432 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_158
timestamp 1608910539
transform 1 0 15640 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_146
timestamp 1608910539
transform 1 0 14536 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 16008 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 1472 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1608910539
transform 1 0 2300 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1608910539
transform 1 0 4692 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_57
timestamp 1608910539
transform 1 0 6348 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 6440 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5520 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7268 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 8096 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_96
timestamp 1608910539
transform 1 0 9936 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10028 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10856 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 11684 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_143
timestamp 1608910539
transform 1 0 14260 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_131
timestamp 1608910539
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_158
timestamp 1608910539
transform 1 0 15640 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1608910539
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1564 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2024 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_21
timestamp 1608910539
transform 1 0 3036 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4232 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 3496 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1608910539
transform 1 0 4232 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_45
timestamp 1608910539
transform 1 0 5244 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608910539
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5060 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 5336 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1608910539
transform 1 0 6992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 7084 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1608910539
transform 1 0 8464 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_14_93
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1608910539
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1608910539
transform 1 0 8924 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_99
timestamp 1608910539
transform 1 0 10212 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10028 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 10304 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_14_116
timestamp 1608910539
transform 1 0 11776 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1608910539
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 11868 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1608910539
transform 1 0 12144 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10856 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_144
timestamp 1608910539
transform 1 0 14352 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1608910539
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1608910539
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1608910539
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1608910539
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_E_FTB01_A
timestamp 1608910539
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  Test_en_E_FTB01
timestamp 1608910539
transform 1 0 14996 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_158
timestamp 1608910539
transform 1 0 15640 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_154
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_157
timestamp 1608910539
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 16008 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 16008 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1608910539
transform 1 0 1472 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1608910539
transform 1 0 2300 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3128 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1608910539
transform 1 0 3956 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1608910539
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1608910539
transform 1 0 6164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 6440 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 7636 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8464 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 9936 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1608910539
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11408 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1608910539
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1608910539
transform 1 0 13248 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1608910539
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 16008 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_13
timestamp 1608910539
transform 1 0 2300 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1608910539
transform 1 0 1472 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2392 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1608910539
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_46
timestamp 1608910539
transform 1 0 5336 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6440 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5428 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_76
timestamp 1608910539
transform 1 0 8096 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8372 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1608910539
transform 1 0 7268 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_96
timestamp 1608910539
transform 1 0 9936 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10212 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_108
timestamp 1608910539
transform 1 0 11040 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11316 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_139
timestamp 1608910539
transform 1 0 13892 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_127
timestamp 1608910539
transform 1 0 12788 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_158
timestamp 1608910539
transform 1 0 15640 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1608910539
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 16008 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_20
timestamp 1608910539
transform 1 0 2944 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_16
timestamp 1608910539
transform 1 0 2576 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 2024 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4692 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3220 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_55
timestamp 1608910539
transform 1 0 6164 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1608910539
transform 1 0 7084 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7176 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_17_100
timestamp 1608910539
transform 1 0 10304 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_84
timestamp 1608910539
transform 1 0 8832 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9936 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1608910539
transform 1 0 9108 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1608910539
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_112
timestamp 1608910539
transform 1 0 11408 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1608910539
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1608910539
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 16008 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_10
timestamp 1608910539
transform 1 0 2024 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_40
timestamp 1608910539
transform 1 0 4784 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_32
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1608910539
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_22
timestamp 1608910539
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5060 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5888 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_71
timestamp 1608910539
transform 1 0 7636 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 7360 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1608910539
transform 1 0 7912 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8740 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9844 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_125
timestamp 1608910539
transform 1 0 12604 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1608910539
transform 1 0 11316 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1608910539
transform 1 0 12144 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_137
timestamp 1608910539
transform 1 0 13708 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_158
timestamp 1608910539
transform 1 0 15640 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1608910539
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 16008 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_15
timestamp 1608910539
transform 1 0 2484 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1748 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_20_23
timestamp 1608910539
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_21
timestamp 1608910539
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1608910539
transform 1 0 3128 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1608910539
transform 1 0 3956 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4324 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 4968 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1608910539
transform 1 0 5244 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_60
timestamp 1608910539
transform 1 0 6624 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1608910539
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 5152 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 6716 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_20_77
timestamp 1608910539
transform 1 0 8188 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7636 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8464 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8464 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_99
timestamp 1608910539
transform 1 0 10212 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_95
timestamp 1608910539
transform 1 0 9844 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1608910539
transform 1 0 10304 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 9292 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_20_118
timestamp 1608910539
transform 1 0 11960 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1608910539
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_105
timestamp 1608910539
transform 1 0 10764 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11132 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1608910539
transform 1 0 10856 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_142
timestamp 1608910539
transform 1 0 14168 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_130
timestamp 1608910539
transform 1 0 13064 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1608910539
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_158
timestamp 1608910539
transform 1 0 15640 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_154
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1608910539
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1608910539
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 16008 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 16008 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_11
timestamp 1608910539
transform 1 0 2116 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2668 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4140 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_62
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1608910539
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_44
timestamp 1608910539
transform 1 0 5152 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 6072 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1608910539
transform 1 0 5244 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_79
timestamp 1608910539
transform 1 0 8372 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6900 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_100
timestamp 1608910539
transform 1 0 10304 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1608910539
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 10120 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1608910539
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_115
timestamp 1608910539
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10856 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1608910539
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_151
timestamp 1608910539
transform 1 0 14996 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 16008 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_16
timestamp 1608910539
transform 1 0 2576 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_10
timestamp 1608910539
transform 1 0 2024 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2668 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1608910539
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_26
timestamp 1608910539
transform 1 0 3496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5336 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1608910539
transform 1 0 6164 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_69
timestamp 1608910539
transform 1 0 7452 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7544 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608910539
transform 1 0 6992 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_102
timestamp 1608910539
transform 1 0 10488 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_88
timestamp 1608910539
transform 1 0 9200 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10580 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608910539
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_119
timestamp 1608910539
transform 1 0 12052 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1608910539
transform 1 0 12328 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1608910539
transform 1 0 13156 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1608910539
transform 1 0 15640 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1608910539
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1608910539
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_146
timestamp 1608910539
transform 1 0 14536 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 16008 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_10
timestamp 1608910539
transform 1 0 2024 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1608910539
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1608910539
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 2300 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1608910539
transform 1 0 3772 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1608910539
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5796 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1608910539
transform 1 0 4968 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1608910539
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8464 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7636 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1608910539
transform 1 0 10120 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1608910539
transform 1 0 9292 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1608910539
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10948 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1608910539
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608910539
transform 1 0 13248 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1608910539
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1608910539
transform -1 0 16008 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_10
timestamp 1608910539
transform 1 0 2024 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1608910539
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1608910539
transform 1 0 2944 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1608910539
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 1472 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608910539
transform 1 0 2576 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_46
timestamp 1608910539
transform 1 0 5336 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_43
timestamp 1608910539
transform 1 0 5060 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 6256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1608910539
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5428 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6440 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_78
timestamp 1608910539
transform 1 0 8280 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_right_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 8372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8648 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_104
timestamp 1608910539
transform 1 0 10672 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1608910539
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1608910539
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 10764 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1608910539
transform 1 0 11776 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10948 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1608910539
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1608910539
transform 1 0 14076 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1608910539
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_154
timestamp 1608910539
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1608910539
transform 1 0 14812 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_N_FTB01_A
timestamp 1608910539
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1608910539
transform -1 0 16008 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_13
timestamp 1608910539
transform 1 0 2300 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1608910539
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_N_FTB01_A
timestamp 1608910539
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1608910539
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clk_2_N_FTB01
timestamp 1608910539
transform 1 0 1564 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_21
timestamp 1608910539
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4600 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3128 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_54
timestamp 1608910539
transform 1 0 6072 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1608910539
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1608910539
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_71
timestamp 1608910539
transform 1 0 7636 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7728 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_25_104
timestamp 1608910539
transform 1 0 10672 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 9200 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_118
timestamp 1608910539
transform 1 0 11960 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1608910539
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10948 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_144
timestamp 1608910539
transform 1 0 14352 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_132
timestamp 1608910539
transform 1 0 13248 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_156
timestamp 1608910539
transform 1 0 15456 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1608910539
transform -1 0 16008 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1608910539
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1608910539
transform 1 0 1748 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1608910539
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1608910539
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1608910539
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  Test_en_W_FTB01
timestamp 1608910539
transform 1 0 1472 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01
timestamp 1608910539
transform 1 0 1840 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_16
timestamp 1608910539
transform 1 0 2576 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_N_FTB01_A
timestamp 1608910539
transform 1 0 2392 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_W_FTB01_A
timestamp 1608910539
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1608910539
transform 1 0 2024 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_20
timestamp 1608910539
transform 1 0 2944 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_20
timestamp 1608910539
transform 1 0 2944 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1608910539
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608910539
transform 1 0 3404 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608910539
transform 1 0 3036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_32
timestamp 1608910539
transform 1 0 4048 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_28
timestamp 1608910539
transform 1 0 3680 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1608910539
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1608910539
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1608910539
transform 1 0 3956 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1608910539
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608910539
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_38
timestamp 1608910539
transform 1 0 4600 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1608910539
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608910539
transform 1 0 4876 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608910539
transform 1 0 4784 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608910539
transform 1 0 4416 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_49
timestamp 1608910539
transform 1 0 5612 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1608910539
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608910539
transform 1 0 5704 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608910539
transform 1 0 5244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1608910539
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1608910539
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1608910539
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1608910539
transform 1 0 6624 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1608910539
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608910539
transform 1 0 6808 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5336 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_26_70
timestamp 1608910539
transform 1 0 7544 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1608910539
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608910539
transform 1 0 7268 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608910539
transform 1 0 6900 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608910539
transform 1 0 7176 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608910539
transform 1 0 7636 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_79
timestamp 1608910539
transform 1 0 8372 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_79
timestamp 1608910539
transform 1 0 8372 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1608910539
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1608910539
transform 1 0 8464 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608910539
transform 1 0 8464 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608910539
transform 1 0 8004 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608910539
transform 1 0 8004 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_92
timestamp 1608910539
transform 1 0 9568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1608910539
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1608910539
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1608910539
transform 1 0 9292 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1608910539
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1608910539
transform 1 0 9660 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1608910539
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608910539
transform 1 0 9200 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_98
timestamp 1608910539
transform 1 0 10120 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1608910539
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1608910539
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608910539
transform 1 0 10672 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1608910539
transform 1 0 12604 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_122
timestamp 1608910539
transform 1 0 12328 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1608910539
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_111
timestamp 1608910539
transform 1 0 11316 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1608910539
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1608910539
transform 1 0 12512 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 11408 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_27_145
timestamp 1608910539
transform 1 0 14444 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_137
timestamp 1608910539
transform 1 0 13708 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_142
timestamp 1608910539
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_134
timestamp 1608910539
transform 1 0 13432 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1608910539
transform 1 0 13248 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1608910539
transform 1 0 14352 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608910539
transform 1 0 12880 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1608910539
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_N_FTB01_A
timestamp 1608910539
transform 1 0 15088 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_N_FTB01_A
timestamp 1608910539
transform 1 0 14904 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1608910539
transform 1 0 14536 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_156
timestamp 1608910539
transform 1 0 15456 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_154
timestamp 1608910539
transform 1 0 15272 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp 1608910539
transform 1 0 15640 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1608910539
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1608910539
transform 1 0 15364 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1608910539
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1608910539
transform -1 0 16008 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1608910539
transform -1 0 16008 0 -1 16864
box -38 -48 314 592
<< labels >>
rlabel metal3 s 16400 16600 17200 16720 6 Test_en_E_in
port 0 nsew signal input
rlabel metal3 s 16400 9936 17200 10056 6 Test_en_E_out
port 1 nsew signal tristate
rlabel metal2 s 2042 19200 2098 20000 6 Test_en_N_out
port 2 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 Test_en_S_in
port 3 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 Test_en_W_in
port 4 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 Test_en_W_out
port 5 nsew signal tristate
rlabel metal3 s 0 416 800 536 6 ccff_head
port 6 nsew signal input
rlabel metal3 s 16400 3272 17200 3392 6 ccff_tail
port 7 nsew signal tristate
rlabel metal2 s 6918 0 6974 800 6 chany_bottom_in[0]
port 8 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 chany_bottom_in[10]
port 9 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 chany_bottom_in[11]
port 10 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[12]
port 11 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[13]
port 12 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[14]
port 13 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_in[15]
port 14 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 chany_bottom_in[16]
port 15 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_in[17]
port 16 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_in[18]
port 17 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_in[19]
port 18 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[1]
port 19 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[2]
port 20 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 chany_bottom_in[3]
port 21 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_in[4]
port 22 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[5]
port 23 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[6]
port 24 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 chany_bottom_in[7]
port 25 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 chany_bottom_in[8]
port 26 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[9]
port 27 nsew signal input
rlabel metal2 s 110 0 166 800 6 chany_bottom_out[0]
port 28 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 chany_bottom_out[10]
port 29 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_out[11]
port 30 nsew signal tristate
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_out[12]
port 31 nsew signal tristate
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_out[13]
port 32 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 chany_bottom_out[14]
port 33 nsew signal tristate
rlabel metal2 s 5262 0 5318 800 6 chany_bottom_out[15]
port 34 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_out[16]
port 35 nsew signal tristate
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_out[17]
port 36 nsew signal tristate
rlabel metal2 s 6274 0 6330 800 6 chany_bottom_out[18]
port 37 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_out[19]
port 38 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 chany_bottom_out[1]
port 39 nsew signal tristate
rlabel metal2 s 754 0 810 800 6 chany_bottom_out[2]
port 40 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 chany_bottom_out[3]
port 41 nsew signal tristate
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_out[4]
port 42 nsew signal tristate
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_out[5]
port 43 nsew signal tristate
rlabel metal2 s 2134 0 2190 800 6 chany_bottom_out[6]
port 44 nsew signal tristate
rlabel metal2 s 2502 0 2558 800 6 chany_bottom_out[7]
port 45 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 chany_bottom_out[8]
port 46 nsew signal tristate
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_out[9]
port 47 nsew signal tristate
rlabel metal2 s 9862 19200 9918 20000 6 chany_top_in[0]
port 48 nsew signal input
rlabel metal2 s 13634 19200 13690 20000 6 chany_top_in[10]
port 49 nsew signal input
rlabel metal2 s 14002 19200 14058 20000 6 chany_top_in[11]
port 50 nsew signal input
rlabel metal2 s 14370 19200 14426 20000 6 chany_top_in[12]
port 51 nsew signal input
rlabel metal2 s 14738 19200 14794 20000 6 chany_top_in[13]
port 52 nsew signal input
rlabel metal2 s 15106 19200 15162 20000 6 chany_top_in[14]
port 53 nsew signal input
rlabel metal2 s 15474 19200 15530 20000 6 chany_top_in[15]
port 54 nsew signal input
rlabel metal2 s 15842 19200 15898 20000 6 chany_top_in[16]
port 55 nsew signal input
rlabel metal2 s 16210 19200 16266 20000 6 chany_top_in[17]
port 56 nsew signal input
rlabel metal2 s 16578 19200 16634 20000 6 chany_top_in[18]
port 57 nsew signal input
rlabel metal2 s 16946 19200 17002 20000 6 chany_top_in[19]
port 58 nsew signal input
rlabel metal2 s 10230 19200 10286 20000 6 chany_top_in[1]
port 59 nsew signal input
rlabel metal2 s 10598 19200 10654 20000 6 chany_top_in[2]
port 60 nsew signal input
rlabel metal2 s 10966 19200 11022 20000 6 chany_top_in[3]
port 61 nsew signal input
rlabel metal2 s 11334 19200 11390 20000 6 chany_top_in[4]
port 62 nsew signal input
rlabel metal2 s 11794 19200 11850 20000 6 chany_top_in[5]
port 63 nsew signal input
rlabel metal2 s 12162 19200 12218 20000 6 chany_top_in[6]
port 64 nsew signal input
rlabel metal2 s 12530 19200 12586 20000 6 chany_top_in[7]
port 65 nsew signal input
rlabel metal2 s 12898 19200 12954 20000 6 chany_top_in[8]
port 66 nsew signal input
rlabel metal2 s 13266 19200 13322 20000 6 chany_top_in[9]
port 67 nsew signal input
rlabel metal2 s 2410 19200 2466 20000 6 chany_top_out[0]
port 68 nsew signal tristate
rlabel metal2 s 6182 19200 6238 20000 6 chany_top_out[10]
port 69 nsew signal tristate
rlabel metal2 s 6550 19200 6606 20000 6 chany_top_out[11]
port 70 nsew signal tristate
rlabel metal2 s 6918 19200 6974 20000 6 chany_top_out[12]
port 71 nsew signal tristate
rlabel metal2 s 7286 19200 7342 20000 6 chany_top_out[13]
port 72 nsew signal tristate
rlabel metal2 s 7654 19200 7710 20000 6 chany_top_out[14]
port 73 nsew signal tristate
rlabel metal2 s 8022 19200 8078 20000 6 chany_top_out[15]
port 74 nsew signal tristate
rlabel metal2 s 8390 19200 8446 20000 6 chany_top_out[16]
port 75 nsew signal tristate
rlabel metal2 s 8758 19200 8814 20000 6 chany_top_out[17]
port 76 nsew signal tristate
rlabel metal2 s 9126 19200 9182 20000 6 chany_top_out[18]
port 77 nsew signal tristate
rlabel metal2 s 9494 19200 9550 20000 6 chany_top_out[19]
port 78 nsew signal tristate
rlabel metal2 s 2778 19200 2834 20000 6 chany_top_out[1]
port 79 nsew signal tristate
rlabel metal2 s 3146 19200 3202 20000 6 chany_top_out[2]
port 80 nsew signal tristate
rlabel metal2 s 3514 19200 3570 20000 6 chany_top_out[3]
port 81 nsew signal tristate
rlabel metal2 s 3882 19200 3938 20000 6 chany_top_out[4]
port 82 nsew signal tristate
rlabel metal2 s 4250 19200 4306 20000 6 chany_top_out[5]
port 83 nsew signal tristate
rlabel metal2 s 4618 19200 4674 20000 6 chany_top_out[6]
port 84 nsew signal tristate
rlabel metal2 s 4986 19200 5042 20000 6 chany_top_out[7]
port 85 nsew signal tristate
rlabel metal2 s 5354 19200 5410 20000 6 chany_top_out[8]
port 86 nsew signal tristate
rlabel metal2 s 5722 19200 5778 20000 6 chany_top_out[9]
port 87 nsew signal tristate
rlabel metal2 s 202 19200 258 20000 6 clk_2_N_out
port 88 nsew signal tristate
rlabel metal2 s 14186 0 14242 800 6 clk_2_S_in
port 89 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 clk_2_S_out
port 90 nsew signal tristate
rlabel metal2 s 570 19200 626 20000 6 clk_3_N_out
port 91 nsew signal tristate
rlabel metal2 s 14554 0 14610 800 6 clk_3_S_in
port 92 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 clk_3_S_out
port 93 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 left_grid_pin_16_
port 94 nsew signal tristate
rlabel metal3 s 0 2320 800 2440 6 left_grid_pin_17_
port 95 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 left_grid_pin_18_
port 96 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 left_grid_pin_19_
port 97 nsew signal tristate
rlabel metal3 s 0 5312 800 5432 6 left_grid_pin_20_
port 98 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 left_grid_pin_21_
port 99 nsew signal tristate
rlabel metal3 s 0 7352 800 7472 6 left_grid_pin_22_
port 100 nsew signal tristate
rlabel metal3 s 0 8304 800 8424 6 left_grid_pin_23_
port 101 nsew signal tristate
rlabel metal3 s 0 9392 800 9512 6 left_grid_pin_24_
port 102 nsew signal tristate
rlabel metal3 s 0 10344 800 10464 6 left_grid_pin_25_
port 103 nsew signal tristate
rlabel metal3 s 0 11296 800 11416 6 left_grid_pin_26_
port 104 nsew signal tristate
rlabel metal3 s 0 12384 800 12504 6 left_grid_pin_27_
port 105 nsew signal tristate
rlabel metal3 s 0 13336 800 13456 6 left_grid_pin_28_
port 106 nsew signal tristate
rlabel metal3 s 0 14288 800 14408 6 left_grid_pin_29_
port 107 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 left_grid_pin_30_
port 108 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 left_grid_pin_31_
port 109 nsew signal tristate
rlabel metal2 s 938 19200 994 20000 6 prog_clk_0_N_out
port 110 nsew signal tristate
rlabel metal2 s 16210 0 16266 800 6 prog_clk_0_S_out
port 111 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 prog_clk_0_W_in
port 112 nsew signal input
rlabel metal2 s 1306 19200 1362 20000 6 prog_clk_2_N_out
port 113 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 prog_clk_2_S_in
port 114 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 prog_clk_2_S_out
port 115 nsew signal tristate
rlabel metal2 s 1674 19200 1730 20000 6 prog_clk_3_N_out
port 116 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 prog_clk_3_S_in
port 117 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 prog_clk_3_S_out
port 118 nsew signal tristate
rlabel metal4 s 13437 2128 13757 17456 6 VPWR
port 119 nsew power bidirectional
rlabel metal4 s 8440 2128 8760 17456 6 VPWR
port 120 nsew power bidirectional
rlabel metal4 s 3443 2128 3763 17456 6 VPWR
port 121 nsew power bidirectional
rlabel metal4 s 10939 2128 11259 17456 6 VGND
port 122 nsew ground bidirectional
rlabel metal4 s 5941 2128 6261 17456 6 VGND
port 123 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
